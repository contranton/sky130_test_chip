magic
tech sky130A
magscale 1 2
timestamp 1640660821
<< nwell >>
rect 82712 687217 85064 687251
rect 119210 593040 120330 593330
rect 119250 583500 120370 583790
rect 119290 574480 120410 574770
rect 119240 566810 120360 567100
rect 312162 561428 312200 561514
rect 437482 561428 437520 561514
rect 119240 560270 120360 560560
rect 312162 560340 312200 560436
rect 437482 560340 437520 560436
rect 435312 559896 435350 559992
rect 560632 559896 560670 559992
rect 312162 559252 312200 559348
rect 437482 559252 437520 559348
rect 435312 558808 435350 558904
rect 560632 558808 560670 558904
rect 312162 558164 312200 558260
rect 437482 558164 437520 558260
rect 435312 557720 435350 557816
rect 560632 557720 560670 557816
rect 312162 557076 312200 557172
rect 437482 557076 437520 557172
rect 435312 556632 435350 556728
rect 560632 556632 560670 556728
rect 312162 555988 312200 556084
rect 437482 555988 437520 556084
rect 435312 555544 435350 555640
rect 560632 555544 560670 555640
rect 312162 554900 312200 554996
rect 437482 554900 437520 554996
rect 435312 554456 435350 554552
rect 560632 554456 560670 554552
rect 312162 553812 312200 553908
rect 437482 553812 437520 553908
rect 119310 553440 120430 553730
rect 435312 553368 435350 553464
rect 560632 553368 560670 553464
rect 312162 552724 312200 552820
rect 437482 552724 437520 552820
rect 435312 552280 435350 552376
rect 560632 552280 560670 552376
rect 312162 551636 312200 551732
rect 437482 551636 437520 551732
rect 435312 551192 435350 551288
rect 560632 551192 560670 551288
rect 312162 550548 312200 550644
rect 437482 550548 437520 550644
rect 435312 550104 435350 550200
rect 560632 550104 560670 550200
rect 312162 549460 312200 549556
rect 437482 549460 437520 549556
rect 435312 549016 435350 549112
rect 560632 549016 560670 549112
rect 312162 548372 312200 548468
rect 437482 548372 437520 548468
rect 435312 547928 435350 548024
rect 560632 547928 560670 548024
rect 312162 547284 312200 547380
rect 437482 547284 437520 547380
rect 435312 546840 435350 546936
rect 560632 546840 560670 546936
rect 312162 546196 312200 546292
rect 437482 546196 437520 546292
rect 119310 545870 120430 546160
rect 435312 545752 435350 545848
rect 560632 545752 560670 545848
rect 312162 545108 312200 545204
rect 437482 545108 437520 545204
rect 435312 544664 435350 544760
rect 560632 544664 560670 544760
rect 312162 544020 312200 544116
rect 437482 544020 437520 544116
rect 435312 543576 435350 543672
rect 560632 543576 560670 543672
rect 312162 542932 312200 543028
rect 437482 542932 437520 543028
rect 435312 542488 435350 542584
rect 560632 542488 560670 542584
rect 312162 541844 312200 541940
rect 437482 541844 437520 541940
rect 435312 541400 435350 541496
rect 560632 541400 560670 541496
rect 312162 540756 312200 540852
rect 437482 540756 437520 540852
rect 435312 540312 435350 540408
rect 560632 540312 560670 540408
rect 312162 539668 312200 539764
rect 437482 539668 437520 539764
rect 435312 539224 435350 539320
rect 560632 539224 560670 539320
rect 312162 538580 312200 538676
rect 437482 538580 437520 538676
rect 435312 538136 435350 538232
rect 560632 538136 560670 538232
rect 119280 537810 120400 538100
rect 312162 537492 312200 537588
rect 437482 537492 437520 537588
rect 435312 537048 435350 537144
rect 560632 537048 560670 537144
rect 312162 536404 312200 536500
rect 437482 536404 437520 536500
rect 435312 535960 435350 536056
rect 560632 535960 560670 536056
rect 312162 535316 312200 535412
rect 437482 535316 437520 535412
rect 435312 534872 435350 534968
rect 560632 534872 560670 534968
rect 312162 534228 312200 534324
rect 437482 534228 437520 534324
rect 435312 533784 435350 533880
rect 560632 533784 560670 533880
rect 312162 533140 312200 533236
rect 437482 533140 437520 533236
rect 435312 532696 435350 532792
rect 560632 532696 560670 532792
rect 312162 532052 312200 532148
rect 437482 532052 437520 532148
rect 435312 531608 435350 531704
rect 560632 531608 560670 531704
rect 312162 530964 312200 531060
rect 437482 530964 437520 531060
rect 435312 530520 435350 530616
rect 560632 530520 560670 530616
rect 312162 529876 312200 529972
rect 437482 529876 437520 529972
rect 435312 529432 435350 529528
rect 560632 529432 560670 529528
rect 312162 528788 312200 528884
rect 437482 528788 437520 528884
rect 435312 528344 435350 528440
rect 560632 528344 560670 528440
rect 312162 527700 312200 527796
rect 437482 527700 437520 527796
rect 435312 527256 435350 527352
rect 560632 527256 560670 527352
rect 312162 526612 312200 526708
rect 437482 526612 437520 526708
rect 435312 526168 435350 526264
rect 560632 526168 560670 526264
rect 312162 525524 312200 525620
rect 437482 525524 437520 525620
rect 435312 525080 435350 525176
rect 560632 525080 560670 525176
rect 312162 524436 312200 524532
rect 437482 524436 437520 524532
rect 435312 523992 435350 524088
rect 560632 523992 560670 524088
rect 312162 523348 312200 523444
rect 437482 523348 437520 523444
rect 435312 522904 435350 523000
rect 560632 522904 560670 523000
rect 312162 522260 312200 522356
rect 437482 522260 437520 522356
rect 435312 521816 435350 521912
rect 560632 521816 560670 521912
rect 312162 521172 312200 521268
rect 437482 521172 437520 521268
rect 435312 520728 435350 520824
rect 560632 520728 560670 520824
rect 312162 520084 312200 520180
rect 437482 520084 437520 520180
rect 435312 519640 435350 519736
rect 560632 519640 560670 519736
rect 312162 518996 312200 519092
rect 437482 518996 437520 519092
rect 435312 518552 435350 518648
rect 560632 518552 560670 518648
rect 312162 517908 312200 518004
rect 437482 517908 437520 518004
rect 435312 517464 435350 517560
rect 560632 517464 560670 517560
rect 312162 516820 312200 516916
rect 437482 516820 437520 516916
rect 435312 516376 435350 516472
rect 560632 516376 560670 516472
rect 312162 515732 312200 515828
rect 437482 515732 437520 515828
rect 435312 515288 435350 515384
rect 560632 515288 560670 515384
rect 312162 514644 312200 514740
rect 437482 514644 437520 514740
rect 435312 514200 435350 514296
rect 560632 514200 560670 514296
rect 312162 513556 312200 513652
rect 437482 513556 437520 513652
rect 435312 513112 435350 513208
rect 560632 513112 560670 513208
rect 312162 512468 312200 512564
rect 437482 512468 437520 512564
rect 435312 512024 435350 512120
rect 560632 512024 560670 512120
rect 312162 511380 312200 511476
rect 437482 511380 437520 511476
rect 435312 510936 435350 511032
rect 560632 510936 560670 511032
rect 312162 510292 312200 510388
rect 437482 510292 437520 510388
rect 435312 509848 435350 509944
rect 560632 509848 560670 509944
rect 312162 509204 312200 509300
rect 437482 509204 437520 509300
rect 435312 508760 435350 508856
rect 560632 508760 560670 508856
rect 312162 508116 312200 508212
rect 437482 508116 437520 508212
rect 435312 507672 435350 507768
rect 560632 507672 560670 507768
rect 312162 507028 312200 507124
rect 437482 507028 437520 507124
rect 435312 506584 435350 506680
rect 560632 506584 560670 506680
rect 312162 505940 312200 506036
rect 437482 505940 437520 506036
rect 435312 505496 435350 505592
rect 560632 505496 560670 505592
rect 312162 504852 312200 504948
rect 437482 504852 437520 504948
rect 435312 504408 435350 504504
rect 560632 504408 560670 504504
rect 435312 503330 435350 503416
rect 560632 503330 560670 503416
rect 312162 498768 312200 498854
rect 437482 498768 437520 498854
rect 312162 497680 312200 497776
rect 437482 497680 437520 497776
rect 435312 497236 435350 497332
rect 560632 497236 560670 497332
rect 312162 496592 312200 496688
rect 437482 496592 437520 496688
rect 435312 496148 435350 496244
rect 560632 496148 560670 496244
rect 312162 495504 312200 495600
rect 437482 495504 437520 495600
rect 435312 495060 435350 495156
rect 560632 495060 560670 495156
rect 312162 494416 312200 494512
rect 437482 494416 437520 494512
rect 435312 493972 435350 494068
rect 560632 493972 560670 494068
rect 312162 493328 312200 493424
rect 437482 493328 437520 493424
rect 435312 492884 435350 492980
rect 560632 492884 560670 492980
rect 312162 492240 312200 492336
rect 437482 492240 437520 492336
rect 435312 491796 435350 491892
rect 560632 491796 560670 491892
rect 312162 491152 312200 491248
rect 437482 491152 437520 491248
rect 435312 490708 435350 490804
rect 560632 490708 560670 490804
rect 312162 490064 312200 490160
rect 437482 490064 437520 490160
rect 435312 489620 435350 489716
rect 560632 489620 560670 489716
rect 312162 488976 312200 489072
rect 437482 488976 437520 489072
rect 435312 488532 435350 488628
rect 560632 488532 560670 488628
rect 312162 487888 312200 487984
rect 437482 487888 437520 487984
rect 435312 487444 435350 487540
rect 560632 487444 560670 487540
rect 312162 486800 312200 486896
rect 437482 486800 437520 486896
rect 435312 486356 435350 486452
rect 560632 486356 560670 486452
rect 312162 485712 312200 485808
rect 437482 485712 437520 485808
rect 435312 485268 435350 485364
rect 560632 485268 560670 485364
rect 312162 484624 312200 484720
rect 437482 484624 437520 484720
rect 435312 484180 435350 484276
rect 560632 484180 560670 484276
rect 312162 483536 312200 483632
rect 437482 483536 437520 483632
rect 435312 483092 435350 483188
rect 560632 483092 560670 483188
rect 312162 482448 312200 482544
rect 437482 482448 437520 482544
rect 435312 482004 435350 482100
rect 560632 482004 560670 482100
rect 312162 481360 312200 481456
rect 437482 481360 437520 481456
rect 435312 480916 435350 481012
rect 560632 480916 560670 481012
rect 312162 480272 312200 480368
rect 437482 480272 437520 480368
rect 435312 479828 435350 479924
rect 560632 479828 560670 479924
rect 312162 479184 312200 479280
rect 437482 479184 437520 479280
rect 435312 478740 435350 478836
rect 560632 478740 560670 478836
rect 312162 478096 312200 478192
rect 437482 478096 437520 478192
rect 435312 477652 435350 477748
rect 560632 477652 560670 477748
rect 312162 477008 312200 477104
rect 437482 477008 437520 477104
rect 435312 476564 435350 476660
rect 560632 476564 560670 476660
rect 312162 475920 312200 476016
rect 437482 475920 437520 476016
rect 435312 475476 435350 475572
rect 560632 475476 560670 475572
rect 312162 474832 312200 474928
rect 437482 474832 437520 474928
rect 435312 474388 435350 474484
rect 560632 474388 560670 474484
rect 312162 473744 312200 473840
rect 437482 473744 437520 473840
rect 435312 473300 435350 473396
rect 560632 473300 560670 473396
rect 312162 472656 312200 472752
rect 437482 472656 437520 472752
rect 435312 472212 435350 472308
rect 560632 472212 560670 472308
rect 312162 471568 312200 471664
rect 437482 471568 437520 471664
rect 435312 471124 435350 471220
rect 560632 471124 560670 471220
rect 312162 470480 312200 470576
rect 437482 470480 437520 470576
rect 435312 470036 435350 470132
rect 560632 470036 560670 470132
rect 312162 469392 312200 469488
rect 437482 469392 437520 469488
rect 435312 468948 435350 469044
rect 560632 468948 560670 469044
rect 312162 468304 312200 468400
rect 437482 468304 437520 468400
rect 435312 467860 435350 467956
rect 560632 467860 560670 467956
rect 312162 467216 312200 467312
rect 437482 467216 437520 467312
rect 435312 466772 435350 466868
rect 560632 466772 560670 466868
rect 312162 466128 312200 466224
rect 437482 466128 437520 466224
rect 435312 465684 435350 465780
rect 560632 465684 560670 465780
rect 312162 465040 312200 465136
rect 437482 465040 437520 465136
rect 435312 464596 435350 464692
rect 560632 464596 560670 464692
rect 312162 463952 312200 464048
rect 437482 463952 437520 464048
rect 435312 463508 435350 463604
rect 560632 463508 560670 463604
rect 312162 462864 312200 462960
rect 437482 462864 437520 462960
rect 435312 462420 435350 462516
rect 560632 462420 560670 462516
rect 312162 461776 312200 461872
rect 437482 461776 437520 461872
rect 435312 461332 435350 461428
rect 560632 461332 560670 461428
rect 312162 460688 312200 460784
rect 437482 460688 437520 460784
rect 435312 460244 435350 460340
rect 560632 460244 560670 460340
rect 312162 459600 312200 459696
rect 437482 459600 437520 459696
rect 435312 459156 435350 459252
rect 560632 459156 560670 459252
rect 312162 458512 312200 458608
rect 437482 458512 437520 458608
rect 435312 458068 435350 458164
rect 560632 458068 560670 458164
rect 312162 457424 312200 457520
rect 437482 457424 437520 457520
rect 435312 456980 435350 457076
rect 560632 456980 560670 457076
rect 312162 456336 312200 456432
rect 437482 456336 437520 456432
rect 435312 455892 435350 455988
rect 560632 455892 560670 455988
rect 312162 455248 312200 455344
rect 437482 455248 437520 455344
rect 435312 454804 435350 454900
rect 560632 454804 560670 454900
rect 312162 454160 312200 454256
rect 437482 454160 437520 454256
rect 435312 453716 435350 453812
rect 560632 453716 560670 453812
rect 312162 453072 312200 453168
rect 437482 453072 437520 453168
rect 435312 452628 435350 452724
rect 560632 452628 560670 452724
rect 312162 451984 312200 452080
rect 437482 451984 437520 452080
rect 435312 451540 435350 451636
rect 560632 451540 560670 451636
rect 312162 450896 312200 450992
rect 437482 450896 437520 450992
rect 435312 450452 435350 450548
rect 560632 450452 560670 450548
rect 312162 449808 312200 449904
rect 437482 449808 437520 449904
rect 435312 449364 435350 449460
rect 560632 449364 560670 449460
rect 312162 448720 312200 448816
rect 437482 448720 437520 448816
rect 435312 448276 435350 448372
rect 560632 448276 560670 448372
rect 312162 447632 312200 447728
rect 437482 447632 437520 447728
rect 435312 447188 435350 447284
rect 560632 447188 560670 447284
rect 312162 446544 312200 446640
rect 437482 446544 437520 446640
rect 435312 446100 435350 446196
rect 560632 446100 560670 446196
rect 312162 445456 312200 445552
rect 437482 445456 437520 445552
rect 435312 445012 435350 445108
rect 560632 445012 560670 445108
rect 312162 444368 312200 444464
rect 437482 444368 437520 444464
rect 435312 443924 435350 444020
rect 560632 443924 560670 444020
rect 312162 443280 312200 443376
rect 437482 443280 437520 443376
rect 435312 442836 435350 442932
rect 560632 442836 560670 442932
rect 312162 442192 312200 442288
rect 437482 442192 437520 442288
rect 435312 441748 435350 441844
rect 560632 441748 560670 441844
rect 435312 440670 435350 440756
rect 560632 440670 560670 440756
rect 312162 436108 312200 436194
rect 437482 436108 437520 436194
rect 312162 435020 312200 435116
rect 437482 435020 437520 435116
rect 435312 434576 435350 434672
rect 560632 434576 560670 434672
rect 312162 433932 312200 434028
rect 437482 433932 437520 434028
rect 435312 433488 435350 433584
rect 560632 433488 560670 433584
rect 312162 432844 312200 432940
rect 437482 432844 437520 432940
rect 435312 432400 435350 432496
rect 560632 432400 560670 432496
rect 312162 431756 312200 431852
rect 437482 431756 437520 431852
rect 435312 431312 435350 431408
rect 560632 431312 560670 431408
rect 312162 430668 312200 430764
rect 437482 430668 437520 430764
rect 435312 430224 435350 430320
rect 560632 430224 560670 430320
rect 312162 429580 312200 429676
rect 437482 429580 437520 429676
rect 435312 429136 435350 429232
rect 560632 429136 560670 429232
rect 312162 428492 312200 428588
rect 437482 428492 437520 428588
rect 435312 428048 435350 428144
rect 560632 428048 560670 428144
rect 312162 427404 312200 427500
rect 437482 427404 437520 427500
rect 435312 426960 435350 427056
rect 560632 426960 560670 427056
rect 312162 426316 312200 426412
rect 437482 426316 437520 426412
rect 435312 425872 435350 425968
rect 560632 425872 560670 425968
rect 312162 425228 312200 425324
rect 437482 425228 437520 425324
rect 435312 424784 435350 424880
rect 560632 424784 560670 424880
rect 312162 424140 312200 424236
rect 437482 424140 437520 424236
rect 435312 423696 435350 423792
rect 560632 423696 560670 423792
rect 312162 423052 312200 423148
rect 437482 423052 437520 423148
rect 435312 422608 435350 422704
rect 560632 422608 560670 422704
rect 312162 421964 312200 422060
rect 437482 421964 437520 422060
rect 435312 421520 435350 421616
rect 560632 421520 560670 421616
rect 312162 420876 312200 420972
rect 437482 420876 437520 420972
rect 435312 420432 435350 420528
rect 560632 420432 560670 420528
rect 312162 419788 312200 419884
rect 437482 419788 437520 419884
rect 435312 419344 435350 419440
rect 560632 419344 560670 419440
rect 312162 418700 312200 418796
rect 437482 418700 437520 418796
rect 435312 418256 435350 418352
rect 560632 418256 560670 418352
rect 312162 417612 312200 417708
rect 437482 417612 437520 417708
rect 435312 417168 435350 417264
rect 560632 417168 560670 417264
rect 312162 416524 312200 416620
rect 437482 416524 437520 416620
rect 435312 416080 435350 416176
rect 560632 416080 560670 416176
rect 312162 415436 312200 415532
rect 437482 415436 437520 415532
rect 435312 414992 435350 415088
rect 560632 414992 560670 415088
rect 312162 414348 312200 414444
rect 437482 414348 437520 414444
rect 435312 413904 435350 414000
rect 560632 413904 560670 414000
rect 312162 413260 312200 413356
rect 437482 413260 437520 413356
rect 435312 412816 435350 412912
rect 560632 412816 560670 412912
rect 312162 412172 312200 412268
rect 437482 412172 437520 412268
rect 435312 411728 435350 411824
rect 560632 411728 560670 411824
rect 312162 411084 312200 411180
rect 437482 411084 437520 411180
rect 435312 410640 435350 410736
rect 560632 410640 560670 410736
rect 312162 409996 312200 410092
rect 437482 409996 437520 410092
rect 435312 409552 435350 409648
rect 560632 409552 560670 409648
rect 312162 408908 312200 409004
rect 437482 408908 437520 409004
rect 435312 408464 435350 408560
rect 560632 408464 560670 408560
rect 312162 407820 312200 407916
rect 437482 407820 437520 407916
rect 435312 407376 435350 407472
rect 560632 407376 560670 407472
rect 312162 406732 312200 406828
rect 437482 406732 437520 406828
rect 435312 406288 435350 406384
rect 560632 406288 560670 406384
rect 312162 405644 312200 405740
rect 437482 405644 437520 405740
rect 435312 405200 435350 405296
rect 560632 405200 560670 405296
rect 312162 404556 312200 404652
rect 437482 404556 437520 404652
rect 435312 404112 435350 404208
rect 560632 404112 560670 404208
rect 312162 403468 312200 403564
rect 437482 403468 437520 403564
rect 435312 403024 435350 403120
rect 560632 403024 560670 403120
rect 312162 402380 312200 402476
rect 437482 402380 437520 402476
rect 435312 401936 435350 402032
rect 560632 401936 560670 402032
rect 312162 401292 312200 401388
rect 437482 401292 437520 401388
rect 435312 400848 435350 400944
rect 560632 400848 560670 400944
rect 312162 400204 312200 400300
rect 437482 400204 437520 400300
rect 435312 399760 435350 399856
rect 560632 399760 560670 399856
rect 312162 399116 312200 399212
rect 437482 399116 437520 399212
rect 435312 398672 435350 398768
rect 560632 398672 560670 398768
rect 312162 398028 312200 398124
rect 437482 398028 437520 398124
rect 435312 397584 435350 397680
rect 560632 397584 560670 397680
rect 312162 396940 312200 397036
rect 437482 396940 437520 397036
rect 435312 396496 435350 396592
rect 560632 396496 560670 396592
rect 312162 395852 312200 395948
rect 437482 395852 437520 395948
rect 435312 395408 435350 395504
rect 560632 395408 560670 395504
rect 312162 394764 312200 394860
rect 437482 394764 437520 394860
rect 435312 394320 435350 394416
rect 560632 394320 560670 394416
rect 312162 393676 312200 393772
rect 437482 393676 437520 393772
rect 435312 393232 435350 393328
rect 560632 393232 560670 393328
rect 312162 392588 312200 392684
rect 437482 392588 437520 392684
rect 435312 392144 435350 392240
rect 560632 392144 560670 392240
rect 312162 391500 312200 391596
rect 437482 391500 437520 391596
rect 435312 391056 435350 391152
rect 560632 391056 560670 391152
rect 312162 390412 312200 390508
rect 437482 390412 437520 390508
rect 435312 389968 435350 390064
rect 560632 389968 560670 390064
rect 312162 389324 312200 389420
rect 437482 389324 437520 389420
rect 435312 388880 435350 388976
rect 560632 388880 560670 388976
rect 312162 388236 312200 388332
rect 437482 388236 437520 388332
rect 435312 387792 435350 387888
rect 560632 387792 560670 387888
rect 312162 387148 312200 387244
rect 437482 387148 437520 387244
rect 435312 386704 435350 386800
rect 560632 386704 560670 386800
rect 312162 386060 312200 386156
rect 437482 386060 437520 386156
rect 435312 385616 435350 385712
rect 560632 385616 560670 385712
rect 312162 384972 312200 385068
rect 437482 384972 437520 385068
rect 435312 384528 435350 384624
rect 560632 384528 560670 384624
rect 312162 383884 312200 383980
rect 437482 383884 437520 383980
rect 435312 383440 435350 383536
rect 560632 383440 560670 383536
rect 312162 382796 312200 382892
rect 437482 382796 437520 382892
rect 435312 382352 435350 382448
rect 560632 382352 560670 382448
rect 312162 381708 312200 381804
rect 437482 381708 437520 381804
rect 435312 381264 435350 381360
rect 560632 381264 560670 381360
rect 312162 380620 312200 380716
rect 437482 380620 437520 380716
rect 435312 380176 435350 380272
rect 560632 380176 560670 380272
rect 312162 379532 312200 379628
rect 437482 379532 437520 379628
rect 435312 379088 435350 379184
rect 560632 379088 560670 379184
rect 435312 378010 435350 378096
rect 560632 378010 560670 378096
rect 312162 373448 312200 373534
rect 437482 373448 437520 373534
rect 312162 372360 312200 372456
rect 437482 372360 437520 372456
rect 435312 371916 435350 372012
rect 560632 371916 560670 372012
rect 312162 371272 312200 371368
rect 437482 371272 437520 371368
rect 435312 370828 435350 370924
rect 560632 370828 560670 370924
rect 312162 370184 312200 370280
rect 437482 370184 437520 370280
rect 435312 369740 435350 369836
rect 560632 369740 560670 369836
rect 312162 369096 312200 369192
rect 437482 369096 437520 369192
rect 435312 368652 435350 368748
rect 560632 368652 560670 368748
rect 312162 368008 312200 368104
rect 437482 368008 437520 368104
rect 435312 367564 435350 367660
rect 560632 367564 560670 367660
rect 312162 366920 312200 367016
rect 437482 366920 437520 367016
rect 435312 366476 435350 366572
rect 560632 366476 560670 366572
rect 312162 365832 312200 365928
rect 437482 365832 437520 365928
rect 435312 365388 435350 365484
rect 560632 365388 560670 365484
rect 312162 364744 312200 364840
rect 437482 364744 437520 364840
rect 435312 364300 435350 364396
rect 560632 364300 560670 364396
rect 312162 363656 312200 363752
rect 437482 363656 437520 363752
rect 435312 363212 435350 363308
rect 560632 363212 560670 363308
rect 312162 362568 312200 362664
rect 437482 362568 437520 362664
rect 435312 362124 435350 362220
rect 560632 362124 560670 362220
rect 312162 361480 312200 361576
rect 437482 361480 437520 361576
rect 435312 361036 435350 361132
rect 560632 361036 560670 361132
rect 312162 360392 312200 360488
rect 437482 360392 437520 360488
rect 435312 359948 435350 360044
rect 560632 359948 560670 360044
rect 312162 359304 312200 359400
rect 437482 359304 437520 359400
rect 435312 358860 435350 358956
rect 560632 358860 560670 358956
rect 312162 358216 312200 358312
rect 437482 358216 437520 358312
rect 435312 357772 435350 357868
rect 560632 357772 560670 357868
rect 312162 357128 312200 357224
rect 437482 357128 437520 357224
rect 435312 356684 435350 356780
rect 560632 356684 560670 356780
rect 312162 356040 312200 356136
rect 437482 356040 437520 356136
rect 435312 355596 435350 355692
rect 560632 355596 560670 355692
rect 312162 354952 312200 355048
rect 437482 354952 437520 355048
rect 435312 354508 435350 354604
rect 560632 354508 560670 354604
rect 312162 353864 312200 353960
rect 437482 353864 437520 353960
rect 435312 353420 435350 353516
rect 560632 353420 560670 353516
rect 312162 352776 312200 352872
rect 437482 352776 437520 352872
rect 435312 352332 435350 352428
rect 560632 352332 560670 352428
rect 312162 351688 312200 351784
rect 437482 351688 437520 351784
rect 435312 351244 435350 351340
rect 560632 351244 560670 351340
rect 312162 350600 312200 350696
rect 437482 350600 437520 350696
rect 435312 350156 435350 350252
rect 560632 350156 560670 350252
rect 312162 349512 312200 349608
rect 437482 349512 437520 349608
rect 435312 349068 435350 349164
rect 560632 349068 560670 349164
rect 312162 348424 312200 348520
rect 437482 348424 437520 348520
rect 435312 347980 435350 348076
rect 560632 347980 560670 348076
rect 312162 347336 312200 347432
rect 437482 347336 437520 347432
rect 435312 346892 435350 346988
rect 560632 346892 560670 346988
rect 312162 346248 312200 346344
rect 437482 346248 437520 346344
rect 435312 345804 435350 345900
rect 560632 345804 560670 345900
rect 312162 345160 312200 345256
rect 437482 345160 437520 345256
rect 435312 344716 435350 344812
rect 560632 344716 560670 344812
rect 312162 344072 312200 344168
rect 437482 344072 437520 344168
rect 435312 343628 435350 343724
rect 560632 343628 560670 343724
rect 312162 342984 312200 343080
rect 437482 342984 437520 343080
rect 435312 342540 435350 342636
rect 560632 342540 560670 342636
rect 312162 341896 312200 341992
rect 437482 341896 437520 341992
rect 435312 341452 435350 341548
rect 560632 341452 560670 341548
rect 312162 340808 312200 340904
rect 437482 340808 437520 340904
rect 435312 340364 435350 340460
rect 560632 340364 560670 340460
rect 312162 339720 312200 339816
rect 437482 339720 437520 339816
rect 435312 339276 435350 339372
rect 560632 339276 560670 339372
rect 312162 338632 312200 338728
rect 437482 338632 437520 338728
rect 435312 338188 435350 338284
rect 560632 338188 560670 338284
rect 312162 337544 312200 337640
rect 437482 337544 437520 337640
rect 435312 337100 435350 337196
rect 560632 337100 560670 337196
rect 312162 336456 312200 336552
rect 437482 336456 437520 336552
rect 435312 336012 435350 336108
rect 560632 336012 560670 336108
rect 312162 335368 312200 335464
rect 437482 335368 437520 335464
rect 435312 334924 435350 335020
rect 560632 334924 560670 335020
rect 312162 334280 312200 334376
rect 437482 334280 437520 334376
rect 435312 333836 435350 333932
rect 560632 333836 560670 333932
rect 312162 333192 312200 333288
rect 437482 333192 437520 333288
rect 435312 332748 435350 332844
rect 560632 332748 560670 332844
rect 312162 332104 312200 332200
rect 437482 332104 437520 332200
rect 435312 331660 435350 331756
rect 560632 331660 560670 331756
rect 312162 331016 312200 331112
rect 437482 331016 437520 331112
rect 435312 330572 435350 330668
rect 560632 330572 560670 330668
rect 312162 329928 312200 330024
rect 437482 329928 437520 330024
rect 435312 329484 435350 329580
rect 560632 329484 560670 329580
rect 312162 328840 312200 328936
rect 437482 328840 437520 328936
rect 435312 328396 435350 328492
rect 560632 328396 560670 328492
rect 312162 327752 312200 327848
rect 437482 327752 437520 327848
rect 435312 327308 435350 327404
rect 560632 327308 560670 327404
rect 312162 326664 312200 326760
rect 437482 326664 437520 326760
rect 435312 326220 435350 326316
rect 560632 326220 560670 326316
rect 312162 325576 312200 325672
rect 437482 325576 437520 325672
rect 435312 325132 435350 325228
rect 560632 325132 560670 325228
rect 312162 324488 312200 324584
rect 437482 324488 437520 324584
rect 435312 324044 435350 324140
rect 560632 324044 560670 324140
rect 312162 323400 312200 323496
rect 437482 323400 437520 323496
rect 435312 322956 435350 323052
rect 560632 322956 560670 323052
rect 312162 322312 312200 322408
rect 437482 322312 437520 322408
rect 435312 321868 435350 321964
rect 560632 321868 560670 321964
rect 312162 321224 312200 321320
rect 437482 321224 437520 321320
rect 435312 320780 435350 320876
rect 560632 320780 560670 320876
rect 312162 320136 312200 320232
rect 437482 320136 437520 320232
rect 435312 319692 435350 319788
rect 560632 319692 560670 319788
rect 312162 319048 312200 319144
rect 437482 319048 437520 319144
rect 435312 318604 435350 318700
rect 560632 318604 560670 318700
rect 312162 317960 312200 318056
rect 437482 317960 437520 318056
rect 435312 317516 435350 317612
rect 560632 317516 560670 317612
rect 312162 316872 312200 316968
rect 437482 316872 437520 316968
rect 435312 316428 435350 316524
rect 560632 316428 560670 316524
rect 435312 315350 435350 315436
rect 560632 315350 560670 315436
rect 312162 310788 312200 310874
rect 437482 310788 437520 310874
rect 312162 309700 312200 309796
rect 437482 309700 437520 309796
rect 435312 309256 435350 309352
rect 560632 309256 560670 309352
rect 312162 308612 312200 308708
rect 437482 308612 437520 308708
rect 435312 308168 435350 308264
rect 560632 308168 560670 308264
rect 312162 307524 312200 307620
rect 437482 307524 437520 307620
rect 435312 307080 435350 307176
rect 560632 307080 560670 307176
rect 312162 306436 312200 306532
rect 437482 306436 437520 306532
rect 435312 305992 435350 306088
rect 560632 305992 560670 306088
rect 312162 305348 312200 305444
rect 437482 305348 437520 305444
rect 435312 304904 435350 305000
rect 560632 304904 560670 305000
rect 312162 304260 312200 304356
rect 437482 304260 437520 304356
rect 435312 303816 435350 303912
rect 560632 303816 560670 303912
rect 312162 303172 312200 303268
rect 437482 303172 437520 303268
rect 435312 302728 435350 302824
rect 560632 302728 560670 302824
rect 312162 302084 312200 302180
rect 437482 302084 437520 302180
rect 435312 301640 435350 301736
rect 560632 301640 560670 301736
rect 312162 300996 312200 301092
rect 437482 300996 437520 301092
rect 435312 300552 435350 300648
rect 560632 300552 560670 300648
rect 312162 299908 312200 300004
rect 437482 299908 437520 300004
rect 435312 299464 435350 299560
rect 560632 299464 560670 299560
rect 312162 298820 312200 298916
rect 437482 298820 437520 298916
rect 435312 298376 435350 298472
rect 560632 298376 560670 298472
rect 312162 297732 312200 297828
rect 437482 297732 437520 297828
rect 435312 297288 435350 297384
rect 560632 297288 560670 297384
rect 312162 296644 312200 296740
rect 437482 296644 437520 296740
rect 435312 296200 435350 296296
rect 560632 296200 560670 296296
rect 312162 295556 312200 295652
rect 437482 295556 437520 295652
rect 435312 295112 435350 295208
rect 560632 295112 560670 295208
rect 312162 294468 312200 294564
rect 437482 294468 437520 294564
rect 435312 294024 435350 294120
rect 560632 294024 560670 294120
rect 312162 293380 312200 293476
rect 437482 293380 437520 293476
rect 435312 292936 435350 293032
rect 560632 292936 560670 293032
rect 312162 292292 312200 292388
rect 437482 292292 437520 292388
rect 435312 291848 435350 291944
rect 560632 291848 560670 291944
rect 312162 291204 312200 291300
rect 437482 291204 437520 291300
rect 435312 290760 435350 290856
rect 560632 290760 560670 290856
rect 312162 290116 312200 290212
rect 437482 290116 437520 290212
rect 435312 289672 435350 289768
rect 560632 289672 560670 289768
rect 312162 289028 312200 289124
rect 437482 289028 437520 289124
rect 435312 288584 435350 288680
rect 560632 288584 560670 288680
rect 312162 287940 312200 288036
rect 437482 287940 437520 288036
rect 435312 287496 435350 287592
rect 560632 287496 560670 287592
rect 312162 286852 312200 286948
rect 437482 286852 437520 286948
rect 435312 286408 435350 286504
rect 560632 286408 560670 286504
rect 312162 285764 312200 285860
rect 437482 285764 437520 285860
rect 435312 285320 435350 285416
rect 560632 285320 560670 285416
rect 312162 284676 312200 284772
rect 437482 284676 437520 284772
rect 435312 284232 435350 284328
rect 560632 284232 560670 284328
rect 312162 283588 312200 283684
rect 437482 283588 437520 283684
rect 435312 283144 435350 283240
rect 560632 283144 560670 283240
rect 312162 282500 312200 282596
rect 437482 282500 437520 282596
rect 435312 282056 435350 282152
rect 560632 282056 560670 282152
rect 312162 281412 312200 281508
rect 437482 281412 437520 281508
rect 435312 280968 435350 281064
rect 560632 280968 560670 281064
rect 312162 280324 312200 280420
rect 437482 280324 437520 280420
rect 435312 279880 435350 279976
rect 560632 279880 560670 279976
rect 312162 279236 312200 279332
rect 437482 279236 437520 279332
rect 435312 278792 435350 278888
rect 560632 278792 560670 278888
rect 312162 278148 312200 278244
rect 437482 278148 437520 278244
rect 435312 277704 435350 277800
rect 560632 277704 560670 277800
rect 312162 277060 312200 277156
rect 437482 277060 437520 277156
rect 435312 276616 435350 276712
rect 560632 276616 560670 276712
rect 312162 275972 312200 276068
rect 437482 275972 437520 276068
rect 435312 275528 435350 275624
rect 560632 275528 560670 275624
rect 312162 274884 312200 274980
rect 437482 274884 437520 274980
rect 435312 274440 435350 274536
rect 560632 274440 560670 274536
rect 312162 273796 312200 273892
rect 437482 273796 437520 273892
rect 435312 273352 435350 273448
rect 560632 273352 560670 273448
rect 312162 272708 312200 272804
rect 437482 272708 437520 272804
rect 435312 272264 435350 272360
rect 560632 272264 560670 272360
rect 312162 271620 312200 271716
rect 437482 271620 437520 271716
rect 435312 271176 435350 271272
rect 560632 271176 560670 271272
rect 312162 270532 312200 270628
rect 437482 270532 437520 270628
rect 435312 270088 435350 270184
rect 560632 270088 560670 270184
rect 312162 269444 312200 269540
rect 437482 269444 437520 269540
rect 435312 269000 435350 269096
rect 560632 269000 560670 269096
rect 312162 268356 312200 268452
rect 437482 268356 437520 268452
rect 435312 267912 435350 268008
rect 560632 267912 560670 268008
rect 312162 267268 312200 267364
rect 437482 267268 437520 267364
rect 435312 266824 435350 266920
rect 560632 266824 560670 266920
rect 312162 266180 312200 266276
rect 437482 266180 437520 266276
rect 435312 265736 435350 265832
rect 560632 265736 560670 265832
rect 312162 265092 312200 265188
rect 437482 265092 437520 265188
rect 435312 264648 435350 264744
rect 560632 264648 560670 264744
rect 312162 264004 312200 264100
rect 437482 264004 437520 264100
rect 435312 263560 435350 263656
rect 560632 263560 560670 263656
rect 312162 262916 312200 263012
rect 437482 262916 437520 263012
rect 435312 262472 435350 262568
rect 560632 262472 560670 262568
rect 312162 261828 312200 261924
rect 437482 261828 437520 261924
rect 435312 261384 435350 261480
rect 560632 261384 560670 261480
rect 312162 260740 312200 260836
rect 437482 260740 437520 260836
rect 435312 260296 435350 260392
rect 560632 260296 560670 260392
rect 312162 259652 312200 259748
rect 437482 259652 437520 259748
rect 435312 259208 435350 259304
rect 560632 259208 560670 259304
rect 312162 258564 312200 258660
rect 437482 258564 437520 258660
rect 435312 258120 435350 258216
rect 560632 258120 560670 258216
rect 312162 257476 312200 257572
rect 437482 257476 437520 257572
rect 435312 257032 435350 257128
rect 560632 257032 560670 257128
rect 312162 256388 312200 256484
rect 437482 256388 437520 256484
rect 435312 255944 435350 256040
rect 560632 255944 560670 256040
rect 312162 255300 312200 255396
rect 437482 255300 437520 255396
rect 435312 254856 435350 254952
rect 560632 254856 560670 254952
rect 312162 254212 312200 254308
rect 437482 254212 437520 254308
rect 435312 253768 435350 253864
rect 560632 253768 560670 253864
rect 435312 252690 435350 252776
rect 560632 252690 560670 252776
rect 312162 248128 312200 248214
rect 437482 248128 437520 248214
rect 312162 247040 312200 247136
rect 437482 247040 437520 247136
rect 435312 246596 435350 246692
rect 560632 246596 560670 246692
rect 312162 245952 312200 246048
rect 437482 245952 437520 246048
rect 435312 245508 435350 245604
rect 560632 245508 560670 245604
rect 312162 244864 312200 244960
rect 437482 244864 437520 244960
rect 435312 244420 435350 244516
rect 560632 244420 560670 244516
rect 312162 243776 312200 243872
rect 437482 243776 437520 243872
rect 435312 243332 435350 243428
rect 560632 243332 560670 243428
rect 312162 242688 312200 242784
rect 437482 242688 437520 242784
rect 435312 242244 435350 242340
rect 560632 242244 560670 242340
rect 312162 241600 312200 241696
rect 437482 241600 437520 241696
rect 435312 241156 435350 241252
rect 560632 241156 560670 241252
rect 312162 240512 312200 240608
rect 437482 240512 437520 240608
rect 435312 240068 435350 240164
rect 560632 240068 560670 240164
rect 312162 239424 312200 239520
rect 437482 239424 437520 239520
rect 435312 238980 435350 239076
rect 560632 238980 560670 239076
rect 312162 238336 312200 238432
rect 437482 238336 437520 238432
rect 435312 237892 435350 237988
rect 560632 237892 560670 237988
rect 312162 237248 312200 237344
rect 437482 237248 437520 237344
rect 435312 236804 435350 236900
rect 560632 236804 560670 236900
rect 312162 236160 312200 236256
rect 437482 236160 437520 236256
rect 435312 235716 435350 235812
rect 560632 235716 560670 235812
rect 312162 235072 312200 235168
rect 437482 235072 437520 235168
rect 435312 234628 435350 234724
rect 560632 234628 560670 234724
rect 312162 233984 312200 234080
rect 437482 233984 437520 234080
rect 435312 233540 435350 233636
rect 560632 233540 560670 233636
rect 312162 232896 312200 232992
rect 437482 232896 437520 232992
rect 435312 232452 435350 232548
rect 560632 232452 560670 232548
rect 312162 231808 312200 231904
rect 437482 231808 437520 231904
rect 435312 231364 435350 231460
rect 560632 231364 560670 231460
rect 312162 230720 312200 230816
rect 437482 230720 437520 230816
rect 435312 230276 435350 230372
rect 560632 230276 560670 230372
rect 312162 229632 312200 229728
rect 437482 229632 437520 229728
rect 435312 229188 435350 229284
rect 560632 229188 560670 229284
rect 312162 228544 312200 228640
rect 437482 228544 437520 228640
rect 435312 228100 435350 228196
rect 560632 228100 560670 228196
rect 312162 227456 312200 227552
rect 437482 227456 437520 227552
rect 435312 227012 435350 227108
rect 560632 227012 560670 227108
rect 312162 226368 312200 226464
rect 437482 226368 437520 226464
rect 435312 225924 435350 226020
rect 560632 225924 560670 226020
rect 312162 225280 312200 225376
rect 437482 225280 437520 225376
rect 435312 224836 435350 224932
rect 560632 224836 560670 224932
rect 312162 224192 312200 224288
rect 437482 224192 437520 224288
rect 435312 223748 435350 223844
rect 560632 223748 560670 223844
rect 312162 223104 312200 223200
rect 437482 223104 437520 223200
rect 435312 222660 435350 222756
rect 560632 222660 560670 222756
rect 312162 222016 312200 222112
rect 437482 222016 437520 222112
rect 435312 221572 435350 221668
rect 560632 221572 560670 221668
rect 312162 220928 312200 221024
rect 437482 220928 437520 221024
rect 435312 220484 435350 220580
rect 560632 220484 560670 220580
rect 312162 219840 312200 219936
rect 437482 219840 437520 219936
rect 435312 219396 435350 219492
rect 560632 219396 560670 219492
rect 312162 218752 312200 218848
rect 437482 218752 437520 218848
rect 435312 218308 435350 218404
rect 560632 218308 560670 218404
rect 312162 217664 312200 217760
rect 437482 217664 437520 217760
rect 435312 217220 435350 217316
rect 560632 217220 560670 217316
rect 312162 216576 312200 216672
rect 437482 216576 437520 216672
rect 435312 216132 435350 216228
rect 560632 216132 560670 216228
rect 312162 215488 312200 215584
rect 437482 215488 437520 215584
rect 435312 215044 435350 215140
rect 560632 215044 560670 215140
rect 312162 214400 312200 214496
rect 437482 214400 437520 214496
rect 435312 213956 435350 214052
rect 560632 213956 560670 214052
rect 312162 213312 312200 213408
rect 437482 213312 437520 213408
rect 435312 212868 435350 212964
rect 560632 212868 560670 212964
rect 312162 212224 312200 212320
rect 437482 212224 437520 212320
rect 435312 211780 435350 211876
rect 560632 211780 560670 211876
rect 312162 211136 312200 211232
rect 437482 211136 437520 211232
rect 435312 210692 435350 210788
rect 560632 210692 560670 210788
rect 312162 210048 312200 210144
rect 437482 210048 437520 210144
rect 435312 209604 435350 209700
rect 560632 209604 560670 209700
rect 312162 208960 312200 209056
rect 437482 208960 437520 209056
rect 435312 208516 435350 208612
rect 560632 208516 560670 208612
rect 312162 207872 312200 207968
rect 437482 207872 437520 207968
rect 435312 207428 435350 207524
rect 560632 207428 560670 207524
rect 312162 206784 312200 206880
rect 437482 206784 437520 206880
rect 435312 206340 435350 206436
rect 560632 206340 560670 206436
rect 312162 205696 312200 205792
rect 437482 205696 437520 205792
rect 435312 205252 435350 205348
rect 560632 205252 560670 205348
rect 312162 204608 312200 204704
rect 437482 204608 437520 204704
rect 435312 204164 435350 204260
rect 560632 204164 560670 204260
rect 312162 203520 312200 203616
rect 437482 203520 437520 203616
rect 435312 203076 435350 203172
rect 560632 203076 560670 203172
rect 312162 202432 312200 202528
rect 437482 202432 437520 202528
rect 435312 201988 435350 202084
rect 560632 201988 560670 202084
rect 312162 201344 312200 201440
rect 437482 201344 437520 201440
rect 435312 200900 435350 200996
rect 560632 200900 560670 200996
rect 312162 200256 312200 200352
rect 437482 200256 437520 200352
rect 435312 199812 435350 199908
rect 560632 199812 560670 199908
rect 312162 199168 312200 199264
rect 437482 199168 437520 199264
rect 435312 198724 435350 198820
rect 560632 198724 560670 198820
rect 312162 198080 312200 198176
rect 437482 198080 437520 198176
rect 435312 197636 435350 197732
rect 560632 197636 560670 197732
rect 312162 196992 312200 197088
rect 437482 196992 437520 197088
rect 435312 196548 435350 196644
rect 560632 196548 560670 196644
rect 312162 195904 312200 196000
rect 437482 195904 437520 196000
rect 435312 195460 435350 195556
rect 560632 195460 560670 195556
rect 312162 194816 312200 194912
rect 437482 194816 437520 194912
rect 435312 194372 435350 194468
rect 560632 194372 560670 194468
rect 312162 193728 312200 193824
rect 437482 193728 437520 193824
rect 435312 193284 435350 193380
rect 560632 193284 560670 193380
rect 312162 192640 312200 192736
rect 437482 192640 437520 192736
rect 435312 192196 435350 192292
rect 560632 192196 560670 192292
rect 312162 191552 312200 191648
rect 437482 191552 437520 191648
rect 435312 191108 435350 191204
rect 560632 191108 560670 191204
rect 435312 190030 435350 190116
rect 560632 190030 560670 190116
rect 312162 185468 312200 185554
rect 437482 185468 437520 185554
rect 312162 184380 312200 184476
rect 437482 184380 437520 184476
rect 435312 183936 435350 184032
rect 560632 183936 560670 184032
rect 312162 183292 312200 183388
rect 437482 183292 437520 183388
rect 435312 182848 435350 182944
rect 560632 182848 560670 182944
rect 312162 182204 312200 182300
rect 437482 182204 437520 182300
rect 435312 181760 435350 181856
rect 560632 181760 560670 181856
rect 312162 181116 312200 181212
rect 437482 181116 437520 181212
rect 435312 180672 435350 180768
rect 560632 180672 560670 180768
rect 312162 180028 312200 180124
rect 437482 180028 437520 180124
rect 435312 179584 435350 179680
rect 560632 179584 560670 179680
rect 312162 178940 312200 179036
rect 437482 178940 437520 179036
rect 435312 178496 435350 178592
rect 560632 178496 560670 178592
rect 312162 177852 312200 177948
rect 437482 177852 437520 177948
rect 435312 177408 435350 177504
rect 560632 177408 560670 177504
rect 312162 176764 312200 176860
rect 437482 176764 437520 176860
rect 435312 176320 435350 176416
rect 560632 176320 560670 176416
rect 312162 175676 312200 175772
rect 437482 175676 437520 175772
rect 435312 175232 435350 175328
rect 560632 175232 560670 175328
rect 312162 174588 312200 174684
rect 437482 174588 437520 174684
rect 435312 174144 435350 174240
rect 560632 174144 560670 174240
rect 312162 173500 312200 173596
rect 437482 173500 437520 173596
rect 435312 173056 435350 173152
rect 560632 173056 560670 173152
rect 312162 172412 312200 172508
rect 437482 172412 437520 172508
rect 435312 171968 435350 172064
rect 560632 171968 560670 172064
rect 312162 171324 312200 171420
rect 437482 171324 437520 171420
rect 435312 170880 435350 170976
rect 560632 170880 560670 170976
rect 312162 170236 312200 170332
rect 437482 170236 437520 170332
rect 435312 169792 435350 169888
rect 560632 169792 560670 169888
rect 312162 169148 312200 169244
rect 437482 169148 437520 169244
rect 435312 168704 435350 168800
rect 560632 168704 560670 168800
rect 312162 168060 312200 168156
rect 437482 168060 437520 168156
rect 435312 167616 435350 167712
rect 560632 167616 560670 167712
rect 312162 166972 312200 167068
rect 437482 166972 437520 167068
rect 435312 166528 435350 166624
rect 560632 166528 560670 166624
rect 312162 165884 312200 165980
rect 437482 165884 437520 165980
rect 435312 165440 435350 165536
rect 560632 165440 560670 165536
rect 312162 164796 312200 164892
rect 437482 164796 437520 164892
rect 435312 164352 435350 164448
rect 560632 164352 560670 164448
rect 312162 163708 312200 163804
rect 437482 163708 437520 163804
rect 435312 163264 435350 163360
rect 560632 163264 560670 163360
rect 312162 162620 312200 162716
rect 437482 162620 437520 162716
rect 435312 162176 435350 162272
rect 560632 162176 560670 162272
rect 312162 161532 312200 161628
rect 437482 161532 437520 161628
rect 435312 161088 435350 161184
rect 560632 161088 560670 161184
rect 312162 160444 312200 160540
rect 437482 160444 437520 160540
rect 435312 160000 435350 160096
rect 560632 160000 560670 160096
rect 312162 159356 312200 159452
rect 437482 159356 437520 159452
rect 435312 158912 435350 159008
rect 560632 158912 560670 159008
rect 312162 158268 312200 158364
rect 437482 158268 437520 158364
rect 435312 157824 435350 157920
rect 560632 157824 560670 157920
rect 312162 157180 312200 157276
rect 437482 157180 437520 157276
rect 435312 156736 435350 156832
rect 560632 156736 560670 156832
rect 312162 156092 312200 156188
rect 437482 156092 437520 156188
rect 435312 155648 435350 155744
rect 560632 155648 560670 155744
rect 312162 155004 312200 155100
rect 437482 155004 437520 155100
rect 435312 154560 435350 154656
rect 560632 154560 560670 154656
rect 312162 153916 312200 154012
rect 437482 153916 437520 154012
rect 435312 153472 435350 153568
rect 560632 153472 560670 153568
rect 312162 152828 312200 152924
rect 437482 152828 437520 152924
rect 435312 152384 435350 152480
rect 560632 152384 560670 152480
rect 312162 151740 312200 151836
rect 437482 151740 437520 151836
rect 435312 151296 435350 151392
rect 560632 151296 560670 151392
rect 312162 150652 312200 150748
rect 437482 150652 437520 150748
rect 435312 150208 435350 150304
rect 560632 150208 560670 150304
rect 312162 149564 312200 149660
rect 437482 149564 437520 149660
rect 435312 149120 435350 149216
rect 560632 149120 560670 149216
rect 312162 148476 312200 148572
rect 437482 148476 437520 148572
rect 435312 148032 435350 148128
rect 560632 148032 560670 148128
rect 312162 147388 312200 147484
rect 437482 147388 437520 147484
rect 435312 146944 435350 147040
rect 560632 146944 560670 147040
rect 312162 146300 312200 146396
rect 437482 146300 437520 146396
rect 435312 145856 435350 145952
rect 560632 145856 560670 145952
rect 312162 145212 312200 145308
rect 437482 145212 437520 145308
rect 435312 144768 435350 144864
rect 560632 144768 560670 144864
rect 312162 144124 312200 144220
rect 437482 144124 437520 144220
rect 435312 143680 435350 143776
rect 560632 143680 560670 143776
rect 312162 143036 312200 143132
rect 437482 143036 437520 143132
rect 435312 142592 435350 142688
rect 560632 142592 560670 142688
rect 312162 141948 312200 142044
rect 437482 141948 437520 142044
rect 435312 141504 435350 141600
rect 560632 141504 560670 141600
rect 312162 140860 312200 140956
rect 437482 140860 437520 140956
rect 435312 140416 435350 140512
rect 560632 140416 560670 140512
rect 312162 139772 312200 139868
rect 437482 139772 437520 139868
rect 435312 139328 435350 139424
rect 560632 139328 560670 139424
rect 312162 138684 312200 138780
rect 437482 138684 437520 138780
rect 435312 138240 435350 138336
rect 560632 138240 560670 138336
rect 312162 137596 312200 137692
rect 437482 137596 437520 137692
rect 435312 137152 435350 137248
rect 560632 137152 560670 137248
rect 312162 136508 312200 136604
rect 437482 136508 437520 136604
rect 435312 136064 435350 136160
rect 560632 136064 560670 136160
rect 312162 135420 312200 135516
rect 437482 135420 437520 135516
rect 435312 134976 435350 135072
rect 560632 134976 560670 135072
rect 312162 134332 312200 134428
rect 437482 134332 437520 134428
rect 435312 133888 435350 133984
rect 560632 133888 560670 133984
rect 312162 133244 312200 133340
rect 437482 133244 437520 133340
rect 435312 132800 435350 132896
rect 560632 132800 560670 132896
rect 312162 132156 312200 132252
rect 437482 132156 437520 132252
rect 435312 131712 435350 131808
rect 560632 131712 560670 131808
rect 312162 131068 312200 131164
rect 437482 131068 437520 131164
rect 435312 130624 435350 130720
rect 560632 130624 560670 130720
rect 312162 129980 312200 130076
rect 437482 129980 437520 130076
rect 435312 129536 435350 129632
rect 560632 129536 560670 129632
rect 312162 128892 312200 128988
rect 437482 128892 437520 128988
rect 435312 128448 435350 128544
rect 560632 128448 560670 128544
rect 435312 127370 435350 127456
rect 560632 127370 560670 127456
rect 312162 122808 312200 122894
rect 437482 122808 437520 122894
rect 312162 121720 312200 121816
rect 437482 121720 437520 121816
rect 435312 121276 435350 121372
rect 560632 121276 560670 121372
rect 312162 120632 312200 120728
rect 437482 120632 437520 120728
rect 435312 120188 435350 120284
rect 560632 120188 560670 120284
rect 312162 119544 312200 119640
rect 437482 119544 437520 119640
rect 435312 119100 435350 119196
rect 560632 119100 560670 119196
rect 312162 118456 312200 118552
rect 437482 118456 437520 118552
rect 435312 118012 435350 118108
rect 560632 118012 560670 118108
rect 312162 117368 312200 117464
rect 437482 117368 437520 117464
rect 435312 116924 435350 117020
rect 560632 116924 560670 117020
rect 312162 116280 312200 116376
rect 437482 116280 437520 116376
rect 435312 115836 435350 115932
rect 560632 115836 560670 115932
rect 312162 115192 312200 115288
rect 437482 115192 437520 115288
rect 435312 114748 435350 114844
rect 560632 114748 560670 114844
rect 312162 114104 312200 114200
rect 437482 114104 437520 114200
rect 435312 113660 435350 113756
rect 560632 113660 560670 113756
rect 312162 113016 312200 113112
rect 437482 113016 437520 113112
rect 435312 112572 435350 112668
rect 560632 112572 560670 112668
rect 312162 111928 312200 112024
rect 437482 111928 437520 112024
rect 435312 111484 435350 111580
rect 560632 111484 560670 111580
rect 312162 110840 312200 110936
rect 437482 110840 437520 110936
rect 435312 110396 435350 110492
rect 560632 110396 560670 110492
rect 312162 109752 312200 109848
rect 437482 109752 437520 109848
rect 435312 109308 435350 109404
rect 560632 109308 560670 109404
rect 312162 108664 312200 108760
rect 437482 108664 437520 108760
rect 435312 108220 435350 108316
rect 560632 108220 560670 108316
rect 312162 107576 312200 107672
rect 437482 107576 437520 107672
rect 435312 107132 435350 107228
rect 560632 107132 560670 107228
rect 312162 106488 312200 106584
rect 437482 106488 437520 106584
rect 435312 106044 435350 106140
rect 560632 106044 560670 106140
rect 312162 105400 312200 105496
rect 437482 105400 437520 105496
rect 435312 104956 435350 105052
rect 560632 104956 560670 105052
rect 312162 104312 312200 104408
rect 437482 104312 437520 104408
rect 435312 103868 435350 103964
rect 560632 103868 560670 103964
rect 312162 103224 312200 103320
rect 437482 103224 437520 103320
rect 435312 102780 435350 102876
rect 560632 102780 560670 102876
rect 312162 102136 312200 102232
rect 437482 102136 437520 102232
rect 435312 101692 435350 101788
rect 560632 101692 560670 101788
rect 312162 101048 312200 101144
rect 437482 101048 437520 101144
rect 435312 100604 435350 100700
rect 560632 100604 560670 100700
rect 312162 99960 312200 100056
rect 437482 99960 437520 100056
rect 435312 99516 435350 99612
rect 560632 99516 560670 99612
rect 312162 98872 312200 98968
rect 437482 98872 437520 98968
rect 435312 98428 435350 98524
rect 560632 98428 560670 98524
rect 312162 97784 312200 97880
rect 437482 97784 437520 97880
rect 435312 97340 435350 97436
rect 560632 97340 560670 97436
rect 312162 96696 312200 96792
rect 437482 96696 437520 96792
rect 435312 96252 435350 96348
rect 560632 96252 560670 96348
rect 312162 95608 312200 95704
rect 437482 95608 437520 95704
rect 435312 95164 435350 95260
rect 560632 95164 560670 95260
rect 312162 94520 312200 94616
rect 437482 94520 437520 94616
rect 435312 94076 435350 94172
rect 560632 94076 560670 94172
rect 312162 93432 312200 93528
rect 437482 93432 437520 93528
rect 435312 92988 435350 93084
rect 560632 92988 560670 93084
rect 312162 92344 312200 92440
rect 437482 92344 437520 92440
rect 435312 91900 435350 91996
rect 560632 91900 560670 91996
rect 312162 91256 312200 91352
rect 437482 91256 437520 91352
rect 435312 90812 435350 90908
rect 560632 90812 560670 90908
rect 312162 90168 312200 90264
rect 437482 90168 437520 90264
rect 435312 89724 435350 89820
rect 560632 89724 560670 89820
rect 312162 89080 312200 89176
rect 437482 89080 437520 89176
rect 435312 88636 435350 88732
rect 560632 88636 560670 88732
rect 312162 87992 312200 88088
rect 437482 87992 437520 88088
rect 435312 87548 435350 87644
rect 560632 87548 560670 87644
rect 312162 86904 312200 87000
rect 437482 86904 437520 87000
rect 435312 86460 435350 86556
rect 560632 86460 560670 86556
rect 312162 85816 312200 85912
rect 437482 85816 437520 85912
rect 435312 85372 435350 85468
rect 560632 85372 560670 85468
rect 312162 84728 312200 84824
rect 437482 84728 437520 84824
rect 435312 84284 435350 84380
rect 560632 84284 560670 84380
rect 312162 83640 312200 83736
rect 437482 83640 437520 83736
rect 435312 83196 435350 83292
rect 560632 83196 560670 83292
rect 312162 82552 312200 82648
rect 437482 82552 437520 82648
rect 435312 82108 435350 82204
rect 560632 82108 560670 82204
rect 312162 81464 312200 81560
rect 437482 81464 437520 81560
rect 435312 81020 435350 81116
rect 560632 81020 560670 81116
rect 312162 80376 312200 80472
rect 437482 80376 437520 80472
rect 435312 79932 435350 80028
rect 560632 79932 560670 80028
rect 312162 79288 312200 79384
rect 437482 79288 437520 79384
rect 435312 78844 435350 78940
rect 560632 78844 560670 78940
rect 312162 78200 312200 78296
rect 437482 78200 437520 78296
rect 435312 77756 435350 77852
rect 560632 77756 560670 77852
rect 312162 77112 312200 77208
rect 437482 77112 437520 77208
rect 435312 76668 435350 76764
rect 560632 76668 560670 76764
rect 312162 76024 312200 76120
rect 437482 76024 437520 76120
rect 435312 75580 435350 75676
rect 560632 75580 560670 75676
rect 312162 74936 312200 75032
rect 437482 74936 437520 75032
rect 435312 74492 435350 74588
rect 560632 74492 560670 74588
rect 312162 73848 312200 73944
rect 437482 73848 437520 73944
rect 435312 73404 435350 73500
rect 560632 73404 560670 73500
rect 312162 72760 312200 72856
rect 437482 72760 437520 72856
rect 435312 72316 435350 72412
rect 560632 72316 560670 72412
rect 312162 71672 312200 71768
rect 437482 71672 437520 71768
rect 435312 71228 435350 71324
rect 560632 71228 560670 71324
rect 312162 70584 312200 70680
rect 437482 70584 437520 70680
rect 435312 70140 435350 70236
rect 560632 70140 560670 70236
rect 312162 69496 312200 69592
rect 437482 69496 437520 69592
rect 435312 69052 435350 69148
rect 560632 69052 560670 69148
rect 312162 68408 312200 68504
rect 437482 68408 437520 68504
rect 435312 67964 435350 68060
rect 560632 67964 560670 68060
rect 312162 67320 312200 67416
rect 437482 67320 437520 67416
rect 435312 66876 435350 66972
rect 560632 66876 560670 66972
rect 312162 66232 312200 66328
rect 437482 66232 437520 66328
rect 435312 65788 435350 65884
rect 560632 65788 560670 65884
rect 435312 64710 435350 64796
rect 560632 64710 560670 64796
<< pwell >>
rect 123720 642790 131790 643240
rect 123620 642690 131790 642790
rect 123720 641500 131790 642690
rect 127380 641490 128420 641500
rect 127860 641170 127960 641210
rect 123710 634960 129470 637430
rect 124030 630260 129710 630990
rect 124000 630000 129710 630260
rect 124030 629310 129710 630000
rect 124280 623960 129360 624470
rect 124260 623740 129360 623960
rect 124250 623480 129360 623740
rect 124280 622790 129360 623480
rect 125040 618990 132070 619080
rect 125040 618120 132080 618990
rect 125040 618060 125370 618120
rect 125730 618060 125870 618120
rect 126230 618060 126370 618120
rect 126730 618060 126870 618120
rect 127230 618060 127370 618120
rect 127730 618060 127870 618120
rect 128230 618060 129020 618120
rect 129230 618060 129370 618120
rect 129730 618060 129870 618120
rect 129950 617520 130390 618120
rect 130730 618060 130870 618120
rect 131230 618060 131370 618120
rect 131730 618060 131870 618120
rect 131940 618060 132080 618120
rect 124690 611540 131720 611630
rect 124690 610670 131730 611540
rect 124690 610610 125020 610670
rect 125380 610610 125520 610670
rect 125880 610610 126020 610670
rect 126380 610610 126520 610670
rect 126880 610610 127020 610670
rect 127380 610610 127520 610670
rect 127880 610610 128670 610670
rect 128880 610610 129020 610670
rect 129380 610610 129520 610670
rect 129600 610070 130040 610670
rect 130380 610610 130520 610670
rect 130880 610610 131020 610670
rect 131380 610610 131520 610670
rect 131590 610610 131730 610670
rect 124820 605490 131850 605580
rect 124820 604520 131860 605490
rect 124820 604460 125150 604520
rect 125510 604460 125650 604520
rect 126010 604460 126150 604520
rect 126510 604460 126650 604520
rect 127010 604460 127150 604520
rect 127510 604460 127650 604520
rect 128010 604460 128800 604520
rect 129010 604460 129150 604520
rect 129510 604460 129650 604520
rect 129730 603920 130170 604520
rect 130510 604460 130650 604520
rect 131010 604460 131150 604520
rect 131510 604460 131650 604520
rect 131720 604460 131860 604520
rect 124620 599230 131650 599320
rect 124620 598160 131660 599230
rect 124620 598100 124950 598160
rect 125310 598100 125450 598160
rect 125810 598100 125950 598160
rect 126310 598100 126450 598160
rect 126810 598100 126950 598160
rect 127310 598100 127450 598160
rect 127810 598100 128600 598160
rect 128810 598100 128950 598160
rect 129310 598100 129450 598160
rect 129530 597560 129970 598160
rect 130310 598100 130450 598160
rect 130810 598100 130950 598160
rect 131310 598100 131450 598160
rect 131520 598100 131660 598160
rect 124580 591680 131610 591770
rect 124580 590510 131620 591680
rect 124580 590450 124910 590510
rect 125270 590450 125410 590510
rect 125770 590450 125910 590510
rect 126270 590450 126410 590510
rect 126770 590450 126910 590510
rect 127270 590450 127410 590510
rect 127770 590450 128560 590510
rect 128770 590450 128910 590510
rect 129270 590450 129410 590510
rect 129490 589910 129930 590510
rect 130270 590450 130410 590510
rect 130770 590450 130910 590510
rect 131270 590450 131410 590510
rect 131480 590450 131620 590510
rect 124880 581620 133080 582830
rect 124920 572500 133120 573810
rect 124870 564730 133070 566140
rect 124870 558090 133070 559600
rect 124940 551560 134090 552770
rect 124940 543790 134090 545200
rect 124910 535530 134060 537140
<< nmos >>
rect 124150 642310 124240 642340
rect 124330 642310 124420 642340
rect 124510 642310 124600 642340
rect 124690 642310 124780 642340
rect 124870 642310 124960 642340
rect 125050 642310 125140 642340
rect 125230 642310 125320 642340
rect 125410 642310 125500 642340
rect 125590 642310 125680 642340
rect 125770 642310 125860 642340
rect 125950 642310 126040 642340
rect 126130 642310 126220 642340
rect 126310 642310 126400 642340
rect 126490 642310 126580 642340
rect 126670 642310 126760 642340
rect 126850 642310 126940 642340
rect 127030 642310 127120 642340
rect 127210 642310 127300 642340
rect 127390 642310 127480 642340
rect 127570 642310 127660 642340
rect 127750 642310 127840 642340
rect 127930 642310 128020 642340
rect 128110 642310 128200 642340
rect 128290 642310 128380 642340
rect 128470 642310 128560 642340
rect 128650 642310 128740 642340
rect 128830 642310 128920 642340
rect 129010 642310 129100 642340
rect 129190 642310 129280 642340
rect 129370 642310 129460 642340
rect 129550 642310 129640 642340
rect 129730 642310 129820 642340
rect 129910 642310 130000 642340
rect 130090 642310 130180 642340
rect 130270 642310 130360 642340
rect 130450 642310 130540 642340
rect 130630 642310 130720 642340
rect 130810 642310 130900 642340
rect 130990 642310 131080 642340
rect 131170 642310 131260 642340
rect 124180 636140 124360 636170
rect 124420 636140 124600 636170
rect 124660 636140 124840 636170
rect 124900 636140 125080 636170
rect 125140 636140 125320 636170
rect 125380 636140 125560 636170
rect 125620 636140 125800 636170
rect 125860 636140 126040 636170
rect 126100 636140 126280 636170
rect 126340 636140 126520 636170
rect 126580 636140 126760 636170
rect 126820 636140 127000 636170
rect 127060 636140 127240 636170
rect 127300 636140 127480 636170
rect 127540 636140 127720 636170
rect 127780 636140 127960 636170
rect 128020 636140 128200 636170
rect 128260 636140 128440 636170
rect 128500 636140 128680 636170
rect 128740 636140 128920 636170
rect 124240 632550 124640 632580
rect 124450 630110 124850 630140
rect 124910 630110 125310 630140
rect 125370 630110 125770 630140
rect 125830 630110 126230 630140
rect 126290 630110 126690 630140
rect 126750 630110 127150 630140
rect 127210 630110 127610 630140
rect 127670 630110 128070 630140
rect 128130 630110 128530 630140
rect 128590 630110 128990 630140
rect 124220 624880 124820 624910
rect 124780 623590 125380 623620
rect 125440 623590 126040 623620
rect 126100 623590 126700 623620
rect 126760 623590 127360 623620
rect 127420 623590 128020 623620
rect 128080 623590 128680 623620
rect 125530 619400 125560 619450
rect 125420 619370 125560 619400
rect 125420 619290 125450 619370
rect 125530 619290 125560 619370
rect 125420 619260 125560 619290
rect 125600 618620 125630 618670
rect 125490 618590 125630 618620
rect 125490 618510 125520 618590
rect 125600 618510 125630 618590
rect 125490 618480 125630 618510
rect 125940 618620 125970 618670
rect 125830 618590 125970 618620
rect 125830 618510 125860 618590
rect 125940 618510 125970 618590
rect 125830 618480 125970 618510
rect 126280 618620 126310 618670
rect 126170 618590 126310 618620
rect 126170 618510 126200 618590
rect 126280 618510 126310 618590
rect 126170 618480 126310 618510
rect 126620 618620 126650 618670
rect 126510 618590 126650 618620
rect 126510 618510 126540 618590
rect 126620 618510 126650 618590
rect 126510 618480 126650 618510
rect 126960 618620 126990 618670
rect 126850 618590 126990 618620
rect 126850 618510 126880 618590
rect 126960 618510 126990 618590
rect 126850 618480 126990 618510
rect 127300 618620 127330 618670
rect 127190 618590 127330 618620
rect 127190 618510 127220 618590
rect 127300 618510 127330 618590
rect 127190 618480 127330 618510
rect 127640 618620 127670 618670
rect 127530 618590 127670 618620
rect 127530 618510 127560 618590
rect 127640 618510 127670 618590
rect 127530 618480 127670 618510
rect 127980 618620 128010 618670
rect 127870 618590 128010 618620
rect 127870 618510 127900 618590
rect 127980 618510 128010 618590
rect 127870 618480 128010 618510
rect 128320 618620 128350 618670
rect 128210 618590 128350 618620
rect 128210 618510 128240 618590
rect 128320 618510 128350 618590
rect 128210 618480 128350 618510
rect 128660 618620 128690 618670
rect 128550 618590 128690 618620
rect 128550 618510 128580 618590
rect 128660 618510 128690 618590
rect 128550 618480 128690 618510
rect 129000 618620 129030 618670
rect 128890 618590 129030 618620
rect 128890 618510 128920 618590
rect 129000 618510 129030 618590
rect 128890 618480 129030 618510
rect 129340 618620 129370 618670
rect 129230 618590 129370 618620
rect 129230 618510 129260 618590
rect 129340 618510 129370 618590
rect 129230 618480 129370 618510
rect 129680 618620 129710 618670
rect 129570 618590 129710 618620
rect 129570 618510 129600 618590
rect 129680 618510 129710 618590
rect 129570 618480 129710 618510
rect 130020 618620 130050 618670
rect 129910 618590 130050 618620
rect 129910 618510 129940 618590
rect 130020 618510 130050 618590
rect 129910 618480 130050 618510
rect 130360 618620 130390 618670
rect 130250 618590 130390 618620
rect 130250 618510 130280 618590
rect 130360 618510 130390 618590
rect 130250 618480 130390 618510
rect 130700 618620 130730 618670
rect 130590 618590 130730 618620
rect 130590 618510 130620 618590
rect 130700 618510 130730 618590
rect 130590 618480 130730 618510
rect 131040 618620 131070 618670
rect 130930 618590 131070 618620
rect 130930 618510 130960 618590
rect 131040 618510 131070 618590
rect 130930 618480 131070 618510
rect 131380 618620 131410 618670
rect 131270 618590 131410 618620
rect 131270 618510 131300 618590
rect 131380 618510 131410 618590
rect 131270 618480 131410 618510
rect 131720 618620 131750 618670
rect 131610 618590 131750 618620
rect 131610 618510 131640 618590
rect 131720 618510 131750 618590
rect 131610 618480 131750 618510
rect 125180 611950 125210 612000
rect 125070 611920 125210 611950
rect 125070 611840 125100 611920
rect 125180 611840 125210 611920
rect 125070 611810 125210 611840
rect 125250 611170 125280 611220
rect 125140 611140 125280 611170
rect 125140 610910 125170 611140
rect 125250 610910 125280 611140
rect 125140 610880 125280 610910
rect 125590 611170 125620 611220
rect 125480 611140 125620 611170
rect 125480 610910 125510 611140
rect 125590 610910 125620 611140
rect 125480 610880 125620 610910
rect 125930 611170 125960 611220
rect 125820 611140 125960 611170
rect 125820 610910 125850 611140
rect 125930 610910 125960 611140
rect 125820 610880 125960 610910
rect 126270 611170 126300 611220
rect 126160 611140 126300 611170
rect 126160 610910 126190 611140
rect 126270 610910 126300 611140
rect 126160 610880 126300 610910
rect 126610 611170 126640 611220
rect 126500 611140 126640 611170
rect 126500 610910 126530 611140
rect 126610 610910 126640 611140
rect 126500 610880 126640 610910
rect 126950 611170 126980 611220
rect 126840 611140 126980 611170
rect 126840 610910 126870 611140
rect 126950 610910 126980 611140
rect 126840 610880 126980 610910
rect 127290 611170 127320 611220
rect 127180 611140 127320 611170
rect 127180 610910 127210 611140
rect 127290 610910 127320 611140
rect 127180 610880 127320 610910
rect 127630 611170 127660 611220
rect 127520 611140 127660 611170
rect 127520 610910 127550 611140
rect 127630 610910 127660 611140
rect 127520 610880 127660 610910
rect 127970 611170 128000 611220
rect 127860 611140 128000 611170
rect 127860 610910 127890 611140
rect 127970 610910 128000 611140
rect 127860 610880 128000 610910
rect 128310 611170 128340 611220
rect 128200 611140 128340 611170
rect 128200 610910 128230 611140
rect 128310 610910 128340 611140
rect 128200 610880 128340 610910
rect 128650 611170 128680 611220
rect 128540 611140 128680 611170
rect 128540 610910 128570 611140
rect 128650 610910 128680 611140
rect 128540 610880 128680 610910
rect 128990 611170 129020 611220
rect 128880 611140 129020 611170
rect 128880 610910 128910 611140
rect 128990 610910 129020 611140
rect 128880 610880 129020 610910
rect 129330 611170 129360 611220
rect 129220 611140 129360 611170
rect 129220 610910 129250 611140
rect 129330 610910 129360 611140
rect 129220 610880 129360 610910
rect 129670 611170 129700 611220
rect 129560 611140 129700 611170
rect 129560 610910 129590 611140
rect 129670 610910 129700 611140
rect 129560 610880 129700 610910
rect 130010 611170 130040 611220
rect 129900 611140 130040 611170
rect 129900 610910 129930 611140
rect 130010 610910 130040 611140
rect 129900 610880 130040 610910
rect 130350 611170 130380 611220
rect 130240 611140 130380 611170
rect 130240 610910 130270 611140
rect 130350 610910 130380 611140
rect 130240 610880 130380 610910
rect 130690 611170 130720 611220
rect 130580 611140 130720 611170
rect 130580 610910 130610 611140
rect 130690 610910 130720 611140
rect 130580 610880 130720 610910
rect 131030 611170 131060 611220
rect 130920 611140 131060 611170
rect 130920 610910 130950 611140
rect 131030 610910 131060 611140
rect 130920 610880 131060 610910
rect 131370 611170 131400 611220
rect 131260 611140 131400 611170
rect 131260 610910 131290 611140
rect 131370 610910 131400 611140
rect 131260 610880 131400 610910
rect 125310 605900 125340 605950
rect 125200 605870 125340 605900
rect 125200 605790 125230 605870
rect 125310 605790 125340 605870
rect 125200 605760 125340 605790
rect 125380 605120 125410 605170
rect 125270 605090 125410 605120
rect 125270 604760 125300 605090
rect 125380 604760 125410 605090
rect 125270 604730 125410 604760
rect 125720 605120 125750 605170
rect 125610 605090 125750 605120
rect 125610 604760 125640 605090
rect 125720 604760 125750 605090
rect 125610 604730 125750 604760
rect 126060 605120 126090 605170
rect 125950 605090 126090 605120
rect 125950 604760 125980 605090
rect 126060 604760 126090 605090
rect 125950 604730 126090 604760
rect 126400 605120 126430 605170
rect 126290 605090 126430 605120
rect 126290 604760 126320 605090
rect 126400 604760 126430 605090
rect 126290 604730 126430 604760
rect 126740 605120 126770 605170
rect 126630 605090 126770 605120
rect 126630 604760 126660 605090
rect 126740 604760 126770 605090
rect 126630 604730 126770 604760
rect 127080 605120 127110 605170
rect 126970 605090 127110 605120
rect 126970 604760 127000 605090
rect 127080 604760 127110 605090
rect 126970 604730 127110 604760
rect 127420 605120 127450 605170
rect 127310 605090 127450 605120
rect 127310 604760 127340 605090
rect 127420 604760 127450 605090
rect 127310 604730 127450 604760
rect 127760 605120 127790 605170
rect 127650 605090 127790 605120
rect 127650 604760 127680 605090
rect 127760 604760 127790 605090
rect 127650 604730 127790 604760
rect 128100 605120 128130 605170
rect 127990 605090 128130 605120
rect 127990 604760 128020 605090
rect 128100 604760 128130 605090
rect 127990 604730 128130 604760
rect 128440 605120 128470 605170
rect 128330 605090 128470 605120
rect 128330 604760 128360 605090
rect 128440 604760 128470 605090
rect 128330 604730 128470 604760
rect 128780 605120 128810 605170
rect 128670 605090 128810 605120
rect 128670 604760 128700 605090
rect 128780 604760 128810 605090
rect 128670 604730 128810 604760
rect 129120 605120 129150 605170
rect 129010 605090 129150 605120
rect 129010 604760 129040 605090
rect 129120 604760 129150 605090
rect 129010 604730 129150 604760
rect 129460 605120 129490 605170
rect 129350 605090 129490 605120
rect 129350 604760 129380 605090
rect 129460 604760 129490 605090
rect 129350 604730 129490 604760
rect 129800 605120 129830 605170
rect 129690 605090 129830 605120
rect 129690 604760 129720 605090
rect 129800 604760 129830 605090
rect 129690 604730 129830 604760
rect 130140 605120 130170 605170
rect 130030 605090 130170 605120
rect 130030 604760 130060 605090
rect 130140 604760 130170 605090
rect 130030 604730 130170 604760
rect 130480 605120 130510 605170
rect 130370 605090 130510 605120
rect 130370 604760 130400 605090
rect 130480 604760 130510 605090
rect 130370 604730 130510 604760
rect 130820 605120 130850 605170
rect 130710 605090 130850 605120
rect 130710 604760 130740 605090
rect 130820 604760 130850 605090
rect 130710 604730 130850 604760
rect 131160 605120 131190 605170
rect 131050 605090 131190 605120
rect 131050 604760 131080 605090
rect 131160 604760 131190 605090
rect 131050 604730 131190 604760
rect 131500 605120 131530 605170
rect 131390 605090 131530 605120
rect 131390 604760 131420 605090
rect 131500 604760 131530 605090
rect 131390 604730 131530 604760
rect 125110 599640 125140 599690
rect 125000 599610 125140 599640
rect 125000 599530 125030 599610
rect 125110 599530 125140 599610
rect 125000 599500 125140 599530
rect 125180 598860 125210 598910
rect 125070 598830 125210 598860
rect 125070 598400 125100 598830
rect 125180 598400 125210 598830
rect 125070 598370 125210 598400
rect 125520 598860 125550 598910
rect 125410 598830 125550 598860
rect 125410 598400 125440 598830
rect 125520 598400 125550 598830
rect 125410 598370 125550 598400
rect 125860 598860 125890 598910
rect 125750 598830 125890 598860
rect 125750 598400 125780 598830
rect 125860 598400 125890 598830
rect 125750 598370 125890 598400
rect 126200 598860 126230 598910
rect 126090 598830 126230 598860
rect 126090 598400 126120 598830
rect 126200 598400 126230 598830
rect 126090 598370 126230 598400
rect 126540 598860 126570 598910
rect 126430 598830 126570 598860
rect 126430 598400 126460 598830
rect 126540 598400 126570 598830
rect 126430 598370 126570 598400
rect 126880 598860 126910 598910
rect 126770 598830 126910 598860
rect 126770 598400 126800 598830
rect 126880 598400 126910 598830
rect 126770 598370 126910 598400
rect 127220 598860 127250 598910
rect 127110 598830 127250 598860
rect 127110 598400 127140 598830
rect 127220 598400 127250 598830
rect 127110 598370 127250 598400
rect 127560 598860 127590 598910
rect 127450 598830 127590 598860
rect 127450 598400 127480 598830
rect 127560 598400 127590 598830
rect 127450 598370 127590 598400
rect 127900 598860 127930 598910
rect 127790 598830 127930 598860
rect 127790 598400 127820 598830
rect 127900 598400 127930 598830
rect 127790 598370 127930 598400
rect 128240 598860 128270 598910
rect 128130 598830 128270 598860
rect 128130 598400 128160 598830
rect 128240 598400 128270 598830
rect 128130 598370 128270 598400
rect 128580 598860 128610 598910
rect 128470 598830 128610 598860
rect 128470 598400 128500 598830
rect 128580 598400 128610 598830
rect 128470 598370 128610 598400
rect 128920 598860 128950 598910
rect 128810 598830 128950 598860
rect 128810 598400 128840 598830
rect 128920 598400 128950 598830
rect 128810 598370 128950 598400
rect 129260 598860 129290 598910
rect 129150 598830 129290 598860
rect 129150 598400 129180 598830
rect 129260 598400 129290 598830
rect 129150 598370 129290 598400
rect 129600 598860 129630 598910
rect 129490 598830 129630 598860
rect 129490 598400 129520 598830
rect 129600 598400 129630 598830
rect 129490 598370 129630 598400
rect 129940 598860 129970 598910
rect 129830 598830 129970 598860
rect 129830 598400 129860 598830
rect 129940 598400 129970 598830
rect 129830 598370 129970 598400
rect 130280 598860 130310 598910
rect 130170 598830 130310 598860
rect 130170 598400 130200 598830
rect 130280 598400 130310 598830
rect 130170 598370 130310 598400
rect 130620 598860 130650 598910
rect 130510 598830 130650 598860
rect 130510 598400 130540 598830
rect 130620 598400 130650 598830
rect 130510 598370 130650 598400
rect 130960 598860 130990 598910
rect 130850 598830 130990 598860
rect 130850 598400 130880 598830
rect 130960 598400 130990 598830
rect 130850 598370 130990 598400
rect 131300 598860 131330 598910
rect 131190 598830 131330 598860
rect 131190 598400 131220 598830
rect 131300 598400 131330 598830
rect 131190 598370 131330 598400
rect 119330 592880 119360 592970
rect 119690 592570 119720 592770
rect 120070 592570 120100 592770
rect 125070 592090 125100 592140
rect 124960 592060 125100 592090
rect 124960 591980 124990 592060
rect 125070 591980 125100 592060
rect 124960 591950 125100 591980
rect 125140 591310 125170 591360
rect 125030 591280 125170 591310
rect 125030 590750 125060 591280
rect 125140 590750 125170 591280
rect 125030 590720 125170 590750
rect 125480 591310 125510 591360
rect 125370 591280 125510 591310
rect 125370 590750 125400 591280
rect 125480 590750 125510 591280
rect 125370 590720 125510 590750
rect 125820 591310 125850 591360
rect 125710 591280 125850 591310
rect 125710 590750 125740 591280
rect 125820 590750 125850 591280
rect 125710 590720 125850 590750
rect 126160 591310 126190 591360
rect 126050 591280 126190 591310
rect 126050 590750 126080 591280
rect 126160 590750 126190 591280
rect 126050 590720 126190 590750
rect 126500 591310 126530 591360
rect 126390 591280 126530 591310
rect 126390 590750 126420 591280
rect 126500 590750 126530 591280
rect 126390 590720 126530 590750
rect 126840 591310 126870 591360
rect 126730 591280 126870 591310
rect 126730 590750 126760 591280
rect 126840 590750 126870 591280
rect 126730 590720 126870 590750
rect 127180 591310 127210 591360
rect 127070 591280 127210 591310
rect 127070 590750 127100 591280
rect 127180 590750 127210 591280
rect 127070 590720 127210 590750
rect 127520 591310 127550 591360
rect 127410 591280 127550 591310
rect 127410 590750 127440 591280
rect 127520 590750 127550 591280
rect 127410 590720 127550 590750
rect 127860 591310 127890 591360
rect 127750 591280 127890 591310
rect 127750 590750 127780 591280
rect 127860 590750 127890 591280
rect 127750 590720 127890 590750
rect 128200 591310 128230 591360
rect 128090 591280 128230 591310
rect 128090 590750 128120 591280
rect 128200 590750 128230 591280
rect 128090 590720 128230 590750
rect 128540 591310 128570 591360
rect 128430 591280 128570 591310
rect 128430 590750 128460 591280
rect 128540 590750 128570 591280
rect 128430 590720 128570 590750
rect 128880 591310 128910 591360
rect 128770 591280 128910 591310
rect 128770 590750 128800 591280
rect 128880 590750 128910 591280
rect 128770 590720 128910 590750
rect 129220 591310 129250 591360
rect 129110 591280 129250 591310
rect 129110 590750 129140 591280
rect 129220 590750 129250 591280
rect 129110 590720 129250 590750
rect 129560 591310 129590 591360
rect 129450 591280 129590 591310
rect 129450 590750 129480 591280
rect 129560 590750 129590 591280
rect 129450 590720 129590 590750
rect 129900 591310 129930 591360
rect 129790 591280 129930 591310
rect 129790 590750 129820 591280
rect 129900 590750 129930 591280
rect 129790 590720 129930 590750
rect 130240 591310 130270 591360
rect 130130 591280 130270 591310
rect 130130 590750 130160 591280
rect 130240 590750 130270 591280
rect 130130 590720 130270 590750
rect 130580 591310 130610 591360
rect 130470 591280 130610 591310
rect 130470 590750 130500 591280
rect 130580 590750 130610 591280
rect 130470 590720 130610 590750
rect 130920 591310 130950 591360
rect 130810 591280 130950 591310
rect 130810 590750 130840 591280
rect 130920 590750 130950 591280
rect 130810 590720 130950 590750
rect 131260 591310 131290 591360
rect 131150 591280 131290 591310
rect 131150 590750 131180 591280
rect 131260 590750 131290 591280
rect 131150 590720 131290 590750
rect 119370 583340 119400 583430
rect 119730 583030 119760 583230
rect 120110 583030 120140 583230
rect 125530 583110 125560 583160
rect 125420 583080 125560 583110
rect 125420 583000 125450 583080
rect 125530 583000 125560 583080
rect 125420 582970 125560 583000
rect 125650 582330 125680 582380
rect 125490 582300 125680 582330
rect 125490 582220 125520 582300
rect 125650 582220 125680 582300
rect 125490 582190 125680 582220
rect 126040 582330 126070 582380
rect 125880 582300 126070 582330
rect 125880 582220 125910 582300
rect 126040 582220 126070 582300
rect 125880 582190 126070 582220
rect 126430 582330 126460 582380
rect 126270 582300 126460 582330
rect 126270 582220 126300 582300
rect 126430 582220 126460 582300
rect 126270 582190 126460 582220
rect 126820 582330 126850 582380
rect 126660 582300 126850 582330
rect 126660 582220 126690 582300
rect 126820 582220 126850 582300
rect 126660 582190 126850 582220
rect 127210 582330 127240 582380
rect 127050 582300 127240 582330
rect 127050 582220 127080 582300
rect 127210 582220 127240 582300
rect 127050 582190 127240 582220
rect 127600 582330 127630 582380
rect 127440 582300 127630 582330
rect 127440 582220 127470 582300
rect 127600 582220 127630 582300
rect 127440 582190 127630 582220
rect 127990 582330 128020 582380
rect 127830 582300 128020 582330
rect 127830 582220 127860 582300
rect 127990 582220 128020 582300
rect 127830 582190 128020 582220
rect 128380 582330 128410 582380
rect 128220 582300 128410 582330
rect 128220 582220 128250 582300
rect 128380 582220 128410 582300
rect 128220 582190 128410 582220
rect 128770 582330 128800 582380
rect 128610 582300 128800 582330
rect 128610 582220 128640 582300
rect 128770 582220 128800 582300
rect 128610 582190 128800 582220
rect 129160 582330 129190 582380
rect 129000 582300 129190 582330
rect 129000 582220 129030 582300
rect 129160 582220 129190 582300
rect 129000 582190 129190 582220
rect 129550 582330 129580 582380
rect 129390 582300 129580 582330
rect 129390 582220 129420 582300
rect 129550 582220 129580 582300
rect 129390 582190 129580 582220
rect 129940 582330 129970 582380
rect 129780 582300 129970 582330
rect 129780 582220 129810 582300
rect 129940 582220 129970 582300
rect 129780 582190 129970 582220
rect 130330 582330 130360 582380
rect 130170 582300 130360 582330
rect 130170 582220 130200 582300
rect 130330 582220 130360 582300
rect 130170 582190 130360 582220
rect 130720 582330 130750 582380
rect 130560 582300 130750 582330
rect 130560 582220 130590 582300
rect 130720 582220 130750 582300
rect 130560 582190 130750 582220
rect 131110 582330 131140 582380
rect 130950 582300 131140 582330
rect 130950 582220 130980 582300
rect 131110 582220 131140 582300
rect 130950 582190 131140 582220
rect 131500 582330 131530 582380
rect 131340 582300 131530 582330
rect 131340 582220 131370 582300
rect 131500 582220 131530 582300
rect 131340 582190 131530 582220
rect 131890 582330 131920 582380
rect 131730 582300 131920 582330
rect 131730 582220 131760 582300
rect 131890 582220 131920 582300
rect 131730 582190 131920 582220
rect 132280 582330 132310 582380
rect 132120 582300 132310 582330
rect 132120 582220 132150 582300
rect 132280 582220 132310 582300
rect 132120 582190 132310 582220
rect 132670 582330 132700 582380
rect 132510 582300 132700 582330
rect 132510 582220 132540 582300
rect 132670 582220 132700 582300
rect 132510 582190 132700 582220
rect 119410 574320 119440 574410
rect 119770 574010 119800 574210
rect 120150 574010 120180 574210
rect 125570 574090 125600 574140
rect 125460 574060 125600 574090
rect 125460 573980 125490 574060
rect 125570 573980 125600 574060
rect 125460 573950 125600 573980
rect 125690 573310 125720 573360
rect 125530 573280 125720 573310
rect 125530 573100 125560 573280
rect 125690 573100 125720 573280
rect 125530 573070 125720 573100
rect 126080 573310 126110 573360
rect 125920 573280 126110 573310
rect 125920 573100 125950 573280
rect 126080 573100 126110 573280
rect 125920 573070 126110 573100
rect 126470 573310 126500 573360
rect 126310 573280 126500 573310
rect 126310 573100 126340 573280
rect 126470 573100 126500 573280
rect 126310 573070 126500 573100
rect 126860 573310 126890 573360
rect 126700 573280 126890 573310
rect 126700 573100 126730 573280
rect 126860 573100 126890 573280
rect 126700 573070 126890 573100
rect 127250 573310 127280 573360
rect 127090 573280 127280 573310
rect 127090 573100 127120 573280
rect 127250 573100 127280 573280
rect 127090 573070 127280 573100
rect 127640 573310 127670 573360
rect 127480 573280 127670 573310
rect 127480 573100 127510 573280
rect 127640 573100 127670 573280
rect 127480 573070 127670 573100
rect 128030 573310 128060 573360
rect 127870 573280 128060 573310
rect 127870 573100 127900 573280
rect 128030 573100 128060 573280
rect 127870 573070 128060 573100
rect 128420 573310 128450 573360
rect 128260 573280 128450 573310
rect 128260 573100 128290 573280
rect 128420 573100 128450 573280
rect 128260 573070 128450 573100
rect 128810 573310 128840 573360
rect 128650 573280 128840 573310
rect 128650 573100 128680 573280
rect 128810 573100 128840 573280
rect 128650 573070 128840 573100
rect 129200 573310 129230 573360
rect 129040 573280 129230 573310
rect 129040 573100 129070 573280
rect 129200 573100 129230 573280
rect 129040 573070 129230 573100
rect 129590 573310 129620 573360
rect 129430 573280 129620 573310
rect 129430 573100 129460 573280
rect 129590 573100 129620 573280
rect 129430 573070 129620 573100
rect 129980 573310 130010 573360
rect 129820 573280 130010 573310
rect 129820 573100 129850 573280
rect 129980 573100 130010 573280
rect 129820 573070 130010 573100
rect 130370 573310 130400 573360
rect 130210 573280 130400 573310
rect 130210 573100 130240 573280
rect 130370 573100 130400 573280
rect 130210 573070 130400 573100
rect 130760 573310 130790 573360
rect 130600 573280 130790 573310
rect 130600 573100 130630 573280
rect 130760 573100 130790 573280
rect 130600 573070 130790 573100
rect 131150 573310 131180 573360
rect 130990 573280 131180 573310
rect 130990 573100 131020 573280
rect 131150 573100 131180 573280
rect 130990 573070 131180 573100
rect 131540 573310 131570 573360
rect 131380 573280 131570 573310
rect 131380 573100 131410 573280
rect 131540 573100 131570 573280
rect 131380 573070 131570 573100
rect 131930 573310 131960 573360
rect 131770 573280 131960 573310
rect 131770 573100 131800 573280
rect 131930 573100 131960 573280
rect 131770 573070 131960 573100
rect 132320 573310 132350 573360
rect 132160 573280 132350 573310
rect 132160 573100 132190 573280
rect 132320 573100 132350 573280
rect 132160 573070 132350 573100
rect 132710 573310 132740 573360
rect 132550 573280 132740 573310
rect 132550 573100 132580 573280
rect 132710 573100 132740 573280
rect 132550 573070 132740 573100
rect 119360 566650 119390 566740
rect 119720 566340 119750 566540
rect 120100 566340 120130 566540
rect 125520 566420 125550 566470
rect 125410 566390 125550 566420
rect 125410 566310 125440 566390
rect 125520 566310 125550 566390
rect 125410 566280 125550 566310
rect 125640 565640 125670 565690
rect 125480 565610 125670 565640
rect 125480 565330 125510 565610
rect 125640 565330 125670 565610
rect 125480 565300 125670 565330
rect 126030 565640 126060 565690
rect 125870 565610 126060 565640
rect 125870 565330 125900 565610
rect 126030 565330 126060 565610
rect 125870 565300 126060 565330
rect 126420 565640 126450 565690
rect 126260 565610 126450 565640
rect 126260 565330 126290 565610
rect 126420 565330 126450 565610
rect 126260 565300 126450 565330
rect 126810 565640 126840 565690
rect 126650 565610 126840 565640
rect 126650 565330 126680 565610
rect 126810 565330 126840 565610
rect 126650 565300 126840 565330
rect 127200 565640 127230 565690
rect 127040 565610 127230 565640
rect 127040 565330 127070 565610
rect 127200 565330 127230 565610
rect 127040 565300 127230 565330
rect 127590 565640 127620 565690
rect 127430 565610 127620 565640
rect 127430 565330 127460 565610
rect 127590 565330 127620 565610
rect 127430 565300 127620 565330
rect 127980 565640 128010 565690
rect 127820 565610 128010 565640
rect 127820 565330 127850 565610
rect 127980 565330 128010 565610
rect 127820 565300 128010 565330
rect 128370 565640 128400 565690
rect 128210 565610 128400 565640
rect 128210 565330 128240 565610
rect 128370 565330 128400 565610
rect 128210 565300 128400 565330
rect 128760 565640 128790 565690
rect 128600 565610 128790 565640
rect 128600 565330 128630 565610
rect 128760 565330 128790 565610
rect 128600 565300 128790 565330
rect 129150 565640 129180 565690
rect 128990 565610 129180 565640
rect 128990 565330 129020 565610
rect 129150 565330 129180 565610
rect 128990 565300 129180 565330
rect 129540 565640 129570 565690
rect 129380 565610 129570 565640
rect 129380 565330 129410 565610
rect 129540 565330 129570 565610
rect 129380 565300 129570 565330
rect 129930 565640 129960 565690
rect 129770 565610 129960 565640
rect 129770 565330 129800 565610
rect 129930 565330 129960 565610
rect 129770 565300 129960 565330
rect 130320 565640 130350 565690
rect 130160 565610 130350 565640
rect 130160 565330 130190 565610
rect 130320 565330 130350 565610
rect 130160 565300 130350 565330
rect 130710 565640 130740 565690
rect 130550 565610 130740 565640
rect 130550 565330 130580 565610
rect 130710 565330 130740 565610
rect 130550 565300 130740 565330
rect 131100 565640 131130 565690
rect 130940 565610 131130 565640
rect 130940 565330 130970 565610
rect 131100 565330 131130 565610
rect 130940 565300 131130 565330
rect 131490 565640 131520 565690
rect 131330 565610 131520 565640
rect 131330 565330 131360 565610
rect 131490 565330 131520 565610
rect 131330 565300 131520 565330
rect 131880 565640 131910 565690
rect 131720 565610 131910 565640
rect 131720 565330 131750 565610
rect 131880 565330 131910 565610
rect 131720 565300 131910 565330
rect 132270 565640 132300 565690
rect 132110 565610 132300 565640
rect 132110 565330 132140 565610
rect 132270 565330 132300 565610
rect 132110 565300 132300 565330
rect 132660 565640 132690 565690
rect 132500 565610 132690 565640
rect 132500 565330 132530 565610
rect 132660 565330 132690 565610
rect 132500 565300 132690 565330
rect 119360 560110 119390 560200
rect 119720 559800 119750 560000
rect 120100 559800 120130 560000
rect 125520 559880 125550 559930
rect 125410 559850 125550 559880
rect 125410 559770 125440 559850
rect 125520 559770 125550 559850
rect 125410 559740 125550 559770
rect 125640 559100 125670 559150
rect 125480 559070 125670 559100
rect 125480 558690 125510 559070
rect 125640 558690 125670 559070
rect 125480 558660 125670 558690
rect 126030 559100 126060 559150
rect 125870 559070 126060 559100
rect 125870 558690 125900 559070
rect 126030 558690 126060 559070
rect 125870 558660 126060 558690
rect 126420 559100 126450 559150
rect 126260 559070 126450 559100
rect 126260 558690 126290 559070
rect 126420 558690 126450 559070
rect 126260 558660 126450 558690
rect 126810 559100 126840 559150
rect 126650 559070 126840 559100
rect 126650 558690 126680 559070
rect 126810 558690 126840 559070
rect 126650 558660 126840 558690
rect 127200 559100 127230 559150
rect 127040 559070 127230 559100
rect 127040 558690 127070 559070
rect 127200 558690 127230 559070
rect 127040 558660 127230 558690
rect 127590 559100 127620 559150
rect 127430 559070 127620 559100
rect 127430 558690 127460 559070
rect 127590 558690 127620 559070
rect 127430 558660 127620 558690
rect 127980 559100 128010 559150
rect 127820 559070 128010 559100
rect 127820 558690 127850 559070
rect 127980 558690 128010 559070
rect 127820 558660 128010 558690
rect 128370 559100 128400 559150
rect 128210 559070 128400 559100
rect 128210 558690 128240 559070
rect 128370 558690 128400 559070
rect 128210 558660 128400 558690
rect 128760 559100 128790 559150
rect 128600 559070 128790 559100
rect 128600 558690 128630 559070
rect 128760 558690 128790 559070
rect 128600 558660 128790 558690
rect 129150 559100 129180 559150
rect 128990 559070 129180 559100
rect 128990 558690 129020 559070
rect 129150 558690 129180 559070
rect 128990 558660 129180 558690
rect 129540 559100 129570 559150
rect 129380 559070 129570 559100
rect 129380 558690 129410 559070
rect 129540 558690 129570 559070
rect 129380 558660 129570 558690
rect 129930 559100 129960 559150
rect 129770 559070 129960 559100
rect 129770 558690 129800 559070
rect 129930 558690 129960 559070
rect 129770 558660 129960 558690
rect 130320 559100 130350 559150
rect 130160 559070 130350 559100
rect 130160 558690 130190 559070
rect 130320 558690 130350 559070
rect 130160 558660 130350 558690
rect 130710 559100 130740 559150
rect 130550 559070 130740 559100
rect 130550 558690 130580 559070
rect 130710 558690 130740 559070
rect 130550 558660 130740 558690
rect 131100 559100 131130 559150
rect 130940 559070 131130 559100
rect 130940 558690 130970 559070
rect 131100 558690 131130 559070
rect 130940 558660 131130 558690
rect 131490 559100 131520 559150
rect 131330 559070 131520 559100
rect 131330 558690 131360 559070
rect 131490 558690 131520 559070
rect 131330 558660 131520 558690
rect 131880 559100 131910 559150
rect 131720 559070 131910 559100
rect 131720 558690 131750 559070
rect 131880 558690 131910 559070
rect 131720 558660 131910 558690
rect 132270 559100 132300 559150
rect 132110 559070 132300 559100
rect 132110 558690 132140 559070
rect 132270 558690 132300 559070
rect 132110 558660 132300 558690
rect 132660 559100 132690 559150
rect 132500 559070 132690 559100
rect 132500 558690 132530 559070
rect 132660 558690 132690 559070
rect 132500 558660 132690 558690
rect 125170 554020 125200 554070
rect 125060 553990 125200 554020
rect 125060 553910 125090 553990
rect 125170 553910 125200 553990
rect 125060 553880 125200 553910
rect 119430 553280 119460 553370
rect 119790 552970 119820 553170
rect 120170 552970 120200 553170
rect 125760 552270 125790 552320
rect 125550 552240 125790 552270
rect 125550 552160 125580 552240
rect 125760 552160 125790 552240
rect 125550 552130 125790 552160
rect 126200 552270 126230 552320
rect 125990 552240 126230 552270
rect 125990 552160 126020 552240
rect 126200 552160 126230 552240
rect 125990 552130 126230 552160
rect 126640 552270 126670 552320
rect 126430 552240 126670 552270
rect 126430 552160 126460 552240
rect 126640 552160 126670 552240
rect 126430 552130 126670 552160
rect 127080 552270 127110 552320
rect 126870 552240 127110 552270
rect 126870 552160 126900 552240
rect 127080 552160 127110 552240
rect 126870 552130 127110 552160
rect 127520 552270 127550 552320
rect 127310 552240 127550 552270
rect 127310 552160 127340 552240
rect 127520 552160 127550 552240
rect 127310 552130 127550 552160
rect 127960 552270 127990 552320
rect 127750 552240 127990 552270
rect 127750 552160 127780 552240
rect 127960 552160 127990 552240
rect 127750 552130 127990 552160
rect 128400 552270 128430 552320
rect 128190 552240 128430 552270
rect 128190 552160 128220 552240
rect 128400 552160 128430 552240
rect 128190 552130 128430 552160
rect 128840 552270 128870 552320
rect 128630 552240 128870 552270
rect 128630 552160 128660 552240
rect 128840 552160 128870 552240
rect 128630 552130 128870 552160
rect 129280 552270 129310 552320
rect 129070 552240 129310 552270
rect 129070 552160 129100 552240
rect 129280 552160 129310 552240
rect 129070 552130 129310 552160
rect 129720 552270 129750 552320
rect 129510 552240 129750 552270
rect 129510 552160 129540 552240
rect 129720 552160 129750 552240
rect 129510 552130 129750 552160
rect 130160 552270 130190 552320
rect 129950 552240 130190 552270
rect 129950 552160 129980 552240
rect 130160 552160 130190 552240
rect 129950 552130 130190 552160
rect 130600 552270 130630 552320
rect 130390 552240 130630 552270
rect 130390 552160 130420 552240
rect 130600 552160 130630 552240
rect 130390 552130 130630 552160
rect 131040 552270 131070 552320
rect 130830 552240 131070 552270
rect 130830 552160 130860 552240
rect 131040 552160 131070 552240
rect 130830 552130 131070 552160
rect 131480 552270 131510 552320
rect 131270 552240 131510 552270
rect 131270 552160 131300 552240
rect 131480 552160 131510 552240
rect 131270 552130 131510 552160
rect 131920 552270 131950 552320
rect 131710 552240 131950 552270
rect 131710 552160 131740 552240
rect 131920 552160 131950 552240
rect 131710 552130 131950 552160
rect 132360 552270 132390 552320
rect 132150 552240 132390 552270
rect 132150 552160 132180 552240
rect 132360 552160 132390 552240
rect 132150 552130 132390 552160
rect 132800 552270 132830 552320
rect 132590 552240 132830 552270
rect 132590 552160 132620 552240
rect 132800 552160 132830 552240
rect 132590 552130 132830 552160
rect 133240 552270 133270 552320
rect 133030 552240 133270 552270
rect 133030 552160 133060 552240
rect 133240 552160 133270 552240
rect 133030 552130 133270 552160
rect 133680 552270 133710 552320
rect 133470 552240 133710 552270
rect 133470 552160 133500 552240
rect 133680 552160 133710 552240
rect 133470 552130 133710 552160
rect 125170 546450 125200 546500
rect 125060 546420 125200 546450
rect 125060 546340 125090 546420
rect 125170 546340 125200 546420
rect 125060 546310 125200 546340
rect 119430 545710 119460 545800
rect 119790 545400 119820 545600
rect 120170 545400 120200 545600
rect 125760 544700 125790 544750
rect 125550 544670 125790 544700
rect 125550 544390 125580 544670
rect 125760 544390 125790 544670
rect 125550 544360 125790 544390
rect 126200 544700 126230 544750
rect 125990 544670 126230 544700
rect 125990 544390 126020 544670
rect 126200 544390 126230 544670
rect 125990 544360 126230 544390
rect 126640 544700 126670 544750
rect 126430 544670 126670 544700
rect 126430 544390 126460 544670
rect 126640 544390 126670 544670
rect 126430 544360 126670 544390
rect 127080 544700 127110 544750
rect 126870 544670 127110 544700
rect 126870 544390 126900 544670
rect 127080 544390 127110 544670
rect 126870 544360 127110 544390
rect 127520 544700 127550 544750
rect 127310 544670 127550 544700
rect 127310 544390 127340 544670
rect 127520 544390 127550 544670
rect 127310 544360 127550 544390
rect 127960 544700 127990 544750
rect 127750 544670 127990 544700
rect 127750 544390 127780 544670
rect 127960 544390 127990 544670
rect 127750 544360 127990 544390
rect 128400 544700 128430 544750
rect 128190 544670 128430 544700
rect 128190 544390 128220 544670
rect 128400 544390 128430 544670
rect 128190 544360 128430 544390
rect 128840 544700 128870 544750
rect 128630 544670 128870 544700
rect 128630 544390 128660 544670
rect 128840 544390 128870 544670
rect 128630 544360 128870 544390
rect 129280 544700 129310 544750
rect 129070 544670 129310 544700
rect 129070 544390 129100 544670
rect 129280 544390 129310 544670
rect 129070 544360 129310 544390
rect 129720 544700 129750 544750
rect 129510 544670 129750 544700
rect 129510 544390 129540 544670
rect 129720 544390 129750 544670
rect 129510 544360 129750 544390
rect 130160 544700 130190 544750
rect 129950 544670 130190 544700
rect 129950 544390 129980 544670
rect 130160 544390 130190 544670
rect 129950 544360 130190 544390
rect 130600 544700 130630 544750
rect 130390 544670 130630 544700
rect 130390 544390 130420 544670
rect 130600 544390 130630 544670
rect 130390 544360 130630 544390
rect 131040 544700 131070 544750
rect 130830 544670 131070 544700
rect 130830 544390 130860 544670
rect 131040 544390 131070 544670
rect 130830 544360 131070 544390
rect 131480 544700 131510 544750
rect 131270 544670 131510 544700
rect 131270 544390 131300 544670
rect 131480 544390 131510 544670
rect 131270 544360 131510 544390
rect 131920 544700 131950 544750
rect 131710 544670 131950 544700
rect 131710 544390 131740 544670
rect 131920 544390 131950 544670
rect 131710 544360 131950 544390
rect 132360 544700 132390 544750
rect 132150 544670 132390 544700
rect 132150 544390 132180 544670
rect 132360 544390 132390 544670
rect 132150 544360 132390 544390
rect 132800 544700 132830 544750
rect 132590 544670 132830 544700
rect 132590 544390 132620 544670
rect 132800 544390 132830 544670
rect 132590 544360 132830 544390
rect 133240 544700 133270 544750
rect 133030 544670 133270 544700
rect 133030 544390 133060 544670
rect 133240 544390 133270 544670
rect 133030 544360 133270 544390
rect 133680 544700 133710 544750
rect 133470 544670 133710 544700
rect 133470 544390 133500 544670
rect 133680 544390 133710 544670
rect 133470 544360 133710 544390
rect 125140 538390 125170 538440
rect 125030 538360 125170 538390
rect 125030 538280 125060 538360
rect 125140 538280 125170 538360
rect 125030 538250 125170 538280
rect 119400 537650 119430 537740
rect 119760 537340 119790 537540
rect 120140 537340 120170 537540
rect 125730 536640 125760 536690
rect 125520 536610 125760 536640
rect 125520 536130 125550 536610
rect 125730 536130 125760 536610
rect 125520 536100 125760 536130
rect 126170 536640 126200 536690
rect 125960 536610 126200 536640
rect 125960 536130 125990 536610
rect 126170 536130 126200 536610
rect 125960 536100 126200 536130
rect 126610 536640 126640 536690
rect 126400 536610 126640 536640
rect 126400 536130 126430 536610
rect 126610 536130 126640 536610
rect 126400 536100 126640 536130
rect 127050 536640 127080 536690
rect 126840 536610 127080 536640
rect 126840 536130 126870 536610
rect 127050 536130 127080 536610
rect 126840 536100 127080 536130
rect 127490 536640 127520 536690
rect 127280 536610 127520 536640
rect 127280 536130 127310 536610
rect 127490 536130 127520 536610
rect 127280 536100 127520 536130
rect 127930 536640 127960 536690
rect 127720 536610 127960 536640
rect 127720 536130 127750 536610
rect 127930 536130 127960 536610
rect 127720 536100 127960 536130
rect 128370 536640 128400 536690
rect 128160 536610 128400 536640
rect 128160 536130 128190 536610
rect 128370 536130 128400 536610
rect 128160 536100 128400 536130
rect 128810 536640 128840 536690
rect 128600 536610 128840 536640
rect 128600 536130 128630 536610
rect 128810 536130 128840 536610
rect 128600 536100 128840 536130
rect 129250 536640 129280 536690
rect 129040 536610 129280 536640
rect 129040 536130 129070 536610
rect 129250 536130 129280 536610
rect 129040 536100 129280 536130
rect 129690 536640 129720 536690
rect 129480 536610 129720 536640
rect 129480 536130 129510 536610
rect 129690 536130 129720 536610
rect 129480 536100 129720 536130
rect 130130 536640 130160 536690
rect 129920 536610 130160 536640
rect 129920 536130 129950 536610
rect 130130 536130 130160 536610
rect 129920 536100 130160 536130
rect 130570 536640 130600 536690
rect 130360 536610 130600 536640
rect 130360 536130 130390 536610
rect 130570 536130 130600 536610
rect 130360 536100 130600 536130
rect 131010 536640 131040 536690
rect 130800 536610 131040 536640
rect 130800 536130 130830 536610
rect 131010 536130 131040 536610
rect 130800 536100 131040 536130
rect 131450 536640 131480 536690
rect 131240 536610 131480 536640
rect 131240 536130 131270 536610
rect 131450 536130 131480 536610
rect 131240 536100 131480 536130
rect 131890 536640 131920 536690
rect 131680 536610 131920 536640
rect 131680 536130 131710 536610
rect 131890 536130 131920 536610
rect 131680 536100 131920 536130
rect 132330 536640 132360 536690
rect 132120 536610 132360 536640
rect 132120 536130 132150 536610
rect 132330 536130 132360 536610
rect 132120 536100 132360 536130
rect 132770 536640 132800 536690
rect 132560 536610 132800 536640
rect 132560 536130 132590 536610
rect 132770 536130 132800 536610
rect 132560 536100 132800 536130
rect 133210 536640 133240 536690
rect 133000 536610 133240 536640
rect 133000 536130 133030 536610
rect 133210 536130 133240 536610
rect 133000 536100 133240 536130
rect 133650 536640 133680 536690
rect 133440 536610 133680 536640
rect 133440 536130 133470 536610
rect 133650 536130 133680 536610
rect 133440 536100 133680 536130
<< pmos >>
rect 119330 593160 119360 593250
rect 119690 593080 119720 593280
rect 120070 593080 120100 593280
rect 119370 583620 119400 583710
rect 119730 583540 119760 583740
rect 120110 583540 120140 583740
rect 119410 574600 119440 574690
rect 119770 574520 119800 574720
rect 120150 574520 120180 574720
rect 119360 566930 119390 567020
rect 119720 566850 119750 567050
rect 120100 566850 120130 567050
rect 119360 560390 119390 560480
rect 119720 560310 119750 560510
rect 120100 560310 120130 560510
rect 119430 553560 119460 553650
rect 119790 553480 119820 553680
rect 120170 553480 120200 553680
rect 119430 545990 119460 546080
rect 119790 545910 119820 546110
rect 120170 545910 120200 546110
rect 119400 537930 119430 538020
rect 119760 537850 119790 538050
rect 120140 537850 120170 538050
<< ndiff >>
rect 124150 642400 124240 642410
rect 124150 642360 124170 642400
rect 124220 642360 124240 642400
rect 124150 642340 124240 642360
rect 124330 642400 124420 642410
rect 124330 642360 124350 642400
rect 124400 642360 124420 642400
rect 124330 642340 124420 642360
rect 124510 642400 124600 642410
rect 124510 642360 124530 642400
rect 124580 642360 124600 642400
rect 124510 642340 124600 642360
rect 124690 642400 124780 642410
rect 124690 642360 124710 642400
rect 124760 642360 124780 642400
rect 124690 642340 124780 642360
rect 124870 642400 124960 642410
rect 124870 642360 124890 642400
rect 124940 642360 124960 642400
rect 124870 642340 124960 642360
rect 125050 642400 125140 642410
rect 125050 642360 125070 642400
rect 125120 642360 125140 642400
rect 125050 642340 125140 642360
rect 125230 642400 125320 642410
rect 125230 642360 125250 642400
rect 125300 642360 125320 642400
rect 125230 642340 125320 642360
rect 125410 642400 125500 642410
rect 125410 642360 125430 642400
rect 125480 642360 125500 642400
rect 125410 642340 125500 642360
rect 125590 642400 125680 642410
rect 125590 642360 125610 642400
rect 125660 642360 125680 642400
rect 125590 642340 125680 642360
rect 125770 642400 125860 642410
rect 125770 642360 125790 642400
rect 125840 642360 125860 642400
rect 125770 642340 125860 642360
rect 125950 642400 126040 642410
rect 125950 642360 125970 642400
rect 126020 642360 126040 642400
rect 125950 642340 126040 642360
rect 126130 642400 126220 642410
rect 126130 642360 126150 642400
rect 126200 642360 126220 642400
rect 126130 642340 126220 642360
rect 126310 642400 126400 642410
rect 126310 642360 126330 642400
rect 126380 642360 126400 642400
rect 126310 642340 126400 642360
rect 126490 642400 126580 642410
rect 126490 642360 126510 642400
rect 126560 642360 126580 642400
rect 126490 642340 126580 642360
rect 126670 642400 126760 642410
rect 126670 642360 126690 642400
rect 126740 642360 126760 642400
rect 126670 642340 126760 642360
rect 126850 642400 126940 642410
rect 126850 642360 126870 642400
rect 126920 642360 126940 642400
rect 126850 642340 126940 642360
rect 127030 642400 127120 642410
rect 127030 642360 127050 642400
rect 127100 642360 127120 642400
rect 127030 642340 127120 642360
rect 127210 642400 127300 642410
rect 127210 642360 127230 642400
rect 127280 642360 127300 642400
rect 127210 642340 127300 642360
rect 127390 642400 127480 642410
rect 127390 642360 127410 642400
rect 127460 642360 127480 642400
rect 127390 642340 127480 642360
rect 127570 642400 127660 642410
rect 127570 642360 127590 642400
rect 127640 642360 127660 642400
rect 127570 642340 127660 642360
rect 127750 642400 127840 642410
rect 127750 642360 127770 642400
rect 127820 642360 127840 642400
rect 127750 642340 127840 642360
rect 127930 642400 128020 642410
rect 127930 642360 127950 642400
rect 128000 642360 128020 642400
rect 127930 642340 128020 642360
rect 128110 642400 128200 642410
rect 128110 642360 128130 642400
rect 128180 642360 128200 642400
rect 128110 642340 128200 642360
rect 128290 642400 128380 642410
rect 128290 642360 128310 642400
rect 128360 642360 128380 642400
rect 128290 642340 128380 642360
rect 128470 642400 128560 642410
rect 128470 642360 128490 642400
rect 128540 642360 128560 642400
rect 128470 642340 128560 642360
rect 128650 642400 128740 642410
rect 128650 642360 128670 642400
rect 128720 642360 128740 642400
rect 128650 642340 128740 642360
rect 128830 642400 128920 642410
rect 128830 642360 128850 642400
rect 128900 642360 128920 642400
rect 128830 642340 128920 642360
rect 129010 642400 129100 642410
rect 129010 642360 129030 642400
rect 129080 642360 129100 642400
rect 129010 642340 129100 642360
rect 129190 642400 129280 642410
rect 129190 642360 129210 642400
rect 129260 642360 129280 642400
rect 129190 642340 129280 642360
rect 129370 642400 129460 642410
rect 129370 642360 129390 642400
rect 129440 642360 129460 642400
rect 129370 642340 129460 642360
rect 129550 642400 129640 642410
rect 129550 642360 129570 642400
rect 129620 642360 129640 642400
rect 129550 642340 129640 642360
rect 129730 642400 129820 642410
rect 129730 642360 129750 642400
rect 129800 642360 129820 642400
rect 129730 642340 129820 642360
rect 129910 642400 130000 642410
rect 129910 642360 129930 642400
rect 129980 642360 130000 642400
rect 129910 642340 130000 642360
rect 130090 642400 130180 642410
rect 130090 642360 130110 642400
rect 130160 642360 130180 642400
rect 130090 642340 130180 642360
rect 130270 642400 130360 642410
rect 130270 642360 130290 642400
rect 130340 642360 130360 642400
rect 130270 642340 130360 642360
rect 130450 642400 130540 642410
rect 130450 642360 130470 642400
rect 130520 642360 130540 642400
rect 130450 642340 130540 642360
rect 130630 642400 130720 642410
rect 130630 642360 130650 642400
rect 130700 642360 130720 642400
rect 130630 642340 130720 642360
rect 130810 642400 130900 642410
rect 130810 642360 130830 642400
rect 130880 642360 130900 642400
rect 130810 642340 130900 642360
rect 130990 642400 131080 642410
rect 130990 642360 131010 642400
rect 131060 642360 131080 642400
rect 130990 642340 131080 642360
rect 131170 642400 131260 642410
rect 131170 642360 131190 642400
rect 131240 642360 131260 642400
rect 131170 642340 131260 642360
rect 124150 642290 124240 642310
rect 124150 642250 124170 642290
rect 124220 642250 124240 642290
rect 124150 642240 124240 642250
rect 124330 642290 124420 642310
rect 124330 642250 124350 642290
rect 124400 642250 124420 642290
rect 124330 642240 124420 642250
rect 124510 642290 124600 642310
rect 124510 642250 124530 642290
rect 124580 642250 124600 642290
rect 124510 642240 124600 642250
rect 124690 642290 124780 642310
rect 124690 642250 124710 642290
rect 124760 642250 124780 642290
rect 124690 642240 124780 642250
rect 124870 642290 124960 642310
rect 124870 642250 124890 642290
rect 124940 642250 124960 642290
rect 124870 642240 124960 642250
rect 125050 642290 125140 642310
rect 125050 642250 125070 642290
rect 125120 642250 125140 642290
rect 125050 642240 125140 642250
rect 125230 642290 125320 642310
rect 125230 642250 125250 642290
rect 125300 642250 125320 642290
rect 125230 642240 125320 642250
rect 125410 642290 125500 642310
rect 125410 642250 125430 642290
rect 125480 642250 125500 642290
rect 125410 642240 125500 642250
rect 125590 642290 125680 642310
rect 125590 642250 125610 642290
rect 125660 642250 125680 642290
rect 125590 642240 125680 642250
rect 125770 642290 125860 642310
rect 125770 642250 125790 642290
rect 125840 642250 125860 642290
rect 125770 642240 125860 642250
rect 125950 642290 126040 642310
rect 125950 642250 125970 642290
rect 126020 642250 126040 642290
rect 125950 642240 126040 642250
rect 126130 642290 126220 642310
rect 126130 642250 126150 642290
rect 126200 642250 126220 642290
rect 126130 642240 126220 642250
rect 126310 642290 126400 642310
rect 126310 642250 126330 642290
rect 126380 642250 126400 642290
rect 126310 642240 126400 642250
rect 126490 642290 126580 642310
rect 126490 642250 126510 642290
rect 126560 642250 126580 642290
rect 126490 642240 126580 642250
rect 126670 642290 126760 642310
rect 126670 642250 126690 642290
rect 126740 642250 126760 642290
rect 126670 642240 126760 642250
rect 126850 642290 126940 642310
rect 126850 642250 126870 642290
rect 126920 642250 126940 642290
rect 126850 642240 126940 642250
rect 127030 642290 127120 642310
rect 127030 642250 127050 642290
rect 127100 642250 127120 642290
rect 127030 642240 127120 642250
rect 127210 642290 127300 642310
rect 127210 642250 127230 642290
rect 127280 642250 127300 642290
rect 127210 642240 127300 642250
rect 127390 642290 127480 642310
rect 127390 642250 127410 642290
rect 127460 642250 127480 642290
rect 127390 642240 127480 642250
rect 127570 642290 127660 642310
rect 127570 642250 127590 642290
rect 127640 642250 127660 642290
rect 127570 642240 127660 642250
rect 127750 642290 127840 642310
rect 127750 642250 127770 642290
rect 127820 642250 127840 642290
rect 127750 642240 127840 642250
rect 127930 642290 128020 642310
rect 127930 642250 127950 642290
rect 128000 642250 128020 642290
rect 127930 642240 128020 642250
rect 128110 642290 128200 642310
rect 128110 642250 128130 642290
rect 128180 642250 128200 642290
rect 128110 642240 128200 642250
rect 128290 642290 128380 642310
rect 128290 642250 128310 642290
rect 128360 642250 128380 642290
rect 128290 642240 128380 642250
rect 128470 642290 128560 642310
rect 128470 642250 128490 642290
rect 128540 642250 128560 642290
rect 128470 642240 128560 642250
rect 128650 642290 128740 642310
rect 128650 642250 128670 642290
rect 128720 642250 128740 642290
rect 128650 642240 128740 642250
rect 128830 642290 128920 642310
rect 128830 642250 128850 642290
rect 128900 642250 128920 642290
rect 128830 642240 128920 642250
rect 129010 642290 129100 642310
rect 129010 642250 129030 642290
rect 129080 642250 129100 642290
rect 129010 642240 129100 642250
rect 129190 642290 129280 642310
rect 129190 642250 129210 642290
rect 129260 642250 129280 642290
rect 129190 642240 129280 642250
rect 129370 642290 129460 642310
rect 129370 642250 129390 642290
rect 129440 642250 129460 642290
rect 129370 642240 129460 642250
rect 129550 642290 129640 642310
rect 129550 642250 129570 642290
rect 129620 642250 129640 642290
rect 129550 642240 129640 642250
rect 129730 642290 129820 642310
rect 129730 642250 129750 642290
rect 129800 642250 129820 642290
rect 129730 642240 129820 642250
rect 129910 642290 130000 642310
rect 129910 642250 129930 642290
rect 129980 642250 130000 642290
rect 129910 642240 130000 642250
rect 130090 642290 130180 642310
rect 130090 642250 130110 642290
rect 130160 642250 130180 642290
rect 130090 642240 130180 642250
rect 130270 642290 130360 642310
rect 130270 642250 130290 642290
rect 130340 642250 130360 642290
rect 130270 642240 130360 642250
rect 130450 642290 130540 642310
rect 130450 642250 130470 642290
rect 130520 642250 130540 642290
rect 130450 642240 130540 642250
rect 130630 642290 130720 642310
rect 130630 642250 130650 642290
rect 130700 642250 130720 642290
rect 130630 642240 130720 642250
rect 130810 642290 130900 642310
rect 130810 642250 130830 642290
rect 130880 642250 130900 642290
rect 130810 642240 130900 642250
rect 130990 642290 131080 642310
rect 130990 642250 131010 642290
rect 131060 642250 131080 642290
rect 130990 642240 131080 642250
rect 131170 642290 131260 642310
rect 131170 642250 131190 642290
rect 131240 642250 131260 642290
rect 131170 642240 131260 642250
rect 124180 636230 124360 636240
rect 124180 636190 124200 636230
rect 124340 636190 124360 636230
rect 124180 636170 124360 636190
rect 124420 636230 124600 636240
rect 124420 636190 124440 636230
rect 124580 636190 124600 636230
rect 124420 636170 124600 636190
rect 124660 636230 124840 636240
rect 124660 636190 124680 636230
rect 124820 636190 124840 636230
rect 124660 636170 124840 636190
rect 124900 636230 125080 636240
rect 124900 636190 124920 636230
rect 125060 636190 125080 636230
rect 124900 636170 125080 636190
rect 125140 636230 125320 636240
rect 125140 636190 125160 636230
rect 125300 636190 125320 636230
rect 125140 636170 125320 636190
rect 125380 636230 125560 636240
rect 125380 636190 125400 636230
rect 125540 636190 125560 636230
rect 125380 636170 125560 636190
rect 125620 636230 125800 636240
rect 125620 636190 125640 636230
rect 125780 636190 125800 636230
rect 125620 636170 125800 636190
rect 125860 636230 126040 636240
rect 125860 636190 125880 636230
rect 126020 636190 126040 636230
rect 125860 636170 126040 636190
rect 126100 636230 126280 636240
rect 126100 636190 126120 636230
rect 126260 636190 126280 636230
rect 126100 636170 126280 636190
rect 126340 636230 126520 636240
rect 126340 636190 126360 636230
rect 126500 636190 126520 636230
rect 126340 636170 126520 636190
rect 126580 636230 126760 636240
rect 126580 636190 126600 636230
rect 126740 636190 126760 636230
rect 126580 636170 126760 636190
rect 126820 636230 127000 636240
rect 126820 636190 126840 636230
rect 126980 636190 127000 636230
rect 126820 636170 127000 636190
rect 127060 636230 127240 636240
rect 127060 636190 127080 636230
rect 127220 636190 127240 636230
rect 127060 636170 127240 636190
rect 127300 636230 127480 636240
rect 127300 636190 127320 636230
rect 127460 636190 127480 636230
rect 127300 636170 127480 636190
rect 127540 636230 127720 636240
rect 127540 636190 127560 636230
rect 127700 636190 127720 636230
rect 127540 636170 127720 636190
rect 127780 636230 127960 636240
rect 127780 636190 127800 636230
rect 127940 636190 127960 636230
rect 127780 636170 127960 636190
rect 128020 636230 128200 636240
rect 128020 636190 128040 636230
rect 128180 636190 128200 636230
rect 128020 636170 128200 636190
rect 128260 636230 128440 636240
rect 128260 636190 128280 636230
rect 128420 636190 128440 636230
rect 128260 636170 128440 636190
rect 128500 636230 128680 636240
rect 128500 636190 128520 636230
rect 128660 636190 128680 636230
rect 128500 636170 128680 636190
rect 128740 636230 128920 636240
rect 128740 636190 128760 636230
rect 128900 636190 128920 636230
rect 128740 636170 128920 636190
rect 124180 636120 124360 636140
rect 124180 636080 124200 636120
rect 124340 636080 124360 636120
rect 124180 636070 124360 636080
rect 124420 636120 124600 636140
rect 124420 636080 124440 636120
rect 124580 636080 124600 636120
rect 124420 636070 124600 636080
rect 124660 636120 124840 636140
rect 124660 636080 124680 636120
rect 124820 636080 124840 636120
rect 124660 636070 124840 636080
rect 124900 636120 125080 636140
rect 124900 636080 124920 636120
rect 125060 636080 125080 636120
rect 124900 636070 125080 636080
rect 125140 636120 125320 636140
rect 125140 636080 125160 636120
rect 125300 636080 125320 636120
rect 125140 636070 125320 636080
rect 125380 636120 125560 636140
rect 125380 636080 125400 636120
rect 125540 636080 125560 636120
rect 125380 636070 125560 636080
rect 125620 636120 125800 636140
rect 125620 636080 125640 636120
rect 125780 636080 125800 636120
rect 125620 636070 125800 636080
rect 125860 636120 126040 636140
rect 125860 636080 125880 636120
rect 126020 636080 126040 636120
rect 125860 636070 126040 636080
rect 126100 636120 126280 636140
rect 126100 636080 126120 636120
rect 126260 636080 126280 636120
rect 126100 636070 126280 636080
rect 126340 636120 126520 636140
rect 126340 636080 126360 636120
rect 126500 636080 126520 636120
rect 126340 636070 126520 636080
rect 126580 636120 126760 636140
rect 126580 636080 126600 636120
rect 126740 636080 126760 636120
rect 126580 636070 126760 636080
rect 126820 636120 127000 636140
rect 126820 636080 126840 636120
rect 126980 636080 127000 636120
rect 126820 636070 127000 636080
rect 127060 636120 127240 636140
rect 127060 636080 127080 636120
rect 127220 636080 127240 636120
rect 127060 636070 127240 636080
rect 127300 636120 127480 636140
rect 127300 636080 127320 636120
rect 127460 636080 127480 636120
rect 127300 636070 127480 636080
rect 127540 636120 127720 636140
rect 127540 636080 127560 636120
rect 127700 636080 127720 636120
rect 127540 636070 127720 636080
rect 127780 636120 127960 636140
rect 127780 636080 127800 636120
rect 127940 636080 127960 636120
rect 127780 636070 127960 636080
rect 128020 636120 128200 636140
rect 128020 636080 128040 636120
rect 128180 636080 128200 636120
rect 128020 636070 128200 636080
rect 128260 636120 128440 636140
rect 128260 636080 128280 636120
rect 128420 636080 128440 636120
rect 128260 636070 128440 636080
rect 128500 636120 128680 636140
rect 128500 636080 128520 636120
rect 128660 636080 128680 636120
rect 128500 636070 128680 636080
rect 128740 636120 128920 636140
rect 128740 636080 128760 636120
rect 128900 636080 128920 636120
rect 128740 636070 128920 636080
rect 124240 632640 124640 632650
rect 124240 632600 124260 632640
rect 124620 632600 124640 632640
rect 124240 632580 124640 632600
rect 124240 632530 124640 632550
rect 124240 632490 124260 632530
rect 124620 632490 124640 632530
rect 124240 632480 124640 632490
rect 124450 630200 124850 630210
rect 124450 630160 124470 630200
rect 124830 630160 124850 630200
rect 124450 630140 124850 630160
rect 124910 630200 125310 630210
rect 124910 630160 124930 630200
rect 125290 630160 125310 630200
rect 124910 630140 125310 630160
rect 125370 630200 125770 630210
rect 125370 630160 125390 630200
rect 125750 630160 125770 630200
rect 125370 630140 125770 630160
rect 125830 630200 126230 630210
rect 125830 630160 125850 630200
rect 126210 630160 126230 630200
rect 125830 630140 126230 630160
rect 126290 630200 126690 630210
rect 126290 630160 126310 630200
rect 126670 630160 126690 630200
rect 126290 630140 126690 630160
rect 126750 630200 127150 630210
rect 126750 630160 126770 630200
rect 127130 630160 127150 630200
rect 126750 630140 127150 630160
rect 127210 630200 127610 630210
rect 127210 630160 127230 630200
rect 127590 630160 127610 630200
rect 127210 630140 127610 630160
rect 127670 630200 128070 630210
rect 127670 630160 127690 630200
rect 128050 630160 128070 630200
rect 127670 630140 128070 630160
rect 128130 630200 128530 630210
rect 128130 630160 128150 630200
rect 128510 630160 128530 630200
rect 128130 630140 128530 630160
rect 128590 630200 128990 630210
rect 128590 630160 128610 630200
rect 128970 630160 128990 630200
rect 128590 630140 128990 630160
rect 124450 630090 124850 630110
rect 124450 630050 124470 630090
rect 124830 630050 124850 630090
rect 124450 630040 124850 630050
rect 124910 630090 125310 630110
rect 124910 630050 124930 630090
rect 125290 630050 125310 630090
rect 124910 630040 125310 630050
rect 125370 630090 125770 630110
rect 125370 630050 125390 630090
rect 125750 630050 125770 630090
rect 125370 630040 125770 630050
rect 125830 630090 126230 630110
rect 125830 630050 125850 630090
rect 126210 630050 126230 630090
rect 125830 630040 126230 630050
rect 126290 630090 126690 630110
rect 126290 630050 126310 630090
rect 126670 630050 126690 630090
rect 126290 630040 126690 630050
rect 126750 630090 127150 630110
rect 126750 630050 126770 630090
rect 127130 630050 127150 630090
rect 126750 630040 127150 630050
rect 127210 630090 127610 630110
rect 127210 630050 127230 630090
rect 127590 630050 127610 630090
rect 127210 630040 127610 630050
rect 127670 630090 128070 630110
rect 127670 630050 127690 630090
rect 128050 630050 128070 630090
rect 127670 630040 128070 630050
rect 128130 630090 128530 630110
rect 128130 630050 128150 630090
rect 128510 630050 128530 630090
rect 128130 630040 128530 630050
rect 128590 630090 128990 630110
rect 128590 630050 128610 630090
rect 128970 630050 128990 630090
rect 128590 630040 128990 630050
rect 124220 624970 124820 624980
rect 124220 624930 124240 624970
rect 124800 624930 124820 624970
rect 124220 624910 124820 624930
rect 124220 624860 124820 624880
rect 124220 624820 124240 624860
rect 124800 624820 124820 624860
rect 124220 624810 124820 624820
rect 124780 623680 125380 623690
rect 124780 623640 124800 623680
rect 125360 623640 125380 623680
rect 124780 623620 125380 623640
rect 125440 623680 126040 623690
rect 125440 623640 125460 623680
rect 126020 623640 126040 623680
rect 125440 623620 126040 623640
rect 126100 623680 126700 623690
rect 126100 623640 126120 623680
rect 126680 623640 126700 623680
rect 126100 623620 126700 623640
rect 126760 623680 127360 623690
rect 126760 623640 126780 623680
rect 127340 623640 127360 623680
rect 126760 623620 127360 623640
rect 127420 623680 128020 623690
rect 127420 623640 127440 623680
rect 128000 623640 128020 623680
rect 127420 623620 128020 623640
rect 128080 623680 128680 623690
rect 128080 623640 128100 623680
rect 128660 623640 128680 623680
rect 128080 623620 128680 623640
rect 124780 623570 125380 623590
rect 124780 623530 124800 623570
rect 125360 623530 125380 623570
rect 124780 623520 125380 623530
rect 125440 623570 126040 623590
rect 125440 623530 125460 623570
rect 126020 623530 126040 623570
rect 125440 623520 126040 623530
rect 126100 623570 126700 623590
rect 126100 623530 126120 623570
rect 126680 623530 126700 623570
rect 126100 623520 126700 623530
rect 126760 623570 127360 623590
rect 126760 623530 126780 623570
rect 127340 623530 127360 623570
rect 126760 623520 127360 623530
rect 127420 623570 128020 623590
rect 127420 623530 127440 623570
rect 128000 623530 128020 623570
rect 127420 623520 128020 623530
rect 128080 623570 128680 623590
rect 128080 623530 128100 623570
rect 128660 623530 128680 623570
rect 128080 623520 128680 623530
rect 125350 619400 125530 619450
rect 125350 619350 125420 619400
rect 125350 619310 125360 619350
rect 125400 619310 125420 619350
rect 125350 619260 125420 619310
rect 125450 619350 125530 619370
rect 125450 619310 125470 619350
rect 125510 619310 125530 619350
rect 125450 619290 125530 619310
rect 125560 619350 125630 619450
rect 125560 619310 125580 619350
rect 125620 619310 125630 619350
rect 125560 619260 125630 619310
rect 125350 619210 125630 619260
rect 125420 618620 125600 618670
rect 125420 618570 125490 618620
rect 125420 618530 125430 618570
rect 125470 618530 125490 618570
rect 125420 618480 125490 618530
rect 125520 618570 125600 618590
rect 125520 618530 125540 618570
rect 125580 618530 125600 618570
rect 125520 618510 125600 618530
rect 125630 618570 125700 618670
rect 125630 618530 125650 618570
rect 125690 618530 125700 618570
rect 125630 618480 125700 618530
rect 125420 618430 125700 618480
rect 125760 618620 125940 618670
rect 125760 618570 125830 618620
rect 125760 618530 125770 618570
rect 125810 618530 125830 618570
rect 125760 618480 125830 618530
rect 125860 618570 125940 618590
rect 125860 618530 125880 618570
rect 125920 618530 125940 618570
rect 125860 618510 125940 618530
rect 125970 618570 126040 618670
rect 125970 618530 125990 618570
rect 126030 618530 126040 618570
rect 125970 618480 126040 618530
rect 125760 618430 126040 618480
rect 126100 618620 126280 618670
rect 126100 618570 126170 618620
rect 126100 618530 126110 618570
rect 126150 618530 126170 618570
rect 126100 618480 126170 618530
rect 126200 618570 126280 618590
rect 126200 618530 126220 618570
rect 126260 618530 126280 618570
rect 126200 618510 126280 618530
rect 126310 618570 126380 618670
rect 126310 618530 126330 618570
rect 126370 618530 126380 618570
rect 126310 618480 126380 618530
rect 126100 618430 126380 618480
rect 126440 618620 126620 618670
rect 126440 618570 126510 618620
rect 126440 618530 126450 618570
rect 126490 618530 126510 618570
rect 126440 618480 126510 618530
rect 126540 618570 126620 618590
rect 126540 618530 126560 618570
rect 126600 618530 126620 618570
rect 126540 618510 126620 618530
rect 126650 618570 126720 618670
rect 126650 618530 126670 618570
rect 126710 618530 126720 618570
rect 126650 618480 126720 618530
rect 126440 618430 126720 618480
rect 126780 618620 126960 618670
rect 126780 618570 126850 618620
rect 126780 618530 126790 618570
rect 126830 618530 126850 618570
rect 126780 618480 126850 618530
rect 126880 618570 126960 618590
rect 126880 618530 126900 618570
rect 126940 618530 126960 618570
rect 126880 618510 126960 618530
rect 126990 618570 127060 618670
rect 126990 618530 127010 618570
rect 127050 618530 127060 618570
rect 126990 618480 127060 618530
rect 126780 618430 127060 618480
rect 127120 618620 127300 618670
rect 127120 618570 127190 618620
rect 127120 618530 127130 618570
rect 127170 618530 127190 618570
rect 127120 618480 127190 618530
rect 127220 618570 127300 618590
rect 127220 618530 127240 618570
rect 127280 618530 127300 618570
rect 127220 618510 127300 618530
rect 127330 618570 127400 618670
rect 127330 618530 127350 618570
rect 127390 618530 127400 618570
rect 127330 618480 127400 618530
rect 127120 618430 127400 618480
rect 127460 618620 127640 618670
rect 127460 618570 127530 618620
rect 127460 618530 127470 618570
rect 127510 618530 127530 618570
rect 127460 618480 127530 618530
rect 127560 618570 127640 618590
rect 127560 618530 127580 618570
rect 127620 618530 127640 618570
rect 127560 618510 127640 618530
rect 127670 618570 127740 618670
rect 127670 618530 127690 618570
rect 127730 618530 127740 618570
rect 127670 618480 127740 618530
rect 127460 618430 127740 618480
rect 127800 618620 127980 618670
rect 127800 618570 127870 618620
rect 127800 618530 127810 618570
rect 127850 618530 127870 618570
rect 127800 618480 127870 618530
rect 127900 618570 127980 618590
rect 127900 618530 127920 618570
rect 127960 618530 127980 618570
rect 127900 618510 127980 618530
rect 128010 618570 128080 618670
rect 128010 618530 128030 618570
rect 128070 618530 128080 618570
rect 128010 618480 128080 618530
rect 127800 618430 128080 618480
rect 128140 618620 128320 618670
rect 128140 618570 128210 618620
rect 128140 618530 128150 618570
rect 128190 618530 128210 618570
rect 128140 618480 128210 618530
rect 128240 618570 128320 618590
rect 128240 618530 128260 618570
rect 128300 618530 128320 618570
rect 128240 618510 128320 618530
rect 128350 618570 128420 618670
rect 128350 618530 128370 618570
rect 128410 618530 128420 618570
rect 128350 618480 128420 618530
rect 128140 618430 128420 618480
rect 128480 618620 128660 618670
rect 128480 618570 128550 618620
rect 128480 618530 128490 618570
rect 128530 618530 128550 618570
rect 128480 618480 128550 618530
rect 128580 618570 128660 618590
rect 128580 618530 128600 618570
rect 128640 618530 128660 618570
rect 128580 618510 128660 618530
rect 128690 618570 128760 618670
rect 128690 618530 128710 618570
rect 128750 618530 128760 618570
rect 128690 618480 128760 618530
rect 128480 618430 128760 618480
rect 128820 618620 129000 618670
rect 128820 618570 128890 618620
rect 128820 618530 128830 618570
rect 128870 618530 128890 618570
rect 128820 618480 128890 618530
rect 128920 618570 129000 618590
rect 128920 618530 128940 618570
rect 128980 618530 129000 618570
rect 128920 618510 129000 618530
rect 129030 618570 129100 618670
rect 129030 618530 129050 618570
rect 129090 618530 129100 618570
rect 129030 618480 129100 618530
rect 128820 618430 129100 618480
rect 129160 618620 129340 618670
rect 129160 618570 129230 618620
rect 129160 618530 129170 618570
rect 129210 618530 129230 618570
rect 129160 618480 129230 618530
rect 129260 618570 129340 618590
rect 129260 618530 129280 618570
rect 129320 618530 129340 618570
rect 129260 618510 129340 618530
rect 129370 618570 129440 618670
rect 129370 618530 129390 618570
rect 129430 618530 129440 618570
rect 129370 618480 129440 618530
rect 129160 618430 129440 618480
rect 129500 618620 129680 618670
rect 129500 618570 129570 618620
rect 129500 618530 129510 618570
rect 129550 618530 129570 618570
rect 129500 618480 129570 618530
rect 129600 618570 129680 618590
rect 129600 618530 129620 618570
rect 129660 618530 129680 618570
rect 129600 618510 129680 618530
rect 129710 618570 129780 618670
rect 129710 618530 129730 618570
rect 129770 618530 129780 618570
rect 129710 618480 129780 618530
rect 129500 618430 129780 618480
rect 129840 618620 130020 618670
rect 129840 618570 129910 618620
rect 129840 618530 129850 618570
rect 129890 618530 129910 618570
rect 129840 618480 129910 618530
rect 129940 618570 130020 618590
rect 129940 618530 129960 618570
rect 130000 618530 130020 618570
rect 129940 618510 130020 618530
rect 130050 618570 130120 618670
rect 130050 618530 130070 618570
rect 130110 618530 130120 618570
rect 130050 618480 130120 618530
rect 129840 618430 130120 618480
rect 130180 618620 130360 618670
rect 130180 618570 130250 618620
rect 130180 618530 130190 618570
rect 130230 618530 130250 618570
rect 130180 618480 130250 618530
rect 130280 618570 130360 618590
rect 130280 618530 130300 618570
rect 130340 618530 130360 618570
rect 130280 618510 130360 618530
rect 130390 618570 130460 618670
rect 130390 618530 130410 618570
rect 130450 618530 130460 618570
rect 130390 618480 130460 618530
rect 130180 618430 130460 618480
rect 130520 618620 130700 618670
rect 130520 618570 130590 618620
rect 130520 618530 130530 618570
rect 130570 618530 130590 618570
rect 130520 618480 130590 618530
rect 130620 618570 130700 618590
rect 130620 618530 130640 618570
rect 130680 618530 130700 618570
rect 130620 618510 130700 618530
rect 130730 618570 130800 618670
rect 130730 618530 130750 618570
rect 130790 618530 130800 618570
rect 130730 618480 130800 618530
rect 130520 618430 130800 618480
rect 130860 618620 131040 618670
rect 130860 618570 130930 618620
rect 130860 618530 130870 618570
rect 130910 618530 130930 618570
rect 130860 618480 130930 618530
rect 130960 618570 131040 618590
rect 130960 618530 130980 618570
rect 131020 618530 131040 618570
rect 130960 618510 131040 618530
rect 131070 618570 131140 618670
rect 131070 618530 131090 618570
rect 131130 618530 131140 618570
rect 131070 618480 131140 618530
rect 130860 618430 131140 618480
rect 131200 618620 131380 618670
rect 131200 618570 131270 618620
rect 131200 618530 131210 618570
rect 131250 618530 131270 618570
rect 131200 618480 131270 618530
rect 131300 618570 131380 618590
rect 131300 618530 131320 618570
rect 131360 618530 131380 618570
rect 131300 618510 131380 618530
rect 131410 618570 131480 618670
rect 131410 618530 131430 618570
rect 131470 618530 131480 618570
rect 131410 618480 131480 618530
rect 131200 618430 131480 618480
rect 131540 618620 131720 618670
rect 131540 618570 131610 618620
rect 131540 618530 131550 618570
rect 131590 618530 131610 618570
rect 131540 618480 131610 618530
rect 131640 618570 131720 618590
rect 131640 618530 131660 618570
rect 131700 618530 131720 618570
rect 131640 618510 131720 618530
rect 131750 618570 131820 618670
rect 131750 618530 131770 618570
rect 131810 618530 131820 618570
rect 131750 618480 131820 618530
rect 131540 618430 131820 618480
rect 125000 611950 125180 612000
rect 125000 611900 125070 611950
rect 125000 611860 125010 611900
rect 125050 611860 125070 611900
rect 125000 611810 125070 611860
rect 125100 611900 125180 611920
rect 125100 611860 125120 611900
rect 125160 611860 125180 611900
rect 125100 611840 125180 611860
rect 125210 611900 125280 612000
rect 125210 611860 125230 611900
rect 125270 611860 125280 611900
rect 125210 611810 125280 611860
rect 125000 611760 125280 611810
rect 125070 611170 125250 611220
rect 125070 611120 125140 611170
rect 125070 610930 125080 611120
rect 125120 610930 125140 611120
rect 125070 610880 125140 610930
rect 125170 611120 125250 611140
rect 125170 610930 125190 611120
rect 125230 610930 125250 611120
rect 125170 610910 125250 610930
rect 125280 611120 125350 611220
rect 125280 610930 125300 611120
rect 125340 610930 125350 611120
rect 125280 610880 125350 610930
rect 125070 610830 125350 610880
rect 125410 611170 125590 611220
rect 125410 611120 125480 611170
rect 125410 610930 125420 611120
rect 125460 610930 125480 611120
rect 125410 610880 125480 610930
rect 125510 611120 125590 611140
rect 125510 610930 125530 611120
rect 125570 610930 125590 611120
rect 125510 610910 125590 610930
rect 125620 611120 125690 611220
rect 125620 610930 125640 611120
rect 125680 610930 125690 611120
rect 125620 610880 125690 610930
rect 125410 610830 125690 610880
rect 125750 611170 125930 611220
rect 125750 611120 125820 611170
rect 125750 610930 125760 611120
rect 125800 610930 125820 611120
rect 125750 610880 125820 610930
rect 125850 611120 125930 611140
rect 125850 610930 125870 611120
rect 125910 610930 125930 611120
rect 125850 610910 125930 610930
rect 125960 611120 126030 611220
rect 125960 610930 125980 611120
rect 126020 610930 126030 611120
rect 125960 610880 126030 610930
rect 125750 610830 126030 610880
rect 126090 611170 126270 611220
rect 126090 611120 126160 611170
rect 126090 610930 126100 611120
rect 126140 610930 126160 611120
rect 126090 610880 126160 610930
rect 126190 611120 126270 611140
rect 126190 610930 126210 611120
rect 126250 610930 126270 611120
rect 126190 610910 126270 610930
rect 126300 611120 126370 611220
rect 126300 610930 126320 611120
rect 126360 610930 126370 611120
rect 126300 610880 126370 610930
rect 126090 610830 126370 610880
rect 126430 611170 126610 611220
rect 126430 611120 126500 611170
rect 126430 610930 126440 611120
rect 126480 610930 126500 611120
rect 126430 610880 126500 610930
rect 126530 611120 126610 611140
rect 126530 610930 126550 611120
rect 126590 610930 126610 611120
rect 126530 610910 126610 610930
rect 126640 611120 126710 611220
rect 126640 610930 126660 611120
rect 126700 610930 126710 611120
rect 126640 610880 126710 610930
rect 126430 610830 126710 610880
rect 126770 611170 126950 611220
rect 126770 611120 126840 611170
rect 126770 610930 126780 611120
rect 126820 610930 126840 611120
rect 126770 610880 126840 610930
rect 126870 611120 126950 611140
rect 126870 610930 126890 611120
rect 126930 610930 126950 611120
rect 126870 610910 126950 610930
rect 126980 611120 127050 611220
rect 126980 610930 127000 611120
rect 127040 610930 127050 611120
rect 126980 610880 127050 610930
rect 126770 610830 127050 610880
rect 127110 611170 127290 611220
rect 127110 611120 127180 611170
rect 127110 610930 127120 611120
rect 127160 610930 127180 611120
rect 127110 610880 127180 610930
rect 127210 611120 127290 611140
rect 127210 610930 127230 611120
rect 127270 610930 127290 611120
rect 127210 610910 127290 610930
rect 127320 611120 127390 611220
rect 127320 610930 127340 611120
rect 127380 610930 127390 611120
rect 127320 610880 127390 610930
rect 127110 610830 127390 610880
rect 127450 611170 127630 611220
rect 127450 611120 127520 611170
rect 127450 610930 127460 611120
rect 127500 610930 127520 611120
rect 127450 610880 127520 610930
rect 127550 611120 127630 611140
rect 127550 610930 127570 611120
rect 127610 610930 127630 611120
rect 127550 610910 127630 610930
rect 127660 611120 127730 611220
rect 127660 610930 127680 611120
rect 127720 610930 127730 611120
rect 127660 610880 127730 610930
rect 127450 610830 127730 610880
rect 127790 611170 127970 611220
rect 127790 611120 127860 611170
rect 127790 610930 127800 611120
rect 127840 610930 127860 611120
rect 127790 610880 127860 610930
rect 127890 611120 127970 611140
rect 127890 610930 127910 611120
rect 127950 610930 127970 611120
rect 127890 610910 127970 610930
rect 128000 611120 128070 611220
rect 128000 610930 128020 611120
rect 128060 610930 128070 611120
rect 128000 610880 128070 610930
rect 127790 610830 128070 610880
rect 128130 611170 128310 611220
rect 128130 611120 128200 611170
rect 128130 610930 128140 611120
rect 128180 610930 128200 611120
rect 128130 610880 128200 610930
rect 128230 611120 128310 611140
rect 128230 610930 128250 611120
rect 128290 610930 128310 611120
rect 128230 610910 128310 610930
rect 128340 611120 128410 611220
rect 128340 610930 128360 611120
rect 128400 610930 128410 611120
rect 128340 610880 128410 610930
rect 128130 610830 128410 610880
rect 128470 611170 128650 611220
rect 128470 611120 128540 611170
rect 128470 610930 128480 611120
rect 128520 610930 128540 611120
rect 128470 610880 128540 610930
rect 128570 611120 128650 611140
rect 128570 610930 128590 611120
rect 128630 610930 128650 611120
rect 128570 610910 128650 610930
rect 128680 611120 128750 611220
rect 128680 610930 128700 611120
rect 128740 610930 128750 611120
rect 128680 610880 128750 610930
rect 128470 610830 128750 610880
rect 128810 611170 128990 611220
rect 128810 611120 128880 611170
rect 128810 610930 128820 611120
rect 128860 610930 128880 611120
rect 128810 610880 128880 610930
rect 128910 611120 128990 611140
rect 128910 610930 128930 611120
rect 128970 610930 128990 611120
rect 128910 610910 128990 610930
rect 129020 611120 129090 611220
rect 129020 610930 129040 611120
rect 129080 610930 129090 611120
rect 129020 610880 129090 610930
rect 128810 610830 129090 610880
rect 129150 611170 129330 611220
rect 129150 611120 129220 611170
rect 129150 610930 129160 611120
rect 129200 610930 129220 611120
rect 129150 610880 129220 610930
rect 129250 611120 129330 611140
rect 129250 610930 129270 611120
rect 129310 610930 129330 611120
rect 129250 610910 129330 610930
rect 129360 611120 129430 611220
rect 129360 610930 129380 611120
rect 129420 610930 129430 611120
rect 129360 610880 129430 610930
rect 129150 610830 129430 610880
rect 129490 611170 129670 611220
rect 129490 611120 129560 611170
rect 129490 610930 129500 611120
rect 129540 610930 129560 611120
rect 129490 610880 129560 610930
rect 129590 611120 129670 611140
rect 129590 610930 129610 611120
rect 129650 610930 129670 611120
rect 129590 610910 129670 610930
rect 129700 611120 129770 611220
rect 129700 610930 129720 611120
rect 129760 610930 129770 611120
rect 129700 610880 129770 610930
rect 129490 610830 129770 610880
rect 129830 611170 130010 611220
rect 129830 611120 129900 611170
rect 129830 610930 129840 611120
rect 129880 610930 129900 611120
rect 129830 610880 129900 610930
rect 129930 611120 130010 611140
rect 129930 610930 129950 611120
rect 129990 610930 130010 611120
rect 129930 610910 130010 610930
rect 130040 611120 130110 611220
rect 130040 610930 130060 611120
rect 130100 610930 130110 611120
rect 130040 610880 130110 610930
rect 129830 610830 130110 610880
rect 130170 611170 130350 611220
rect 130170 611120 130240 611170
rect 130170 610930 130180 611120
rect 130220 610930 130240 611120
rect 130170 610880 130240 610930
rect 130270 611120 130350 611140
rect 130270 610930 130290 611120
rect 130330 610930 130350 611120
rect 130270 610910 130350 610930
rect 130380 611120 130450 611220
rect 130380 610930 130400 611120
rect 130440 610930 130450 611120
rect 130380 610880 130450 610930
rect 130170 610830 130450 610880
rect 130510 611170 130690 611220
rect 130510 611120 130580 611170
rect 130510 610930 130520 611120
rect 130560 610930 130580 611120
rect 130510 610880 130580 610930
rect 130610 611120 130690 611140
rect 130610 610930 130630 611120
rect 130670 610930 130690 611120
rect 130610 610910 130690 610930
rect 130720 611120 130790 611220
rect 130720 610930 130740 611120
rect 130780 610930 130790 611120
rect 130720 610880 130790 610930
rect 130510 610830 130790 610880
rect 130850 611170 131030 611220
rect 130850 611120 130920 611170
rect 130850 610930 130860 611120
rect 130900 610930 130920 611120
rect 130850 610880 130920 610930
rect 130950 611120 131030 611140
rect 130950 610930 130970 611120
rect 131010 610930 131030 611120
rect 130950 610910 131030 610930
rect 131060 611120 131130 611220
rect 131060 610930 131080 611120
rect 131120 610930 131130 611120
rect 131060 610880 131130 610930
rect 130850 610830 131130 610880
rect 131190 611170 131370 611220
rect 131190 611120 131260 611170
rect 131190 610930 131200 611120
rect 131240 610930 131260 611120
rect 131190 610880 131260 610930
rect 131290 611120 131370 611140
rect 131290 610930 131310 611120
rect 131350 610930 131370 611120
rect 131290 610910 131370 610930
rect 131400 611120 131470 611220
rect 131400 610930 131420 611120
rect 131460 610930 131470 611120
rect 131400 610880 131470 610930
rect 131190 610830 131470 610880
rect 125130 605900 125310 605950
rect 125130 605850 125200 605900
rect 125130 605810 125140 605850
rect 125180 605810 125200 605850
rect 125130 605760 125200 605810
rect 125230 605850 125310 605870
rect 125230 605810 125250 605850
rect 125290 605810 125310 605850
rect 125230 605790 125310 605810
rect 125340 605850 125410 605950
rect 125340 605810 125360 605850
rect 125400 605810 125410 605850
rect 125340 605760 125410 605810
rect 125130 605710 125410 605760
rect 125200 605120 125380 605170
rect 125200 605070 125270 605120
rect 125200 604780 125210 605070
rect 125250 604780 125270 605070
rect 125200 604730 125270 604780
rect 125300 605070 125380 605090
rect 125300 604780 125320 605070
rect 125360 604780 125380 605070
rect 125300 604760 125380 604780
rect 125410 605070 125480 605170
rect 125410 604780 125430 605070
rect 125470 604780 125480 605070
rect 125410 604730 125480 604780
rect 125200 604680 125480 604730
rect 125540 605120 125720 605170
rect 125540 605070 125610 605120
rect 125540 604780 125550 605070
rect 125590 604780 125610 605070
rect 125540 604730 125610 604780
rect 125640 605070 125720 605090
rect 125640 604780 125660 605070
rect 125700 604780 125720 605070
rect 125640 604760 125720 604780
rect 125750 605070 125820 605170
rect 125750 604780 125770 605070
rect 125810 604780 125820 605070
rect 125750 604730 125820 604780
rect 125540 604680 125820 604730
rect 125880 605120 126060 605170
rect 125880 605070 125950 605120
rect 125880 604780 125890 605070
rect 125930 604780 125950 605070
rect 125880 604730 125950 604780
rect 125980 605070 126060 605090
rect 125980 604780 126000 605070
rect 126040 604780 126060 605070
rect 125980 604760 126060 604780
rect 126090 605070 126160 605170
rect 126090 604780 126110 605070
rect 126150 604780 126160 605070
rect 126090 604730 126160 604780
rect 125880 604680 126160 604730
rect 126220 605120 126400 605170
rect 126220 605070 126290 605120
rect 126220 604780 126230 605070
rect 126270 604780 126290 605070
rect 126220 604730 126290 604780
rect 126320 605070 126400 605090
rect 126320 604780 126340 605070
rect 126380 604780 126400 605070
rect 126320 604760 126400 604780
rect 126430 605070 126500 605170
rect 126430 604780 126450 605070
rect 126490 604780 126500 605070
rect 126430 604730 126500 604780
rect 126220 604680 126500 604730
rect 126560 605120 126740 605170
rect 126560 605070 126630 605120
rect 126560 604780 126570 605070
rect 126610 604780 126630 605070
rect 126560 604730 126630 604780
rect 126660 605070 126740 605090
rect 126660 604780 126680 605070
rect 126720 604780 126740 605070
rect 126660 604760 126740 604780
rect 126770 605070 126840 605170
rect 126770 604780 126790 605070
rect 126830 604780 126840 605070
rect 126770 604730 126840 604780
rect 126560 604680 126840 604730
rect 126900 605120 127080 605170
rect 126900 605070 126970 605120
rect 126900 604780 126910 605070
rect 126950 604780 126970 605070
rect 126900 604730 126970 604780
rect 127000 605070 127080 605090
rect 127000 604780 127020 605070
rect 127060 604780 127080 605070
rect 127000 604760 127080 604780
rect 127110 605070 127180 605170
rect 127110 604780 127130 605070
rect 127170 604780 127180 605070
rect 127110 604730 127180 604780
rect 126900 604680 127180 604730
rect 127240 605120 127420 605170
rect 127240 605070 127310 605120
rect 127240 604780 127250 605070
rect 127290 604780 127310 605070
rect 127240 604730 127310 604780
rect 127340 605070 127420 605090
rect 127340 604780 127360 605070
rect 127400 604780 127420 605070
rect 127340 604760 127420 604780
rect 127450 605070 127520 605170
rect 127450 604780 127470 605070
rect 127510 604780 127520 605070
rect 127450 604730 127520 604780
rect 127240 604680 127520 604730
rect 127580 605120 127760 605170
rect 127580 605070 127650 605120
rect 127580 604780 127590 605070
rect 127630 604780 127650 605070
rect 127580 604730 127650 604780
rect 127680 605070 127760 605090
rect 127680 604780 127700 605070
rect 127740 604780 127760 605070
rect 127680 604760 127760 604780
rect 127790 605070 127860 605170
rect 127790 604780 127810 605070
rect 127850 604780 127860 605070
rect 127790 604730 127860 604780
rect 127580 604680 127860 604730
rect 127920 605120 128100 605170
rect 127920 605070 127990 605120
rect 127920 604780 127930 605070
rect 127970 604780 127990 605070
rect 127920 604730 127990 604780
rect 128020 605070 128100 605090
rect 128020 604780 128040 605070
rect 128080 604780 128100 605070
rect 128020 604760 128100 604780
rect 128130 605070 128200 605170
rect 128130 604780 128150 605070
rect 128190 604780 128200 605070
rect 128130 604730 128200 604780
rect 127920 604680 128200 604730
rect 128260 605120 128440 605170
rect 128260 605070 128330 605120
rect 128260 604780 128270 605070
rect 128310 604780 128330 605070
rect 128260 604730 128330 604780
rect 128360 605070 128440 605090
rect 128360 604780 128380 605070
rect 128420 604780 128440 605070
rect 128360 604760 128440 604780
rect 128470 605070 128540 605170
rect 128470 604780 128490 605070
rect 128530 604780 128540 605070
rect 128470 604730 128540 604780
rect 128260 604680 128540 604730
rect 128600 605120 128780 605170
rect 128600 605070 128670 605120
rect 128600 604780 128610 605070
rect 128650 604780 128670 605070
rect 128600 604730 128670 604780
rect 128700 605070 128780 605090
rect 128700 604780 128720 605070
rect 128760 604780 128780 605070
rect 128700 604760 128780 604780
rect 128810 605070 128880 605170
rect 128810 604780 128830 605070
rect 128870 604780 128880 605070
rect 128810 604730 128880 604780
rect 128600 604680 128880 604730
rect 128940 605120 129120 605170
rect 128940 605070 129010 605120
rect 128940 604780 128950 605070
rect 128990 604780 129010 605070
rect 128940 604730 129010 604780
rect 129040 605070 129120 605090
rect 129040 604780 129060 605070
rect 129100 604780 129120 605070
rect 129040 604760 129120 604780
rect 129150 605070 129220 605170
rect 129150 604780 129170 605070
rect 129210 604780 129220 605070
rect 129150 604730 129220 604780
rect 128940 604680 129220 604730
rect 129280 605120 129460 605170
rect 129280 605070 129350 605120
rect 129280 604780 129290 605070
rect 129330 604780 129350 605070
rect 129280 604730 129350 604780
rect 129380 605070 129460 605090
rect 129380 604780 129400 605070
rect 129440 604780 129460 605070
rect 129380 604760 129460 604780
rect 129490 605070 129560 605170
rect 129490 604780 129510 605070
rect 129550 604780 129560 605070
rect 129490 604730 129560 604780
rect 129280 604680 129560 604730
rect 129620 605120 129800 605170
rect 129620 605070 129690 605120
rect 129620 604780 129630 605070
rect 129670 604780 129690 605070
rect 129620 604730 129690 604780
rect 129720 605070 129800 605090
rect 129720 604780 129740 605070
rect 129780 604780 129800 605070
rect 129720 604760 129800 604780
rect 129830 605070 129900 605170
rect 129830 604780 129850 605070
rect 129890 604780 129900 605070
rect 129830 604730 129900 604780
rect 129620 604680 129900 604730
rect 129960 605120 130140 605170
rect 129960 605070 130030 605120
rect 129960 604780 129970 605070
rect 130010 604780 130030 605070
rect 129960 604730 130030 604780
rect 130060 605070 130140 605090
rect 130060 604780 130080 605070
rect 130120 604780 130140 605070
rect 130060 604760 130140 604780
rect 130170 605070 130240 605170
rect 130170 604780 130190 605070
rect 130230 604780 130240 605070
rect 130170 604730 130240 604780
rect 129960 604680 130240 604730
rect 130300 605120 130480 605170
rect 130300 605070 130370 605120
rect 130300 604780 130310 605070
rect 130350 604780 130370 605070
rect 130300 604730 130370 604780
rect 130400 605070 130480 605090
rect 130400 604780 130420 605070
rect 130460 604780 130480 605070
rect 130400 604760 130480 604780
rect 130510 605070 130580 605170
rect 130510 604780 130530 605070
rect 130570 604780 130580 605070
rect 130510 604730 130580 604780
rect 130300 604680 130580 604730
rect 130640 605120 130820 605170
rect 130640 605070 130710 605120
rect 130640 604780 130650 605070
rect 130690 604780 130710 605070
rect 130640 604730 130710 604780
rect 130740 605070 130820 605090
rect 130740 604780 130760 605070
rect 130800 604780 130820 605070
rect 130740 604760 130820 604780
rect 130850 605070 130920 605170
rect 130850 604780 130870 605070
rect 130910 604780 130920 605070
rect 130850 604730 130920 604780
rect 130640 604680 130920 604730
rect 130980 605120 131160 605170
rect 130980 605070 131050 605120
rect 130980 604780 130990 605070
rect 131030 604780 131050 605070
rect 130980 604730 131050 604780
rect 131080 605070 131160 605090
rect 131080 604780 131100 605070
rect 131140 604780 131160 605070
rect 131080 604760 131160 604780
rect 131190 605070 131260 605170
rect 131190 604780 131210 605070
rect 131250 604780 131260 605070
rect 131190 604730 131260 604780
rect 130980 604680 131260 604730
rect 131320 605120 131500 605170
rect 131320 605070 131390 605120
rect 131320 604780 131330 605070
rect 131370 604780 131390 605070
rect 131320 604730 131390 604780
rect 131420 605070 131500 605090
rect 131420 604780 131440 605070
rect 131480 604780 131500 605070
rect 131420 604760 131500 604780
rect 131530 605070 131600 605170
rect 131530 604780 131550 605070
rect 131590 604780 131600 605070
rect 131530 604730 131600 604780
rect 131320 604680 131600 604730
rect 124930 599640 125110 599690
rect 124930 599590 125000 599640
rect 124930 599550 124940 599590
rect 124980 599550 125000 599590
rect 124930 599500 125000 599550
rect 125030 599590 125110 599610
rect 125030 599550 125050 599590
rect 125090 599550 125110 599590
rect 125030 599530 125110 599550
rect 125140 599590 125210 599690
rect 125140 599550 125160 599590
rect 125200 599550 125210 599590
rect 125140 599500 125210 599550
rect 124930 599450 125210 599500
rect 125000 598860 125180 598910
rect 125000 598810 125070 598860
rect 125000 598420 125010 598810
rect 125050 598420 125070 598810
rect 125000 598370 125070 598420
rect 125100 598810 125180 598830
rect 125100 598420 125120 598810
rect 125160 598420 125180 598810
rect 125100 598400 125180 598420
rect 125210 598810 125280 598910
rect 125210 598420 125230 598810
rect 125270 598420 125280 598810
rect 125210 598370 125280 598420
rect 125000 598320 125280 598370
rect 125340 598860 125520 598910
rect 125340 598810 125410 598860
rect 125340 598420 125350 598810
rect 125390 598420 125410 598810
rect 125340 598370 125410 598420
rect 125440 598810 125520 598830
rect 125440 598420 125460 598810
rect 125500 598420 125520 598810
rect 125440 598400 125520 598420
rect 125550 598810 125620 598910
rect 125550 598420 125570 598810
rect 125610 598420 125620 598810
rect 125550 598370 125620 598420
rect 125340 598320 125620 598370
rect 125680 598860 125860 598910
rect 125680 598810 125750 598860
rect 125680 598420 125690 598810
rect 125730 598420 125750 598810
rect 125680 598370 125750 598420
rect 125780 598810 125860 598830
rect 125780 598420 125800 598810
rect 125840 598420 125860 598810
rect 125780 598400 125860 598420
rect 125890 598810 125960 598910
rect 125890 598420 125910 598810
rect 125950 598420 125960 598810
rect 125890 598370 125960 598420
rect 125680 598320 125960 598370
rect 126020 598860 126200 598910
rect 126020 598810 126090 598860
rect 126020 598420 126030 598810
rect 126070 598420 126090 598810
rect 126020 598370 126090 598420
rect 126120 598810 126200 598830
rect 126120 598420 126140 598810
rect 126180 598420 126200 598810
rect 126120 598400 126200 598420
rect 126230 598810 126300 598910
rect 126230 598420 126250 598810
rect 126290 598420 126300 598810
rect 126230 598370 126300 598420
rect 126020 598320 126300 598370
rect 126360 598860 126540 598910
rect 126360 598810 126430 598860
rect 126360 598420 126370 598810
rect 126410 598420 126430 598810
rect 126360 598370 126430 598420
rect 126460 598810 126540 598830
rect 126460 598420 126480 598810
rect 126520 598420 126540 598810
rect 126460 598400 126540 598420
rect 126570 598810 126640 598910
rect 126570 598420 126590 598810
rect 126630 598420 126640 598810
rect 126570 598370 126640 598420
rect 126360 598320 126640 598370
rect 126700 598860 126880 598910
rect 126700 598810 126770 598860
rect 126700 598420 126710 598810
rect 126750 598420 126770 598810
rect 126700 598370 126770 598420
rect 126800 598810 126880 598830
rect 126800 598420 126820 598810
rect 126860 598420 126880 598810
rect 126800 598400 126880 598420
rect 126910 598810 126980 598910
rect 126910 598420 126930 598810
rect 126970 598420 126980 598810
rect 126910 598370 126980 598420
rect 126700 598320 126980 598370
rect 127040 598860 127220 598910
rect 127040 598810 127110 598860
rect 127040 598420 127050 598810
rect 127090 598420 127110 598810
rect 127040 598370 127110 598420
rect 127140 598810 127220 598830
rect 127140 598420 127160 598810
rect 127200 598420 127220 598810
rect 127140 598400 127220 598420
rect 127250 598810 127320 598910
rect 127250 598420 127270 598810
rect 127310 598420 127320 598810
rect 127250 598370 127320 598420
rect 127040 598320 127320 598370
rect 127380 598860 127560 598910
rect 127380 598810 127450 598860
rect 127380 598420 127390 598810
rect 127430 598420 127450 598810
rect 127380 598370 127450 598420
rect 127480 598810 127560 598830
rect 127480 598420 127500 598810
rect 127540 598420 127560 598810
rect 127480 598400 127560 598420
rect 127590 598810 127660 598910
rect 127590 598420 127610 598810
rect 127650 598420 127660 598810
rect 127590 598370 127660 598420
rect 127380 598320 127660 598370
rect 127720 598860 127900 598910
rect 127720 598810 127790 598860
rect 127720 598420 127730 598810
rect 127770 598420 127790 598810
rect 127720 598370 127790 598420
rect 127820 598810 127900 598830
rect 127820 598420 127840 598810
rect 127880 598420 127900 598810
rect 127820 598400 127900 598420
rect 127930 598810 128000 598910
rect 127930 598420 127950 598810
rect 127990 598420 128000 598810
rect 127930 598370 128000 598420
rect 127720 598320 128000 598370
rect 128060 598860 128240 598910
rect 128060 598810 128130 598860
rect 128060 598420 128070 598810
rect 128110 598420 128130 598810
rect 128060 598370 128130 598420
rect 128160 598810 128240 598830
rect 128160 598420 128180 598810
rect 128220 598420 128240 598810
rect 128160 598400 128240 598420
rect 128270 598810 128340 598910
rect 128270 598420 128290 598810
rect 128330 598420 128340 598810
rect 128270 598370 128340 598420
rect 128060 598320 128340 598370
rect 128400 598860 128580 598910
rect 128400 598810 128470 598860
rect 128400 598420 128410 598810
rect 128450 598420 128470 598810
rect 128400 598370 128470 598420
rect 128500 598810 128580 598830
rect 128500 598420 128520 598810
rect 128560 598420 128580 598810
rect 128500 598400 128580 598420
rect 128610 598810 128680 598910
rect 128610 598420 128630 598810
rect 128670 598420 128680 598810
rect 128610 598370 128680 598420
rect 128400 598320 128680 598370
rect 128740 598860 128920 598910
rect 128740 598810 128810 598860
rect 128740 598420 128750 598810
rect 128790 598420 128810 598810
rect 128740 598370 128810 598420
rect 128840 598810 128920 598830
rect 128840 598420 128860 598810
rect 128900 598420 128920 598810
rect 128840 598400 128920 598420
rect 128950 598810 129020 598910
rect 128950 598420 128970 598810
rect 129010 598420 129020 598810
rect 128950 598370 129020 598420
rect 128740 598320 129020 598370
rect 129080 598860 129260 598910
rect 129080 598810 129150 598860
rect 129080 598420 129090 598810
rect 129130 598420 129150 598810
rect 129080 598370 129150 598420
rect 129180 598810 129260 598830
rect 129180 598420 129200 598810
rect 129240 598420 129260 598810
rect 129180 598400 129260 598420
rect 129290 598810 129360 598910
rect 129290 598420 129310 598810
rect 129350 598420 129360 598810
rect 129290 598370 129360 598420
rect 129080 598320 129360 598370
rect 129420 598860 129600 598910
rect 129420 598810 129490 598860
rect 129420 598420 129430 598810
rect 129470 598420 129490 598810
rect 129420 598370 129490 598420
rect 129520 598810 129600 598830
rect 129520 598420 129540 598810
rect 129580 598420 129600 598810
rect 129520 598400 129600 598420
rect 129630 598810 129700 598910
rect 129630 598420 129650 598810
rect 129690 598420 129700 598810
rect 129630 598370 129700 598420
rect 129420 598320 129700 598370
rect 129760 598860 129940 598910
rect 129760 598810 129830 598860
rect 129760 598420 129770 598810
rect 129810 598420 129830 598810
rect 129760 598370 129830 598420
rect 129860 598810 129940 598830
rect 129860 598420 129880 598810
rect 129920 598420 129940 598810
rect 129860 598400 129940 598420
rect 129970 598810 130040 598910
rect 129970 598420 129990 598810
rect 130030 598420 130040 598810
rect 129970 598370 130040 598420
rect 129760 598320 130040 598370
rect 130100 598860 130280 598910
rect 130100 598810 130170 598860
rect 130100 598420 130110 598810
rect 130150 598420 130170 598810
rect 130100 598370 130170 598420
rect 130200 598810 130280 598830
rect 130200 598420 130220 598810
rect 130260 598420 130280 598810
rect 130200 598400 130280 598420
rect 130310 598810 130380 598910
rect 130310 598420 130330 598810
rect 130370 598420 130380 598810
rect 130310 598370 130380 598420
rect 130100 598320 130380 598370
rect 130440 598860 130620 598910
rect 130440 598810 130510 598860
rect 130440 598420 130450 598810
rect 130490 598420 130510 598810
rect 130440 598370 130510 598420
rect 130540 598810 130620 598830
rect 130540 598420 130560 598810
rect 130600 598420 130620 598810
rect 130540 598400 130620 598420
rect 130650 598810 130720 598910
rect 130650 598420 130670 598810
rect 130710 598420 130720 598810
rect 130650 598370 130720 598420
rect 130440 598320 130720 598370
rect 130780 598860 130960 598910
rect 130780 598810 130850 598860
rect 130780 598420 130790 598810
rect 130830 598420 130850 598810
rect 130780 598370 130850 598420
rect 130880 598810 130960 598830
rect 130880 598420 130900 598810
rect 130940 598420 130960 598810
rect 130880 598400 130960 598420
rect 130990 598810 131060 598910
rect 130990 598420 131010 598810
rect 131050 598420 131060 598810
rect 130990 598370 131060 598420
rect 130780 598320 131060 598370
rect 131120 598860 131300 598910
rect 131120 598810 131190 598860
rect 131120 598420 131130 598810
rect 131170 598420 131190 598810
rect 131120 598370 131190 598420
rect 131220 598810 131300 598830
rect 131220 598420 131240 598810
rect 131280 598420 131300 598810
rect 131220 598400 131300 598420
rect 131330 598810 131400 598910
rect 131330 598420 131350 598810
rect 131390 598420 131400 598810
rect 131330 598370 131400 598420
rect 131120 598320 131400 598370
rect 119260 592950 119330 592970
rect 119260 592900 119270 592950
rect 119310 592900 119330 592950
rect 119260 592880 119330 592900
rect 119360 592950 119430 592970
rect 119360 592900 119380 592950
rect 119420 592900 119430 592950
rect 119360 592880 119430 592900
rect 119620 592750 119690 592770
rect 119620 592590 119630 592750
rect 119670 592590 119690 592750
rect 119620 592570 119690 592590
rect 119720 592750 119790 592770
rect 119720 592590 119740 592750
rect 119780 592590 119790 592750
rect 119720 592570 119790 592590
rect 120000 592750 120070 592770
rect 120000 592590 120010 592750
rect 120050 592590 120070 592750
rect 120000 592570 120070 592590
rect 120100 592750 120170 592770
rect 120100 592590 120120 592750
rect 120160 592590 120170 592750
rect 120100 592570 120170 592590
rect 124890 592090 125070 592140
rect 124890 592040 124960 592090
rect 124890 592000 124900 592040
rect 124940 592000 124960 592040
rect 124890 591950 124960 592000
rect 124990 592040 125070 592060
rect 124990 592000 125010 592040
rect 125050 592000 125070 592040
rect 124990 591980 125070 592000
rect 125100 592040 125170 592140
rect 125100 592000 125120 592040
rect 125160 592000 125170 592040
rect 125100 591950 125170 592000
rect 124890 591900 125170 591950
rect 124960 591310 125140 591360
rect 124960 591260 125030 591310
rect 124960 590770 124970 591260
rect 125010 590770 125030 591260
rect 124960 590720 125030 590770
rect 125060 591260 125140 591280
rect 125060 590770 125080 591260
rect 125120 590770 125140 591260
rect 125060 590750 125140 590770
rect 125170 591260 125240 591360
rect 125170 590770 125190 591260
rect 125230 590770 125240 591260
rect 125170 590720 125240 590770
rect 124960 590670 125240 590720
rect 125300 591310 125480 591360
rect 125300 591260 125370 591310
rect 125300 590770 125310 591260
rect 125350 590770 125370 591260
rect 125300 590720 125370 590770
rect 125400 591260 125480 591280
rect 125400 590770 125420 591260
rect 125460 590770 125480 591260
rect 125400 590750 125480 590770
rect 125510 591260 125580 591360
rect 125510 590770 125530 591260
rect 125570 590770 125580 591260
rect 125510 590720 125580 590770
rect 125300 590670 125580 590720
rect 125640 591310 125820 591360
rect 125640 591260 125710 591310
rect 125640 590770 125650 591260
rect 125690 590770 125710 591260
rect 125640 590720 125710 590770
rect 125740 591260 125820 591280
rect 125740 590770 125760 591260
rect 125800 590770 125820 591260
rect 125740 590750 125820 590770
rect 125850 591260 125920 591360
rect 125850 590770 125870 591260
rect 125910 590770 125920 591260
rect 125850 590720 125920 590770
rect 125640 590670 125920 590720
rect 125980 591310 126160 591360
rect 125980 591260 126050 591310
rect 125980 590770 125990 591260
rect 126030 590770 126050 591260
rect 125980 590720 126050 590770
rect 126080 591260 126160 591280
rect 126080 590770 126100 591260
rect 126140 590770 126160 591260
rect 126080 590750 126160 590770
rect 126190 591260 126260 591360
rect 126190 590770 126210 591260
rect 126250 590770 126260 591260
rect 126190 590720 126260 590770
rect 125980 590670 126260 590720
rect 126320 591310 126500 591360
rect 126320 591260 126390 591310
rect 126320 590770 126330 591260
rect 126370 590770 126390 591260
rect 126320 590720 126390 590770
rect 126420 591260 126500 591280
rect 126420 590770 126440 591260
rect 126480 590770 126500 591260
rect 126420 590750 126500 590770
rect 126530 591260 126600 591360
rect 126530 590770 126550 591260
rect 126590 590770 126600 591260
rect 126530 590720 126600 590770
rect 126320 590670 126600 590720
rect 126660 591310 126840 591360
rect 126660 591260 126730 591310
rect 126660 590770 126670 591260
rect 126710 590770 126730 591260
rect 126660 590720 126730 590770
rect 126760 591260 126840 591280
rect 126760 590770 126780 591260
rect 126820 590770 126840 591260
rect 126760 590750 126840 590770
rect 126870 591260 126940 591360
rect 126870 590770 126890 591260
rect 126930 590770 126940 591260
rect 126870 590720 126940 590770
rect 126660 590670 126940 590720
rect 127000 591310 127180 591360
rect 127000 591260 127070 591310
rect 127000 590770 127010 591260
rect 127050 590770 127070 591260
rect 127000 590720 127070 590770
rect 127100 591260 127180 591280
rect 127100 590770 127120 591260
rect 127160 590770 127180 591260
rect 127100 590750 127180 590770
rect 127210 591260 127280 591360
rect 127210 590770 127230 591260
rect 127270 590770 127280 591260
rect 127210 590720 127280 590770
rect 127000 590670 127280 590720
rect 127340 591310 127520 591360
rect 127340 591260 127410 591310
rect 127340 590770 127350 591260
rect 127390 590770 127410 591260
rect 127340 590720 127410 590770
rect 127440 591260 127520 591280
rect 127440 590770 127460 591260
rect 127500 590770 127520 591260
rect 127440 590750 127520 590770
rect 127550 591260 127620 591360
rect 127550 590770 127570 591260
rect 127610 590770 127620 591260
rect 127550 590720 127620 590770
rect 127340 590670 127620 590720
rect 127680 591310 127860 591360
rect 127680 591260 127750 591310
rect 127680 590770 127690 591260
rect 127730 590770 127750 591260
rect 127680 590720 127750 590770
rect 127780 591260 127860 591280
rect 127780 590770 127800 591260
rect 127840 590770 127860 591260
rect 127780 590750 127860 590770
rect 127890 591260 127960 591360
rect 127890 590770 127910 591260
rect 127950 590770 127960 591260
rect 127890 590720 127960 590770
rect 127680 590670 127960 590720
rect 128020 591310 128200 591360
rect 128020 591260 128090 591310
rect 128020 590770 128030 591260
rect 128070 590770 128090 591260
rect 128020 590720 128090 590770
rect 128120 591260 128200 591280
rect 128120 590770 128140 591260
rect 128180 590770 128200 591260
rect 128120 590750 128200 590770
rect 128230 591260 128300 591360
rect 128230 590770 128250 591260
rect 128290 590770 128300 591260
rect 128230 590720 128300 590770
rect 128020 590670 128300 590720
rect 128360 591310 128540 591360
rect 128360 591260 128430 591310
rect 128360 590770 128370 591260
rect 128410 590770 128430 591260
rect 128360 590720 128430 590770
rect 128460 591260 128540 591280
rect 128460 590770 128480 591260
rect 128520 590770 128540 591260
rect 128460 590750 128540 590770
rect 128570 591260 128640 591360
rect 128570 590770 128590 591260
rect 128630 590770 128640 591260
rect 128570 590720 128640 590770
rect 128360 590670 128640 590720
rect 128700 591310 128880 591360
rect 128700 591260 128770 591310
rect 128700 590770 128710 591260
rect 128750 590770 128770 591260
rect 128700 590720 128770 590770
rect 128800 591260 128880 591280
rect 128800 590770 128820 591260
rect 128860 590770 128880 591260
rect 128800 590750 128880 590770
rect 128910 591260 128980 591360
rect 128910 590770 128930 591260
rect 128970 590770 128980 591260
rect 128910 590720 128980 590770
rect 128700 590670 128980 590720
rect 129040 591310 129220 591360
rect 129040 591260 129110 591310
rect 129040 590770 129050 591260
rect 129090 590770 129110 591260
rect 129040 590720 129110 590770
rect 129140 591260 129220 591280
rect 129140 590770 129160 591260
rect 129200 590770 129220 591260
rect 129140 590750 129220 590770
rect 129250 591260 129320 591360
rect 129250 590770 129270 591260
rect 129310 590770 129320 591260
rect 129250 590720 129320 590770
rect 129040 590670 129320 590720
rect 129380 591310 129560 591360
rect 129380 591260 129450 591310
rect 129380 590770 129390 591260
rect 129430 590770 129450 591260
rect 129380 590720 129450 590770
rect 129480 591260 129560 591280
rect 129480 590770 129500 591260
rect 129540 590770 129560 591260
rect 129480 590750 129560 590770
rect 129590 591260 129660 591360
rect 129590 590770 129610 591260
rect 129650 590770 129660 591260
rect 129590 590720 129660 590770
rect 129380 590670 129660 590720
rect 129720 591310 129900 591360
rect 129720 591260 129790 591310
rect 129720 590770 129730 591260
rect 129770 590770 129790 591260
rect 129720 590720 129790 590770
rect 129820 591260 129900 591280
rect 129820 590770 129840 591260
rect 129880 590770 129900 591260
rect 129820 590750 129900 590770
rect 129930 591260 130000 591360
rect 129930 590770 129950 591260
rect 129990 590770 130000 591260
rect 129930 590720 130000 590770
rect 129720 590670 130000 590720
rect 130060 591310 130240 591360
rect 130060 591260 130130 591310
rect 130060 590770 130070 591260
rect 130110 590770 130130 591260
rect 130060 590720 130130 590770
rect 130160 591260 130240 591280
rect 130160 590770 130180 591260
rect 130220 590770 130240 591260
rect 130160 590750 130240 590770
rect 130270 591260 130340 591360
rect 130270 590770 130290 591260
rect 130330 590770 130340 591260
rect 130270 590720 130340 590770
rect 130060 590670 130340 590720
rect 130400 591310 130580 591360
rect 130400 591260 130470 591310
rect 130400 590770 130410 591260
rect 130450 590770 130470 591260
rect 130400 590720 130470 590770
rect 130500 591260 130580 591280
rect 130500 590770 130520 591260
rect 130560 590770 130580 591260
rect 130500 590750 130580 590770
rect 130610 591260 130680 591360
rect 130610 590770 130630 591260
rect 130670 590770 130680 591260
rect 130610 590720 130680 590770
rect 130400 590670 130680 590720
rect 130740 591310 130920 591360
rect 130740 591260 130810 591310
rect 130740 590770 130750 591260
rect 130790 590770 130810 591260
rect 130740 590720 130810 590770
rect 130840 591260 130920 591280
rect 130840 590770 130860 591260
rect 130900 590770 130920 591260
rect 130840 590750 130920 590770
rect 130950 591260 131020 591360
rect 130950 590770 130970 591260
rect 131010 590770 131020 591260
rect 130950 590720 131020 590770
rect 130740 590670 131020 590720
rect 131080 591310 131260 591360
rect 131080 591260 131150 591310
rect 131080 590770 131090 591260
rect 131130 590770 131150 591260
rect 131080 590720 131150 590770
rect 131180 591260 131260 591280
rect 131180 590770 131200 591260
rect 131240 590770 131260 591260
rect 131180 590750 131260 590770
rect 131290 591260 131360 591360
rect 131290 590770 131310 591260
rect 131350 590770 131360 591260
rect 131290 590720 131360 590770
rect 131080 590670 131360 590720
rect 119300 583410 119370 583430
rect 119300 583360 119310 583410
rect 119350 583360 119370 583410
rect 119300 583340 119370 583360
rect 119400 583410 119470 583430
rect 119400 583360 119420 583410
rect 119460 583360 119470 583410
rect 119400 583340 119470 583360
rect 119660 583210 119730 583230
rect 119660 583050 119670 583210
rect 119710 583050 119730 583210
rect 119660 583030 119730 583050
rect 119760 583210 119830 583230
rect 119760 583050 119780 583210
rect 119820 583050 119830 583210
rect 119760 583030 119830 583050
rect 120040 583210 120110 583230
rect 120040 583050 120050 583210
rect 120090 583050 120110 583210
rect 120040 583030 120110 583050
rect 120140 583210 120210 583230
rect 120140 583050 120160 583210
rect 120200 583050 120210 583210
rect 120140 583030 120210 583050
rect 125350 583110 125530 583160
rect 125350 583060 125420 583110
rect 125350 583020 125360 583060
rect 125400 583020 125420 583060
rect 125350 582970 125420 583020
rect 125450 583060 125530 583080
rect 125450 583020 125470 583060
rect 125510 583020 125530 583060
rect 125450 583000 125530 583020
rect 125560 583060 125630 583160
rect 125560 583020 125580 583060
rect 125620 583020 125630 583060
rect 125560 582970 125630 583020
rect 125350 582920 125630 582970
rect 125420 582330 125650 582380
rect 125420 582280 125490 582330
rect 125420 582240 125430 582280
rect 125470 582240 125490 582280
rect 125420 582190 125490 582240
rect 125520 582280 125650 582300
rect 125520 582240 125540 582280
rect 125630 582240 125650 582280
rect 125520 582220 125650 582240
rect 125680 582280 125750 582380
rect 125680 582240 125700 582280
rect 125740 582240 125750 582280
rect 125680 582190 125750 582240
rect 125420 582140 125750 582190
rect 125810 582330 126040 582380
rect 125810 582280 125880 582330
rect 125810 582240 125820 582280
rect 125860 582240 125880 582280
rect 125810 582190 125880 582240
rect 125910 582280 126040 582300
rect 125910 582240 125930 582280
rect 126020 582240 126040 582280
rect 125910 582220 126040 582240
rect 126070 582280 126140 582380
rect 126070 582240 126090 582280
rect 126130 582240 126140 582280
rect 126070 582190 126140 582240
rect 125810 582140 126140 582190
rect 126200 582330 126430 582380
rect 126200 582280 126270 582330
rect 126200 582240 126210 582280
rect 126250 582240 126270 582280
rect 126200 582190 126270 582240
rect 126300 582280 126430 582300
rect 126300 582240 126320 582280
rect 126410 582240 126430 582280
rect 126300 582220 126430 582240
rect 126460 582280 126530 582380
rect 126460 582240 126480 582280
rect 126520 582240 126530 582280
rect 126460 582190 126530 582240
rect 126200 582140 126530 582190
rect 126590 582330 126820 582380
rect 126590 582280 126660 582330
rect 126590 582240 126600 582280
rect 126640 582240 126660 582280
rect 126590 582190 126660 582240
rect 126690 582280 126820 582300
rect 126690 582240 126710 582280
rect 126800 582240 126820 582280
rect 126690 582220 126820 582240
rect 126850 582280 126920 582380
rect 126850 582240 126870 582280
rect 126910 582240 126920 582280
rect 126850 582190 126920 582240
rect 126590 582140 126920 582190
rect 126980 582330 127210 582380
rect 126980 582280 127050 582330
rect 126980 582240 126990 582280
rect 127030 582240 127050 582280
rect 126980 582190 127050 582240
rect 127080 582280 127210 582300
rect 127080 582240 127100 582280
rect 127190 582240 127210 582280
rect 127080 582220 127210 582240
rect 127240 582280 127310 582380
rect 127240 582240 127260 582280
rect 127300 582240 127310 582280
rect 127240 582190 127310 582240
rect 126980 582140 127310 582190
rect 127370 582330 127600 582380
rect 127370 582280 127440 582330
rect 127370 582240 127380 582280
rect 127420 582240 127440 582280
rect 127370 582190 127440 582240
rect 127470 582280 127600 582300
rect 127470 582240 127490 582280
rect 127580 582240 127600 582280
rect 127470 582220 127600 582240
rect 127630 582280 127700 582380
rect 127630 582240 127650 582280
rect 127690 582240 127700 582280
rect 127630 582190 127700 582240
rect 127370 582140 127700 582190
rect 127760 582330 127990 582380
rect 127760 582280 127830 582330
rect 127760 582240 127770 582280
rect 127810 582240 127830 582280
rect 127760 582190 127830 582240
rect 127860 582280 127990 582300
rect 127860 582240 127880 582280
rect 127970 582240 127990 582280
rect 127860 582220 127990 582240
rect 128020 582280 128090 582380
rect 128020 582240 128040 582280
rect 128080 582240 128090 582280
rect 128020 582190 128090 582240
rect 127760 582140 128090 582190
rect 128150 582330 128380 582380
rect 128150 582280 128220 582330
rect 128150 582240 128160 582280
rect 128200 582240 128220 582280
rect 128150 582190 128220 582240
rect 128250 582280 128380 582300
rect 128250 582240 128270 582280
rect 128360 582240 128380 582280
rect 128250 582220 128380 582240
rect 128410 582280 128480 582380
rect 128410 582240 128430 582280
rect 128470 582240 128480 582280
rect 128410 582190 128480 582240
rect 128150 582140 128480 582190
rect 128540 582330 128770 582380
rect 128540 582280 128610 582330
rect 128540 582240 128550 582280
rect 128590 582240 128610 582280
rect 128540 582190 128610 582240
rect 128640 582280 128770 582300
rect 128640 582240 128660 582280
rect 128750 582240 128770 582280
rect 128640 582220 128770 582240
rect 128800 582280 128870 582380
rect 128800 582240 128820 582280
rect 128860 582240 128870 582280
rect 128800 582190 128870 582240
rect 128540 582140 128870 582190
rect 128930 582330 129160 582380
rect 128930 582280 129000 582330
rect 128930 582240 128940 582280
rect 128980 582240 129000 582280
rect 128930 582190 129000 582240
rect 129030 582280 129160 582300
rect 129030 582240 129050 582280
rect 129140 582240 129160 582280
rect 129030 582220 129160 582240
rect 129190 582280 129260 582380
rect 129190 582240 129210 582280
rect 129250 582240 129260 582280
rect 129190 582190 129260 582240
rect 128930 582140 129260 582190
rect 129320 582330 129550 582380
rect 129320 582280 129390 582330
rect 129320 582240 129330 582280
rect 129370 582240 129390 582280
rect 129320 582190 129390 582240
rect 129420 582280 129550 582300
rect 129420 582240 129440 582280
rect 129530 582240 129550 582280
rect 129420 582220 129550 582240
rect 129580 582280 129650 582380
rect 129580 582240 129600 582280
rect 129640 582240 129650 582280
rect 129580 582190 129650 582240
rect 129320 582140 129650 582190
rect 129710 582330 129940 582380
rect 129710 582280 129780 582330
rect 129710 582240 129720 582280
rect 129760 582240 129780 582280
rect 129710 582190 129780 582240
rect 129810 582280 129940 582300
rect 129810 582240 129830 582280
rect 129920 582240 129940 582280
rect 129810 582220 129940 582240
rect 129970 582280 130040 582380
rect 129970 582240 129990 582280
rect 130030 582240 130040 582280
rect 129970 582190 130040 582240
rect 129710 582140 130040 582190
rect 130100 582330 130330 582380
rect 130100 582280 130170 582330
rect 130100 582240 130110 582280
rect 130150 582240 130170 582280
rect 130100 582190 130170 582240
rect 130200 582280 130330 582300
rect 130200 582240 130220 582280
rect 130310 582240 130330 582280
rect 130200 582220 130330 582240
rect 130360 582280 130430 582380
rect 130360 582240 130380 582280
rect 130420 582240 130430 582280
rect 130360 582190 130430 582240
rect 130100 582140 130430 582190
rect 130490 582330 130720 582380
rect 130490 582280 130560 582330
rect 130490 582240 130500 582280
rect 130540 582240 130560 582280
rect 130490 582190 130560 582240
rect 130590 582280 130720 582300
rect 130590 582240 130610 582280
rect 130700 582240 130720 582280
rect 130590 582220 130720 582240
rect 130750 582280 130820 582380
rect 130750 582240 130770 582280
rect 130810 582240 130820 582280
rect 130750 582190 130820 582240
rect 130490 582140 130820 582190
rect 130880 582330 131110 582380
rect 130880 582280 130950 582330
rect 130880 582240 130890 582280
rect 130930 582240 130950 582280
rect 130880 582190 130950 582240
rect 130980 582280 131110 582300
rect 130980 582240 131000 582280
rect 131090 582240 131110 582280
rect 130980 582220 131110 582240
rect 131140 582280 131210 582380
rect 131140 582240 131160 582280
rect 131200 582240 131210 582280
rect 131140 582190 131210 582240
rect 130880 582140 131210 582190
rect 131270 582330 131500 582380
rect 131270 582280 131340 582330
rect 131270 582240 131280 582280
rect 131320 582240 131340 582280
rect 131270 582190 131340 582240
rect 131370 582280 131500 582300
rect 131370 582240 131390 582280
rect 131480 582240 131500 582280
rect 131370 582220 131500 582240
rect 131530 582280 131600 582380
rect 131530 582240 131550 582280
rect 131590 582240 131600 582280
rect 131530 582190 131600 582240
rect 131270 582140 131600 582190
rect 131660 582330 131890 582380
rect 131660 582280 131730 582330
rect 131660 582240 131670 582280
rect 131710 582240 131730 582280
rect 131660 582190 131730 582240
rect 131760 582280 131890 582300
rect 131760 582240 131780 582280
rect 131870 582240 131890 582280
rect 131760 582220 131890 582240
rect 131920 582280 131990 582380
rect 131920 582240 131940 582280
rect 131980 582240 131990 582280
rect 131920 582190 131990 582240
rect 131660 582140 131990 582190
rect 132050 582330 132280 582380
rect 132050 582280 132120 582330
rect 132050 582240 132060 582280
rect 132100 582240 132120 582280
rect 132050 582190 132120 582240
rect 132150 582280 132280 582300
rect 132150 582240 132170 582280
rect 132260 582240 132280 582280
rect 132150 582220 132280 582240
rect 132310 582280 132380 582380
rect 132310 582240 132330 582280
rect 132370 582240 132380 582280
rect 132310 582190 132380 582240
rect 132050 582140 132380 582190
rect 132440 582330 132670 582380
rect 132440 582280 132510 582330
rect 132440 582240 132450 582280
rect 132490 582240 132510 582280
rect 132440 582190 132510 582240
rect 132540 582280 132670 582300
rect 132540 582240 132560 582280
rect 132650 582240 132670 582280
rect 132540 582220 132670 582240
rect 132700 582280 132770 582380
rect 132700 582240 132720 582280
rect 132760 582240 132770 582280
rect 132700 582190 132770 582240
rect 132440 582140 132770 582190
rect 119340 574390 119410 574410
rect 119340 574340 119350 574390
rect 119390 574340 119410 574390
rect 119340 574320 119410 574340
rect 119440 574390 119510 574410
rect 119440 574340 119460 574390
rect 119500 574340 119510 574390
rect 119440 574320 119510 574340
rect 119700 574190 119770 574210
rect 119700 574030 119710 574190
rect 119750 574030 119770 574190
rect 119700 574010 119770 574030
rect 119800 574190 119870 574210
rect 119800 574030 119820 574190
rect 119860 574030 119870 574190
rect 119800 574010 119870 574030
rect 120080 574190 120150 574210
rect 120080 574030 120090 574190
rect 120130 574030 120150 574190
rect 120080 574010 120150 574030
rect 120180 574190 120250 574210
rect 120180 574030 120200 574190
rect 120240 574030 120250 574190
rect 120180 574010 120250 574030
rect 125390 574090 125570 574140
rect 125390 574040 125460 574090
rect 125390 574000 125400 574040
rect 125440 574000 125460 574040
rect 125390 573950 125460 574000
rect 125490 574040 125570 574060
rect 125490 574000 125510 574040
rect 125550 574000 125570 574040
rect 125490 573980 125570 574000
rect 125600 574040 125670 574140
rect 125600 574000 125620 574040
rect 125660 574000 125670 574040
rect 125600 573950 125670 574000
rect 125390 573900 125670 573950
rect 125460 573310 125690 573360
rect 125460 573260 125530 573310
rect 125460 573120 125470 573260
rect 125510 573120 125530 573260
rect 125460 573070 125530 573120
rect 125560 573260 125690 573280
rect 125560 573120 125580 573260
rect 125670 573120 125690 573260
rect 125560 573100 125690 573120
rect 125720 573260 125790 573360
rect 125720 573120 125740 573260
rect 125780 573120 125790 573260
rect 125720 573070 125790 573120
rect 125460 573020 125790 573070
rect 125850 573310 126080 573360
rect 125850 573260 125920 573310
rect 125850 573120 125860 573260
rect 125900 573120 125920 573260
rect 125850 573070 125920 573120
rect 125950 573260 126080 573280
rect 125950 573120 125970 573260
rect 126060 573120 126080 573260
rect 125950 573100 126080 573120
rect 126110 573260 126180 573360
rect 126110 573120 126130 573260
rect 126170 573120 126180 573260
rect 126110 573070 126180 573120
rect 125850 573020 126180 573070
rect 126240 573310 126470 573360
rect 126240 573260 126310 573310
rect 126240 573120 126250 573260
rect 126290 573120 126310 573260
rect 126240 573070 126310 573120
rect 126340 573260 126470 573280
rect 126340 573120 126360 573260
rect 126450 573120 126470 573260
rect 126340 573100 126470 573120
rect 126500 573260 126570 573360
rect 126500 573120 126520 573260
rect 126560 573120 126570 573260
rect 126500 573070 126570 573120
rect 126240 573020 126570 573070
rect 126630 573310 126860 573360
rect 126630 573260 126700 573310
rect 126630 573120 126640 573260
rect 126680 573120 126700 573260
rect 126630 573070 126700 573120
rect 126730 573260 126860 573280
rect 126730 573120 126750 573260
rect 126840 573120 126860 573260
rect 126730 573100 126860 573120
rect 126890 573260 126960 573360
rect 126890 573120 126910 573260
rect 126950 573120 126960 573260
rect 126890 573070 126960 573120
rect 126630 573020 126960 573070
rect 127020 573310 127250 573360
rect 127020 573260 127090 573310
rect 127020 573120 127030 573260
rect 127070 573120 127090 573260
rect 127020 573070 127090 573120
rect 127120 573260 127250 573280
rect 127120 573120 127140 573260
rect 127230 573120 127250 573260
rect 127120 573100 127250 573120
rect 127280 573260 127350 573360
rect 127280 573120 127300 573260
rect 127340 573120 127350 573260
rect 127280 573070 127350 573120
rect 127020 573020 127350 573070
rect 127410 573310 127640 573360
rect 127410 573260 127480 573310
rect 127410 573120 127420 573260
rect 127460 573120 127480 573260
rect 127410 573070 127480 573120
rect 127510 573260 127640 573280
rect 127510 573120 127530 573260
rect 127620 573120 127640 573260
rect 127510 573100 127640 573120
rect 127670 573260 127740 573360
rect 127670 573120 127690 573260
rect 127730 573120 127740 573260
rect 127670 573070 127740 573120
rect 127410 573020 127740 573070
rect 127800 573310 128030 573360
rect 127800 573260 127870 573310
rect 127800 573120 127810 573260
rect 127850 573120 127870 573260
rect 127800 573070 127870 573120
rect 127900 573260 128030 573280
rect 127900 573120 127920 573260
rect 128010 573120 128030 573260
rect 127900 573100 128030 573120
rect 128060 573260 128130 573360
rect 128060 573120 128080 573260
rect 128120 573120 128130 573260
rect 128060 573070 128130 573120
rect 127800 573020 128130 573070
rect 128190 573310 128420 573360
rect 128190 573260 128260 573310
rect 128190 573120 128200 573260
rect 128240 573120 128260 573260
rect 128190 573070 128260 573120
rect 128290 573260 128420 573280
rect 128290 573120 128310 573260
rect 128400 573120 128420 573260
rect 128290 573100 128420 573120
rect 128450 573260 128520 573360
rect 128450 573120 128470 573260
rect 128510 573120 128520 573260
rect 128450 573070 128520 573120
rect 128190 573020 128520 573070
rect 128580 573310 128810 573360
rect 128580 573260 128650 573310
rect 128580 573120 128590 573260
rect 128630 573120 128650 573260
rect 128580 573070 128650 573120
rect 128680 573260 128810 573280
rect 128680 573120 128700 573260
rect 128790 573120 128810 573260
rect 128680 573100 128810 573120
rect 128840 573260 128910 573360
rect 128840 573120 128860 573260
rect 128900 573120 128910 573260
rect 128840 573070 128910 573120
rect 128580 573020 128910 573070
rect 128970 573310 129200 573360
rect 128970 573260 129040 573310
rect 128970 573120 128980 573260
rect 129020 573120 129040 573260
rect 128970 573070 129040 573120
rect 129070 573260 129200 573280
rect 129070 573120 129090 573260
rect 129180 573120 129200 573260
rect 129070 573100 129200 573120
rect 129230 573260 129300 573360
rect 129230 573120 129250 573260
rect 129290 573120 129300 573260
rect 129230 573070 129300 573120
rect 128970 573020 129300 573070
rect 129360 573310 129590 573360
rect 129360 573260 129430 573310
rect 129360 573120 129370 573260
rect 129410 573120 129430 573260
rect 129360 573070 129430 573120
rect 129460 573260 129590 573280
rect 129460 573120 129480 573260
rect 129570 573120 129590 573260
rect 129460 573100 129590 573120
rect 129620 573260 129690 573360
rect 129620 573120 129640 573260
rect 129680 573120 129690 573260
rect 129620 573070 129690 573120
rect 129360 573020 129690 573070
rect 129750 573310 129980 573360
rect 129750 573260 129820 573310
rect 129750 573120 129760 573260
rect 129800 573120 129820 573260
rect 129750 573070 129820 573120
rect 129850 573260 129980 573280
rect 129850 573120 129870 573260
rect 129960 573120 129980 573260
rect 129850 573100 129980 573120
rect 130010 573260 130080 573360
rect 130010 573120 130030 573260
rect 130070 573120 130080 573260
rect 130010 573070 130080 573120
rect 129750 573020 130080 573070
rect 130140 573310 130370 573360
rect 130140 573260 130210 573310
rect 130140 573120 130150 573260
rect 130190 573120 130210 573260
rect 130140 573070 130210 573120
rect 130240 573260 130370 573280
rect 130240 573120 130260 573260
rect 130350 573120 130370 573260
rect 130240 573100 130370 573120
rect 130400 573260 130470 573360
rect 130400 573120 130420 573260
rect 130460 573120 130470 573260
rect 130400 573070 130470 573120
rect 130140 573020 130470 573070
rect 130530 573310 130760 573360
rect 130530 573260 130600 573310
rect 130530 573120 130540 573260
rect 130580 573120 130600 573260
rect 130530 573070 130600 573120
rect 130630 573260 130760 573280
rect 130630 573120 130650 573260
rect 130740 573120 130760 573260
rect 130630 573100 130760 573120
rect 130790 573260 130860 573360
rect 130790 573120 130810 573260
rect 130850 573120 130860 573260
rect 130790 573070 130860 573120
rect 130530 573020 130860 573070
rect 130920 573310 131150 573360
rect 130920 573260 130990 573310
rect 130920 573120 130930 573260
rect 130970 573120 130990 573260
rect 130920 573070 130990 573120
rect 131020 573260 131150 573280
rect 131020 573120 131040 573260
rect 131130 573120 131150 573260
rect 131020 573100 131150 573120
rect 131180 573260 131250 573360
rect 131180 573120 131200 573260
rect 131240 573120 131250 573260
rect 131180 573070 131250 573120
rect 130920 573020 131250 573070
rect 131310 573310 131540 573360
rect 131310 573260 131380 573310
rect 131310 573120 131320 573260
rect 131360 573120 131380 573260
rect 131310 573070 131380 573120
rect 131410 573260 131540 573280
rect 131410 573120 131430 573260
rect 131520 573120 131540 573260
rect 131410 573100 131540 573120
rect 131570 573260 131640 573360
rect 131570 573120 131590 573260
rect 131630 573120 131640 573260
rect 131570 573070 131640 573120
rect 131310 573020 131640 573070
rect 131700 573310 131930 573360
rect 131700 573260 131770 573310
rect 131700 573120 131710 573260
rect 131750 573120 131770 573260
rect 131700 573070 131770 573120
rect 131800 573260 131930 573280
rect 131800 573120 131820 573260
rect 131910 573120 131930 573260
rect 131800 573100 131930 573120
rect 131960 573260 132030 573360
rect 131960 573120 131980 573260
rect 132020 573120 132030 573260
rect 131960 573070 132030 573120
rect 131700 573020 132030 573070
rect 132090 573310 132320 573360
rect 132090 573260 132160 573310
rect 132090 573120 132100 573260
rect 132140 573120 132160 573260
rect 132090 573070 132160 573120
rect 132190 573260 132320 573280
rect 132190 573120 132210 573260
rect 132300 573120 132320 573260
rect 132190 573100 132320 573120
rect 132350 573260 132420 573360
rect 132350 573120 132370 573260
rect 132410 573120 132420 573260
rect 132350 573070 132420 573120
rect 132090 573020 132420 573070
rect 132480 573310 132710 573360
rect 132480 573260 132550 573310
rect 132480 573120 132490 573260
rect 132530 573120 132550 573260
rect 132480 573070 132550 573120
rect 132580 573260 132710 573280
rect 132580 573120 132600 573260
rect 132690 573120 132710 573260
rect 132580 573100 132710 573120
rect 132740 573260 132810 573360
rect 132740 573120 132760 573260
rect 132800 573120 132810 573260
rect 132740 573070 132810 573120
rect 132480 573020 132810 573070
rect 119290 566720 119360 566740
rect 119290 566670 119300 566720
rect 119340 566670 119360 566720
rect 119290 566650 119360 566670
rect 119390 566720 119460 566740
rect 119390 566670 119410 566720
rect 119450 566670 119460 566720
rect 119390 566650 119460 566670
rect 119650 566520 119720 566540
rect 119650 566360 119660 566520
rect 119700 566360 119720 566520
rect 119650 566340 119720 566360
rect 119750 566520 119820 566540
rect 119750 566360 119770 566520
rect 119810 566360 119820 566520
rect 119750 566340 119820 566360
rect 120030 566520 120100 566540
rect 120030 566360 120040 566520
rect 120080 566360 120100 566520
rect 120030 566340 120100 566360
rect 120130 566520 120200 566540
rect 120130 566360 120150 566520
rect 120190 566360 120200 566520
rect 120130 566340 120200 566360
rect 125340 566420 125520 566470
rect 125340 566370 125410 566420
rect 125340 566330 125350 566370
rect 125390 566330 125410 566370
rect 125340 566280 125410 566330
rect 125440 566370 125520 566390
rect 125440 566330 125460 566370
rect 125500 566330 125520 566370
rect 125440 566310 125520 566330
rect 125550 566370 125620 566470
rect 125550 566330 125570 566370
rect 125610 566330 125620 566370
rect 125550 566280 125620 566330
rect 125340 566230 125620 566280
rect 125410 565640 125640 565690
rect 125410 565590 125480 565640
rect 125410 565350 125420 565590
rect 125460 565350 125480 565590
rect 125410 565300 125480 565350
rect 125510 565590 125640 565610
rect 125510 565350 125530 565590
rect 125620 565350 125640 565590
rect 125510 565330 125640 565350
rect 125670 565590 125740 565690
rect 125670 565350 125690 565590
rect 125730 565350 125740 565590
rect 125670 565300 125740 565350
rect 125410 565250 125740 565300
rect 125800 565640 126030 565690
rect 125800 565590 125870 565640
rect 125800 565350 125810 565590
rect 125850 565350 125870 565590
rect 125800 565300 125870 565350
rect 125900 565590 126030 565610
rect 125900 565350 125920 565590
rect 126010 565350 126030 565590
rect 125900 565330 126030 565350
rect 126060 565590 126130 565690
rect 126060 565350 126080 565590
rect 126120 565350 126130 565590
rect 126060 565300 126130 565350
rect 125800 565250 126130 565300
rect 126190 565640 126420 565690
rect 126190 565590 126260 565640
rect 126190 565350 126200 565590
rect 126240 565350 126260 565590
rect 126190 565300 126260 565350
rect 126290 565590 126420 565610
rect 126290 565350 126310 565590
rect 126400 565350 126420 565590
rect 126290 565330 126420 565350
rect 126450 565590 126520 565690
rect 126450 565350 126470 565590
rect 126510 565350 126520 565590
rect 126450 565300 126520 565350
rect 126190 565250 126520 565300
rect 126580 565640 126810 565690
rect 126580 565590 126650 565640
rect 126580 565350 126590 565590
rect 126630 565350 126650 565590
rect 126580 565300 126650 565350
rect 126680 565590 126810 565610
rect 126680 565350 126700 565590
rect 126790 565350 126810 565590
rect 126680 565330 126810 565350
rect 126840 565590 126910 565690
rect 126840 565350 126860 565590
rect 126900 565350 126910 565590
rect 126840 565300 126910 565350
rect 126580 565250 126910 565300
rect 126970 565640 127200 565690
rect 126970 565590 127040 565640
rect 126970 565350 126980 565590
rect 127020 565350 127040 565590
rect 126970 565300 127040 565350
rect 127070 565590 127200 565610
rect 127070 565350 127090 565590
rect 127180 565350 127200 565590
rect 127070 565330 127200 565350
rect 127230 565590 127300 565690
rect 127230 565350 127250 565590
rect 127290 565350 127300 565590
rect 127230 565300 127300 565350
rect 126970 565250 127300 565300
rect 127360 565640 127590 565690
rect 127360 565590 127430 565640
rect 127360 565350 127370 565590
rect 127410 565350 127430 565590
rect 127360 565300 127430 565350
rect 127460 565590 127590 565610
rect 127460 565350 127480 565590
rect 127570 565350 127590 565590
rect 127460 565330 127590 565350
rect 127620 565590 127690 565690
rect 127620 565350 127640 565590
rect 127680 565350 127690 565590
rect 127620 565300 127690 565350
rect 127360 565250 127690 565300
rect 127750 565640 127980 565690
rect 127750 565590 127820 565640
rect 127750 565350 127760 565590
rect 127800 565350 127820 565590
rect 127750 565300 127820 565350
rect 127850 565590 127980 565610
rect 127850 565350 127870 565590
rect 127960 565350 127980 565590
rect 127850 565330 127980 565350
rect 128010 565590 128080 565690
rect 128010 565350 128030 565590
rect 128070 565350 128080 565590
rect 128010 565300 128080 565350
rect 127750 565250 128080 565300
rect 128140 565640 128370 565690
rect 128140 565590 128210 565640
rect 128140 565350 128150 565590
rect 128190 565350 128210 565590
rect 128140 565300 128210 565350
rect 128240 565590 128370 565610
rect 128240 565350 128260 565590
rect 128350 565350 128370 565590
rect 128240 565330 128370 565350
rect 128400 565590 128470 565690
rect 128400 565350 128420 565590
rect 128460 565350 128470 565590
rect 128400 565300 128470 565350
rect 128140 565250 128470 565300
rect 128530 565640 128760 565690
rect 128530 565590 128600 565640
rect 128530 565350 128540 565590
rect 128580 565350 128600 565590
rect 128530 565300 128600 565350
rect 128630 565590 128760 565610
rect 128630 565350 128650 565590
rect 128740 565350 128760 565590
rect 128630 565330 128760 565350
rect 128790 565590 128860 565690
rect 128790 565350 128810 565590
rect 128850 565350 128860 565590
rect 128790 565300 128860 565350
rect 128530 565250 128860 565300
rect 128920 565640 129150 565690
rect 128920 565590 128990 565640
rect 128920 565350 128930 565590
rect 128970 565350 128990 565590
rect 128920 565300 128990 565350
rect 129020 565590 129150 565610
rect 129020 565350 129040 565590
rect 129130 565350 129150 565590
rect 129020 565330 129150 565350
rect 129180 565590 129250 565690
rect 129180 565350 129200 565590
rect 129240 565350 129250 565590
rect 129180 565300 129250 565350
rect 128920 565250 129250 565300
rect 129310 565640 129540 565690
rect 129310 565590 129380 565640
rect 129310 565350 129320 565590
rect 129360 565350 129380 565590
rect 129310 565300 129380 565350
rect 129410 565590 129540 565610
rect 129410 565350 129430 565590
rect 129520 565350 129540 565590
rect 129410 565330 129540 565350
rect 129570 565590 129640 565690
rect 129570 565350 129590 565590
rect 129630 565350 129640 565590
rect 129570 565300 129640 565350
rect 129310 565250 129640 565300
rect 129700 565640 129930 565690
rect 129700 565590 129770 565640
rect 129700 565350 129710 565590
rect 129750 565350 129770 565590
rect 129700 565300 129770 565350
rect 129800 565590 129930 565610
rect 129800 565350 129820 565590
rect 129910 565350 129930 565590
rect 129800 565330 129930 565350
rect 129960 565590 130030 565690
rect 129960 565350 129980 565590
rect 130020 565350 130030 565590
rect 129960 565300 130030 565350
rect 129700 565250 130030 565300
rect 130090 565640 130320 565690
rect 130090 565590 130160 565640
rect 130090 565350 130100 565590
rect 130140 565350 130160 565590
rect 130090 565300 130160 565350
rect 130190 565590 130320 565610
rect 130190 565350 130210 565590
rect 130300 565350 130320 565590
rect 130190 565330 130320 565350
rect 130350 565590 130420 565690
rect 130350 565350 130370 565590
rect 130410 565350 130420 565590
rect 130350 565300 130420 565350
rect 130090 565250 130420 565300
rect 130480 565640 130710 565690
rect 130480 565590 130550 565640
rect 130480 565350 130490 565590
rect 130530 565350 130550 565590
rect 130480 565300 130550 565350
rect 130580 565590 130710 565610
rect 130580 565350 130600 565590
rect 130690 565350 130710 565590
rect 130580 565330 130710 565350
rect 130740 565590 130810 565690
rect 130740 565350 130760 565590
rect 130800 565350 130810 565590
rect 130740 565300 130810 565350
rect 130480 565250 130810 565300
rect 130870 565640 131100 565690
rect 130870 565590 130940 565640
rect 130870 565350 130880 565590
rect 130920 565350 130940 565590
rect 130870 565300 130940 565350
rect 130970 565590 131100 565610
rect 130970 565350 130990 565590
rect 131080 565350 131100 565590
rect 130970 565330 131100 565350
rect 131130 565590 131200 565690
rect 131130 565350 131150 565590
rect 131190 565350 131200 565590
rect 131130 565300 131200 565350
rect 130870 565250 131200 565300
rect 131260 565640 131490 565690
rect 131260 565590 131330 565640
rect 131260 565350 131270 565590
rect 131310 565350 131330 565590
rect 131260 565300 131330 565350
rect 131360 565590 131490 565610
rect 131360 565350 131380 565590
rect 131470 565350 131490 565590
rect 131360 565330 131490 565350
rect 131520 565590 131590 565690
rect 131520 565350 131540 565590
rect 131580 565350 131590 565590
rect 131520 565300 131590 565350
rect 131260 565250 131590 565300
rect 131650 565640 131880 565690
rect 131650 565590 131720 565640
rect 131650 565350 131660 565590
rect 131700 565350 131720 565590
rect 131650 565300 131720 565350
rect 131750 565590 131880 565610
rect 131750 565350 131770 565590
rect 131860 565350 131880 565590
rect 131750 565330 131880 565350
rect 131910 565590 131980 565690
rect 131910 565350 131930 565590
rect 131970 565350 131980 565590
rect 131910 565300 131980 565350
rect 131650 565250 131980 565300
rect 132040 565640 132270 565690
rect 132040 565590 132110 565640
rect 132040 565350 132050 565590
rect 132090 565350 132110 565590
rect 132040 565300 132110 565350
rect 132140 565590 132270 565610
rect 132140 565350 132160 565590
rect 132250 565350 132270 565590
rect 132140 565330 132270 565350
rect 132300 565590 132370 565690
rect 132300 565350 132320 565590
rect 132360 565350 132370 565590
rect 132300 565300 132370 565350
rect 132040 565250 132370 565300
rect 132430 565640 132660 565690
rect 132430 565590 132500 565640
rect 132430 565350 132440 565590
rect 132480 565350 132500 565590
rect 132430 565300 132500 565350
rect 132530 565590 132660 565610
rect 132530 565350 132550 565590
rect 132640 565350 132660 565590
rect 132530 565330 132660 565350
rect 132690 565590 132760 565690
rect 132690 565350 132710 565590
rect 132750 565350 132760 565590
rect 132690 565300 132760 565350
rect 132430 565250 132760 565300
rect 119290 560180 119360 560200
rect 119290 560130 119300 560180
rect 119340 560130 119360 560180
rect 119290 560110 119360 560130
rect 119390 560180 119460 560200
rect 119390 560130 119410 560180
rect 119450 560130 119460 560180
rect 119390 560110 119460 560130
rect 119650 559980 119720 560000
rect 119650 559820 119660 559980
rect 119700 559820 119720 559980
rect 119650 559800 119720 559820
rect 119750 559980 119820 560000
rect 119750 559820 119770 559980
rect 119810 559820 119820 559980
rect 119750 559800 119820 559820
rect 120030 559980 120100 560000
rect 120030 559820 120040 559980
rect 120080 559820 120100 559980
rect 120030 559800 120100 559820
rect 120130 559980 120200 560000
rect 120130 559820 120150 559980
rect 120190 559820 120200 559980
rect 120130 559800 120200 559820
rect 125340 559880 125520 559930
rect 125340 559830 125410 559880
rect 125340 559790 125350 559830
rect 125390 559790 125410 559830
rect 125340 559740 125410 559790
rect 125440 559830 125520 559850
rect 125440 559790 125460 559830
rect 125500 559790 125520 559830
rect 125440 559770 125520 559790
rect 125550 559830 125620 559930
rect 125550 559790 125570 559830
rect 125610 559790 125620 559830
rect 125550 559740 125620 559790
rect 125340 559690 125620 559740
rect 125410 559100 125640 559150
rect 125410 559050 125480 559100
rect 125410 558710 125420 559050
rect 125460 558710 125480 559050
rect 125410 558660 125480 558710
rect 125510 559050 125640 559070
rect 125510 558710 125530 559050
rect 125620 558710 125640 559050
rect 125510 558690 125640 558710
rect 125670 559050 125740 559150
rect 125670 558710 125690 559050
rect 125730 558710 125740 559050
rect 125670 558660 125740 558710
rect 125410 558610 125740 558660
rect 125800 559100 126030 559150
rect 125800 559050 125870 559100
rect 125800 558710 125810 559050
rect 125850 558710 125870 559050
rect 125800 558660 125870 558710
rect 125900 559050 126030 559070
rect 125900 558710 125920 559050
rect 126010 558710 126030 559050
rect 125900 558690 126030 558710
rect 126060 559050 126130 559150
rect 126060 558710 126080 559050
rect 126120 558710 126130 559050
rect 126060 558660 126130 558710
rect 125800 558610 126130 558660
rect 126190 559100 126420 559150
rect 126190 559050 126260 559100
rect 126190 558710 126200 559050
rect 126240 558710 126260 559050
rect 126190 558660 126260 558710
rect 126290 559050 126420 559070
rect 126290 558710 126310 559050
rect 126400 558710 126420 559050
rect 126290 558690 126420 558710
rect 126450 559050 126520 559150
rect 126450 558710 126470 559050
rect 126510 558710 126520 559050
rect 126450 558660 126520 558710
rect 126190 558610 126520 558660
rect 126580 559100 126810 559150
rect 126580 559050 126650 559100
rect 126580 558710 126590 559050
rect 126630 558710 126650 559050
rect 126580 558660 126650 558710
rect 126680 559050 126810 559070
rect 126680 558710 126700 559050
rect 126790 558710 126810 559050
rect 126680 558690 126810 558710
rect 126840 559050 126910 559150
rect 126840 558710 126860 559050
rect 126900 558710 126910 559050
rect 126840 558660 126910 558710
rect 126580 558610 126910 558660
rect 126970 559100 127200 559150
rect 126970 559050 127040 559100
rect 126970 558710 126980 559050
rect 127020 558710 127040 559050
rect 126970 558660 127040 558710
rect 127070 559050 127200 559070
rect 127070 558710 127090 559050
rect 127180 558710 127200 559050
rect 127070 558690 127200 558710
rect 127230 559050 127300 559150
rect 127230 558710 127250 559050
rect 127290 558710 127300 559050
rect 127230 558660 127300 558710
rect 126970 558610 127300 558660
rect 127360 559100 127590 559150
rect 127360 559050 127430 559100
rect 127360 558710 127370 559050
rect 127410 558710 127430 559050
rect 127360 558660 127430 558710
rect 127460 559050 127590 559070
rect 127460 558710 127480 559050
rect 127570 558710 127590 559050
rect 127460 558690 127590 558710
rect 127620 559050 127690 559150
rect 127620 558710 127640 559050
rect 127680 558710 127690 559050
rect 127620 558660 127690 558710
rect 127360 558610 127690 558660
rect 127750 559100 127980 559150
rect 127750 559050 127820 559100
rect 127750 558710 127760 559050
rect 127800 558710 127820 559050
rect 127750 558660 127820 558710
rect 127850 559050 127980 559070
rect 127850 558710 127870 559050
rect 127960 558710 127980 559050
rect 127850 558690 127980 558710
rect 128010 559050 128080 559150
rect 128010 558710 128030 559050
rect 128070 558710 128080 559050
rect 128010 558660 128080 558710
rect 127750 558610 128080 558660
rect 128140 559100 128370 559150
rect 128140 559050 128210 559100
rect 128140 558710 128150 559050
rect 128190 558710 128210 559050
rect 128140 558660 128210 558710
rect 128240 559050 128370 559070
rect 128240 558710 128260 559050
rect 128350 558710 128370 559050
rect 128240 558690 128370 558710
rect 128400 559050 128470 559150
rect 128400 558710 128420 559050
rect 128460 558710 128470 559050
rect 128400 558660 128470 558710
rect 128140 558610 128470 558660
rect 128530 559100 128760 559150
rect 128530 559050 128600 559100
rect 128530 558710 128540 559050
rect 128580 558710 128600 559050
rect 128530 558660 128600 558710
rect 128630 559050 128760 559070
rect 128630 558710 128650 559050
rect 128740 558710 128760 559050
rect 128630 558690 128760 558710
rect 128790 559050 128860 559150
rect 128790 558710 128810 559050
rect 128850 558710 128860 559050
rect 128790 558660 128860 558710
rect 128530 558610 128860 558660
rect 128920 559100 129150 559150
rect 128920 559050 128990 559100
rect 128920 558710 128930 559050
rect 128970 558710 128990 559050
rect 128920 558660 128990 558710
rect 129020 559050 129150 559070
rect 129020 558710 129040 559050
rect 129130 558710 129150 559050
rect 129020 558690 129150 558710
rect 129180 559050 129250 559150
rect 129180 558710 129200 559050
rect 129240 558710 129250 559050
rect 129180 558660 129250 558710
rect 128920 558610 129250 558660
rect 129310 559100 129540 559150
rect 129310 559050 129380 559100
rect 129310 558710 129320 559050
rect 129360 558710 129380 559050
rect 129310 558660 129380 558710
rect 129410 559050 129540 559070
rect 129410 558710 129430 559050
rect 129520 558710 129540 559050
rect 129410 558690 129540 558710
rect 129570 559050 129640 559150
rect 129570 558710 129590 559050
rect 129630 558710 129640 559050
rect 129570 558660 129640 558710
rect 129310 558610 129640 558660
rect 129700 559100 129930 559150
rect 129700 559050 129770 559100
rect 129700 558710 129710 559050
rect 129750 558710 129770 559050
rect 129700 558660 129770 558710
rect 129800 559050 129930 559070
rect 129800 558710 129820 559050
rect 129910 558710 129930 559050
rect 129800 558690 129930 558710
rect 129960 559050 130030 559150
rect 129960 558710 129980 559050
rect 130020 558710 130030 559050
rect 129960 558660 130030 558710
rect 129700 558610 130030 558660
rect 130090 559100 130320 559150
rect 130090 559050 130160 559100
rect 130090 558710 130100 559050
rect 130140 558710 130160 559050
rect 130090 558660 130160 558710
rect 130190 559050 130320 559070
rect 130190 558710 130210 559050
rect 130300 558710 130320 559050
rect 130190 558690 130320 558710
rect 130350 559050 130420 559150
rect 130350 558710 130370 559050
rect 130410 558710 130420 559050
rect 130350 558660 130420 558710
rect 130090 558610 130420 558660
rect 130480 559100 130710 559150
rect 130480 559050 130550 559100
rect 130480 558710 130490 559050
rect 130530 558710 130550 559050
rect 130480 558660 130550 558710
rect 130580 559050 130710 559070
rect 130580 558710 130600 559050
rect 130690 558710 130710 559050
rect 130580 558690 130710 558710
rect 130740 559050 130810 559150
rect 130740 558710 130760 559050
rect 130800 558710 130810 559050
rect 130740 558660 130810 558710
rect 130480 558610 130810 558660
rect 130870 559100 131100 559150
rect 130870 559050 130940 559100
rect 130870 558710 130880 559050
rect 130920 558710 130940 559050
rect 130870 558660 130940 558710
rect 130970 559050 131100 559070
rect 130970 558710 130990 559050
rect 131080 558710 131100 559050
rect 130970 558690 131100 558710
rect 131130 559050 131200 559150
rect 131130 558710 131150 559050
rect 131190 558710 131200 559050
rect 131130 558660 131200 558710
rect 130870 558610 131200 558660
rect 131260 559100 131490 559150
rect 131260 559050 131330 559100
rect 131260 558710 131270 559050
rect 131310 558710 131330 559050
rect 131260 558660 131330 558710
rect 131360 559050 131490 559070
rect 131360 558710 131380 559050
rect 131470 558710 131490 559050
rect 131360 558690 131490 558710
rect 131520 559050 131590 559150
rect 131520 558710 131540 559050
rect 131580 558710 131590 559050
rect 131520 558660 131590 558710
rect 131260 558610 131590 558660
rect 131650 559100 131880 559150
rect 131650 559050 131720 559100
rect 131650 558710 131660 559050
rect 131700 558710 131720 559050
rect 131650 558660 131720 558710
rect 131750 559050 131880 559070
rect 131750 558710 131770 559050
rect 131860 558710 131880 559050
rect 131750 558690 131880 558710
rect 131910 559050 131980 559150
rect 131910 558710 131930 559050
rect 131970 558710 131980 559050
rect 131910 558660 131980 558710
rect 131650 558610 131980 558660
rect 132040 559100 132270 559150
rect 132040 559050 132110 559100
rect 132040 558710 132050 559050
rect 132090 558710 132110 559050
rect 132040 558660 132110 558710
rect 132140 559050 132270 559070
rect 132140 558710 132160 559050
rect 132250 558710 132270 559050
rect 132140 558690 132270 558710
rect 132300 559050 132370 559150
rect 132300 558710 132320 559050
rect 132360 558710 132370 559050
rect 132300 558660 132370 558710
rect 132040 558610 132370 558660
rect 132430 559100 132660 559150
rect 132430 559050 132500 559100
rect 132430 558710 132440 559050
rect 132480 558710 132500 559050
rect 132430 558660 132500 558710
rect 132530 559050 132660 559070
rect 132530 558710 132550 559050
rect 132640 558710 132660 559050
rect 132530 558690 132660 558710
rect 132690 559050 132760 559150
rect 132690 558710 132710 559050
rect 132750 558710 132760 559050
rect 132690 558660 132760 558710
rect 132430 558610 132760 558660
rect 124990 554020 125170 554070
rect 124990 553970 125060 554020
rect 124990 553930 125000 553970
rect 125040 553930 125060 553970
rect 124990 553880 125060 553930
rect 125090 553970 125170 553990
rect 125090 553930 125110 553970
rect 125150 553930 125170 553970
rect 125090 553910 125170 553930
rect 125200 553970 125270 554070
rect 125200 553930 125220 553970
rect 125260 553930 125270 553970
rect 125200 553880 125270 553930
rect 124990 553830 125270 553880
rect 119360 553350 119430 553370
rect 119360 553300 119370 553350
rect 119410 553300 119430 553350
rect 119360 553280 119430 553300
rect 119460 553350 119530 553370
rect 119460 553300 119480 553350
rect 119520 553300 119530 553350
rect 119460 553280 119530 553300
rect 119720 553150 119790 553170
rect 119720 552990 119730 553150
rect 119770 552990 119790 553150
rect 119720 552970 119790 552990
rect 119820 553150 119890 553170
rect 119820 552990 119840 553150
rect 119880 552990 119890 553150
rect 119820 552970 119890 552990
rect 120100 553150 120170 553170
rect 120100 552990 120110 553150
rect 120150 552990 120170 553150
rect 120100 552970 120170 552990
rect 120200 553150 120270 553170
rect 120200 552990 120220 553150
rect 120260 552990 120270 553150
rect 120200 552970 120270 552990
rect 125480 552270 125760 552320
rect 125480 552220 125550 552270
rect 125480 552180 125490 552220
rect 125530 552180 125550 552220
rect 125480 552130 125550 552180
rect 125580 552220 125760 552240
rect 125580 552180 125600 552220
rect 125740 552180 125760 552220
rect 125580 552160 125760 552180
rect 125790 552220 125860 552320
rect 125790 552180 125810 552220
rect 125850 552180 125860 552220
rect 125790 552130 125860 552180
rect 125480 552080 125860 552130
rect 125920 552270 126200 552320
rect 125920 552220 125990 552270
rect 125920 552180 125930 552220
rect 125970 552180 125990 552220
rect 125920 552130 125990 552180
rect 126020 552220 126200 552240
rect 126020 552180 126040 552220
rect 126180 552180 126200 552220
rect 126020 552160 126200 552180
rect 126230 552220 126300 552320
rect 126230 552180 126250 552220
rect 126290 552180 126300 552220
rect 126230 552130 126300 552180
rect 125920 552080 126300 552130
rect 126360 552270 126640 552320
rect 126360 552220 126430 552270
rect 126360 552180 126370 552220
rect 126410 552180 126430 552220
rect 126360 552130 126430 552180
rect 126460 552220 126640 552240
rect 126460 552180 126480 552220
rect 126620 552180 126640 552220
rect 126460 552160 126640 552180
rect 126670 552220 126740 552320
rect 126670 552180 126690 552220
rect 126730 552180 126740 552220
rect 126670 552130 126740 552180
rect 126360 552080 126740 552130
rect 126800 552270 127080 552320
rect 126800 552220 126870 552270
rect 126800 552180 126810 552220
rect 126850 552180 126870 552220
rect 126800 552130 126870 552180
rect 126900 552220 127080 552240
rect 126900 552180 126920 552220
rect 127060 552180 127080 552220
rect 126900 552160 127080 552180
rect 127110 552220 127180 552320
rect 127110 552180 127130 552220
rect 127170 552180 127180 552220
rect 127110 552130 127180 552180
rect 126800 552080 127180 552130
rect 127240 552270 127520 552320
rect 127240 552220 127310 552270
rect 127240 552180 127250 552220
rect 127290 552180 127310 552220
rect 127240 552130 127310 552180
rect 127340 552220 127520 552240
rect 127340 552180 127360 552220
rect 127500 552180 127520 552220
rect 127340 552160 127520 552180
rect 127550 552220 127620 552320
rect 127550 552180 127570 552220
rect 127610 552180 127620 552220
rect 127550 552130 127620 552180
rect 127240 552080 127620 552130
rect 127680 552270 127960 552320
rect 127680 552220 127750 552270
rect 127680 552180 127690 552220
rect 127730 552180 127750 552220
rect 127680 552130 127750 552180
rect 127780 552220 127960 552240
rect 127780 552180 127800 552220
rect 127940 552180 127960 552220
rect 127780 552160 127960 552180
rect 127990 552220 128060 552320
rect 127990 552180 128010 552220
rect 128050 552180 128060 552220
rect 127990 552130 128060 552180
rect 127680 552080 128060 552130
rect 128120 552270 128400 552320
rect 128120 552220 128190 552270
rect 128120 552180 128130 552220
rect 128170 552180 128190 552220
rect 128120 552130 128190 552180
rect 128220 552220 128400 552240
rect 128220 552180 128240 552220
rect 128380 552180 128400 552220
rect 128220 552160 128400 552180
rect 128430 552220 128500 552320
rect 128430 552180 128450 552220
rect 128490 552180 128500 552220
rect 128430 552130 128500 552180
rect 128120 552080 128500 552130
rect 128560 552270 128840 552320
rect 128560 552220 128630 552270
rect 128560 552180 128570 552220
rect 128610 552180 128630 552220
rect 128560 552130 128630 552180
rect 128660 552220 128840 552240
rect 128660 552180 128680 552220
rect 128820 552180 128840 552220
rect 128660 552160 128840 552180
rect 128870 552220 128940 552320
rect 128870 552180 128890 552220
rect 128930 552180 128940 552220
rect 128870 552130 128940 552180
rect 128560 552080 128940 552130
rect 129000 552270 129280 552320
rect 129000 552220 129070 552270
rect 129000 552180 129010 552220
rect 129050 552180 129070 552220
rect 129000 552130 129070 552180
rect 129100 552220 129280 552240
rect 129100 552180 129120 552220
rect 129260 552180 129280 552220
rect 129100 552160 129280 552180
rect 129310 552220 129380 552320
rect 129310 552180 129330 552220
rect 129370 552180 129380 552220
rect 129310 552130 129380 552180
rect 129000 552080 129380 552130
rect 129440 552270 129720 552320
rect 129440 552220 129510 552270
rect 129440 552180 129450 552220
rect 129490 552180 129510 552220
rect 129440 552130 129510 552180
rect 129540 552220 129720 552240
rect 129540 552180 129560 552220
rect 129700 552180 129720 552220
rect 129540 552160 129720 552180
rect 129750 552220 129820 552320
rect 129750 552180 129770 552220
rect 129810 552180 129820 552220
rect 129750 552130 129820 552180
rect 129440 552080 129820 552130
rect 129880 552270 130160 552320
rect 129880 552220 129950 552270
rect 129880 552180 129890 552220
rect 129930 552180 129950 552220
rect 129880 552130 129950 552180
rect 129980 552220 130160 552240
rect 129980 552180 130000 552220
rect 130140 552180 130160 552220
rect 129980 552160 130160 552180
rect 130190 552220 130260 552320
rect 130190 552180 130210 552220
rect 130250 552180 130260 552220
rect 130190 552130 130260 552180
rect 129880 552080 130260 552130
rect 130320 552270 130600 552320
rect 130320 552220 130390 552270
rect 130320 552180 130330 552220
rect 130370 552180 130390 552220
rect 130320 552130 130390 552180
rect 130420 552220 130600 552240
rect 130420 552180 130440 552220
rect 130580 552180 130600 552220
rect 130420 552160 130600 552180
rect 130630 552220 130700 552320
rect 130630 552180 130650 552220
rect 130690 552180 130700 552220
rect 130630 552130 130700 552180
rect 130320 552080 130700 552130
rect 130760 552270 131040 552320
rect 130760 552220 130830 552270
rect 130760 552180 130770 552220
rect 130810 552180 130830 552220
rect 130760 552130 130830 552180
rect 130860 552220 131040 552240
rect 130860 552180 130880 552220
rect 131020 552180 131040 552220
rect 130860 552160 131040 552180
rect 131070 552220 131140 552320
rect 131070 552180 131090 552220
rect 131130 552180 131140 552220
rect 131070 552130 131140 552180
rect 130760 552080 131140 552130
rect 131200 552270 131480 552320
rect 131200 552220 131270 552270
rect 131200 552180 131210 552220
rect 131250 552180 131270 552220
rect 131200 552130 131270 552180
rect 131300 552220 131480 552240
rect 131300 552180 131320 552220
rect 131460 552180 131480 552220
rect 131300 552160 131480 552180
rect 131510 552220 131580 552320
rect 131510 552180 131530 552220
rect 131570 552180 131580 552220
rect 131510 552130 131580 552180
rect 131200 552080 131580 552130
rect 131640 552270 131920 552320
rect 131640 552220 131710 552270
rect 131640 552180 131650 552220
rect 131690 552180 131710 552220
rect 131640 552130 131710 552180
rect 131740 552220 131920 552240
rect 131740 552180 131760 552220
rect 131900 552180 131920 552220
rect 131740 552160 131920 552180
rect 131950 552220 132020 552320
rect 131950 552180 131970 552220
rect 132010 552180 132020 552220
rect 131950 552130 132020 552180
rect 131640 552080 132020 552130
rect 132080 552270 132360 552320
rect 132080 552220 132150 552270
rect 132080 552180 132090 552220
rect 132130 552180 132150 552220
rect 132080 552130 132150 552180
rect 132180 552220 132360 552240
rect 132180 552180 132200 552220
rect 132340 552180 132360 552220
rect 132180 552160 132360 552180
rect 132390 552220 132460 552320
rect 132390 552180 132410 552220
rect 132450 552180 132460 552220
rect 132390 552130 132460 552180
rect 132080 552080 132460 552130
rect 132520 552270 132800 552320
rect 132520 552220 132590 552270
rect 132520 552180 132530 552220
rect 132570 552180 132590 552220
rect 132520 552130 132590 552180
rect 132620 552220 132800 552240
rect 132620 552180 132640 552220
rect 132780 552180 132800 552220
rect 132620 552160 132800 552180
rect 132830 552220 132900 552320
rect 132830 552180 132850 552220
rect 132890 552180 132900 552220
rect 132830 552130 132900 552180
rect 132520 552080 132900 552130
rect 132960 552270 133240 552320
rect 132960 552220 133030 552270
rect 132960 552180 132970 552220
rect 133010 552180 133030 552220
rect 132960 552130 133030 552180
rect 133060 552220 133240 552240
rect 133060 552180 133080 552220
rect 133220 552180 133240 552220
rect 133060 552160 133240 552180
rect 133270 552220 133340 552320
rect 133270 552180 133290 552220
rect 133330 552180 133340 552220
rect 133270 552130 133340 552180
rect 132960 552080 133340 552130
rect 133400 552270 133680 552320
rect 133400 552220 133470 552270
rect 133400 552180 133410 552220
rect 133450 552180 133470 552220
rect 133400 552130 133470 552180
rect 133500 552220 133680 552240
rect 133500 552180 133520 552220
rect 133660 552180 133680 552220
rect 133500 552160 133680 552180
rect 133710 552220 133780 552320
rect 133710 552180 133730 552220
rect 133770 552180 133780 552220
rect 133710 552130 133780 552180
rect 133400 552080 133780 552130
rect 124990 546450 125170 546500
rect 124990 546400 125060 546450
rect 124990 546360 125000 546400
rect 125040 546360 125060 546400
rect 124990 546310 125060 546360
rect 125090 546400 125170 546420
rect 125090 546360 125110 546400
rect 125150 546360 125170 546400
rect 125090 546340 125170 546360
rect 125200 546400 125270 546500
rect 125200 546360 125220 546400
rect 125260 546360 125270 546400
rect 125200 546310 125270 546360
rect 124990 546260 125270 546310
rect 119360 545780 119430 545800
rect 119360 545730 119370 545780
rect 119410 545730 119430 545780
rect 119360 545710 119430 545730
rect 119460 545780 119530 545800
rect 119460 545730 119480 545780
rect 119520 545730 119530 545780
rect 119460 545710 119530 545730
rect 119720 545580 119790 545600
rect 119720 545420 119730 545580
rect 119770 545420 119790 545580
rect 119720 545400 119790 545420
rect 119820 545580 119890 545600
rect 119820 545420 119840 545580
rect 119880 545420 119890 545580
rect 119820 545400 119890 545420
rect 120100 545580 120170 545600
rect 120100 545420 120110 545580
rect 120150 545420 120170 545580
rect 120100 545400 120170 545420
rect 120200 545580 120270 545600
rect 120200 545420 120220 545580
rect 120260 545420 120270 545580
rect 120200 545400 120270 545420
rect 125480 544700 125760 544750
rect 125480 544650 125550 544700
rect 125480 544410 125490 544650
rect 125530 544410 125550 544650
rect 125480 544360 125550 544410
rect 125580 544650 125760 544670
rect 125580 544410 125600 544650
rect 125740 544410 125760 544650
rect 125580 544390 125760 544410
rect 125790 544650 125860 544750
rect 125790 544410 125810 544650
rect 125850 544410 125860 544650
rect 125790 544360 125860 544410
rect 125480 544310 125860 544360
rect 125920 544700 126200 544750
rect 125920 544650 125990 544700
rect 125920 544410 125930 544650
rect 125970 544410 125990 544650
rect 125920 544360 125990 544410
rect 126020 544650 126200 544670
rect 126020 544410 126040 544650
rect 126180 544410 126200 544650
rect 126020 544390 126200 544410
rect 126230 544650 126300 544750
rect 126230 544410 126250 544650
rect 126290 544410 126300 544650
rect 126230 544360 126300 544410
rect 125920 544310 126300 544360
rect 126360 544700 126640 544750
rect 126360 544650 126430 544700
rect 126360 544410 126370 544650
rect 126410 544410 126430 544650
rect 126360 544360 126430 544410
rect 126460 544650 126640 544670
rect 126460 544410 126480 544650
rect 126620 544410 126640 544650
rect 126460 544390 126640 544410
rect 126670 544650 126740 544750
rect 126670 544410 126690 544650
rect 126730 544410 126740 544650
rect 126670 544360 126740 544410
rect 126360 544310 126740 544360
rect 126800 544700 127080 544750
rect 126800 544650 126870 544700
rect 126800 544410 126810 544650
rect 126850 544410 126870 544650
rect 126800 544360 126870 544410
rect 126900 544650 127080 544670
rect 126900 544410 126920 544650
rect 127060 544410 127080 544650
rect 126900 544390 127080 544410
rect 127110 544650 127180 544750
rect 127110 544410 127130 544650
rect 127170 544410 127180 544650
rect 127110 544360 127180 544410
rect 126800 544310 127180 544360
rect 127240 544700 127520 544750
rect 127240 544650 127310 544700
rect 127240 544410 127250 544650
rect 127290 544410 127310 544650
rect 127240 544360 127310 544410
rect 127340 544650 127520 544670
rect 127340 544410 127360 544650
rect 127500 544410 127520 544650
rect 127340 544390 127520 544410
rect 127550 544650 127620 544750
rect 127550 544410 127570 544650
rect 127610 544410 127620 544650
rect 127550 544360 127620 544410
rect 127240 544310 127620 544360
rect 127680 544700 127960 544750
rect 127680 544650 127750 544700
rect 127680 544410 127690 544650
rect 127730 544410 127750 544650
rect 127680 544360 127750 544410
rect 127780 544650 127960 544670
rect 127780 544410 127800 544650
rect 127940 544410 127960 544650
rect 127780 544390 127960 544410
rect 127990 544650 128060 544750
rect 127990 544410 128010 544650
rect 128050 544410 128060 544650
rect 127990 544360 128060 544410
rect 127680 544310 128060 544360
rect 128120 544700 128400 544750
rect 128120 544650 128190 544700
rect 128120 544410 128130 544650
rect 128170 544410 128190 544650
rect 128120 544360 128190 544410
rect 128220 544650 128400 544670
rect 128220 544410 128240 544650
rect 128380 544410 128400 544650
rect 128220 544390 128400 544410
rect 128430 544650 128500 544750
rect 128430 544410 128450 544650
rect 128490 544410 128500 544650
rect 128430 544360 128500 544410
rect 128120 544310 128500 544360
rect 128560 544700 128840 544750
rect 128560 544650 128630 544700
rect 128560 544410 128570 544650
rect 128610 544410 128630 544650
rect 128560 544360 128630 544410
rect 128660 544650 128840 544670
rect 128660 544410 128680 544650
rect 128820 544410 128840 544650
rect 128660 544390 128840 544410
rect 128870 544650 128940 544750
rect 128870 544410 128890 544650
rect 128930 544410 128940 544650
rect 128870 544360 128940 544410
rect 128560 544310 128940 544360
rect 129000 544700 129280 544750
rect 129000 544650 129070 544700
rect 129000 544410 129010 544650
rect 129050 544410 129070 544650
rect 129000 544360 129070 544410
rect 129100 544650 129280 544670
rect 129100 544410 129120 544650
rect 129260 544410 129280 544650
rect 129100 544390 129280 544410
rect 129310 544650 129380 544750
rect 129310 544410 129330 544650
rect 129370 544410 129380 544650
rect 129310 544360 129380 544410
rect 129000 544310 129380 544360
rect 129440 544700 129720 544750
rect 129440 544650 129510 544700
rect 129440 544410 129450 544650
rect 129490 544410 129510 544650
rect 129440 544360 129510 544410
rect 129540 544650 129720 544670
rect 129540 544410 129560 544650
rect 129700 544410 129720 544650
rect 129540 544390 129720 544410
rect 129750 544650 129820 544750
rect 129750 544410 129770 544650
rect 129810 544410 129820 544650
rect 129750 544360 129820 544410
rect 129440 544310 129820 544360
rect 129880 544700 130160 544750
rect 129880 544650 129950 544700
rect 129880 544410 129890 544650
rect 129930 544410 129950 544650
rect 129880 544360 129950 544410
rect 129980 544650 130160 544670
rect 129980 544410 130000 544650
rect 130140 544410 130160 544650
rect 129980 544390 130160 544410
rect 130190 544650 130260 544750
rect 130190 544410 130210 544650
rect 130250 544410 130260 544650
rect 130190 544360 130260 544410
rect 129880 544310 130260 544360
rect 130320 544700 130600 544750
rect 130320 544650 130390 544700
rect 130320 544410 130330 544650
rect 130370 544410 130390 544650
rect 130320 544360 130390 544410
rect 130420 544650 130600 544670
rect 130420 544410 130440 544650
rect 130580 544410 130600 544650
rect 130420 544390 130600 544410
rect 130630 544650 130700 544750
rect 130630 544410 130650 544650
rect 130690 544410 130700 544650
rect 130630 544360 130700 544410
rect 130320 544310 130700 544360
rect 130760 544700 131040 544750
rect 130760 544650 130830 544700
rect 130760 544410 130770 544650
rect 130810 544410 130830 544650
rect 130760 544360 130830 544410
rect 130860 544650 131040 544670
rect 130860 544410 130880 544650
rect 131020 544410 131040 544650
rect 130860 544390 131040 544410
rect 131070 544650 131140 544750
rect 131070 544410 131090 544650
rect 131130 544410 131140 544650
rect 131070 544360 131140 544410
rect 130760 544310 131140 544360
rect 131200 544700 131480 544750
rect 131200 544650 131270 544700
rect 131200 544410 131210 544650
rect 131250 544410 131270 544650
rect 131200 544360 131270 544410
rect 131300 544650 131480 544670
rect 131300 544410 131320 544650
rect 131460 544410 131480 544650
rect 131300 544390 131480 544410
rect 131510 544650 131580 544750
rect 131510 544410 131530 544650
rect 131570 544410 131580 544650
rect 131510 544360 131580 544410
rect 131200 544310 131580 544360
rect 131640 544700 131920 544750
rect 131640 544650 131710 544700
rect 131640 544410 131650 544650
rect 131690 544410 131710 544650
rect 131640 544360 131710 544410
rect 131740 544650 131920 544670
rect 131740 544410 131760 544650
rect 131900 544410 131920 544650
rect 131740 544390 131920 544410
rect 131950 544650 132020 544750
rect 131950 544410 131970 544650
rect 132010 544410 132020 544650
rect 131950 544360 132020 544410
rect 131640 544310 132020 544360
rect 132080 544700 132360 544750
rect 132080 544650 132150 544700
rect 132080 544410 132090 544650
rect 132130 544410 132150 544650
rect 132080 544360 132150 544410
rect 132180 544650 132360 544670
rect 132180 544410 132200 544650
rect 132340 544410 132360 544650
rect 132180 544390 132360 544410
rect 132390 544650 132460 544750
rect 132390 544410 132410 544650
rect 132450 544410 132460 544650
rect 132390 544360 132460 544410
rect 132080 544310 132460 544360
rect 132520 544700 132800 544750
rect 132520 544650 132590 544700
rect 132520 544410 132530 544650
rect 132570 544410 132590 544650
rect 132520 544360 132590 544410
rect 132620 544650 132800 544670
rect 132620 544410 132640 544650
rect 132780 544410 132800 544650
rect 132620 544390 132800 544410
rect 132830 544650 132900 544750
rect 132830 544410 132850 544650
rect 132890 544410 132900 544650
rect 132830 544360 132900 544410
rect 132520 544310 132900 544360
rect 132960 544700 133240 544750
rect 132960 544650 133030 544700
rect 132960 544410 132970 544650
rect 133010 544410 133030 544650
rect 132960 544360 133030 544410
rect 133060 544650 133240 544670
rect 133060 544410 133080 544650
rect 133220 544410 133240 544650
rect 133060 544390 133240 544410
rect 133270 544650 133340 544750
rect 133270 544410 133290 544650
rect 133330 544410 133340 544650
rect 133270 544360 133340 544410
rect 132960 544310 133340 544360
rect 133400 544700 133680 544750
rect 133400 544650 133470 544700
rect 133400 544410 133410 544650
rect 133450 544410 133470 544650
rect 133400 544360 133470 544410
rect 133500 544650 133680 544670
rect 133500 544410 133520 544650
rect 133660 544410 133680 544650
rect 133500 544390 133680 544410
rect 133710 544650 133780 544750
rect 133710 544410 133730 544650
rect 133770 544410 133780 544650
rect 133710 544360 133780 544410
rect 133400 544310 133780 544360
rect 124960 538390 125140 538440
rect 124960 538340 125030 538390
rect 124960 538300 124970 538340
rect 125010 538300 125030 538340
rect 124960 538250 125030 538300
rect 125060 538340 125140 538360
rect 125060 538300 125080 538340
rect 125120 538300 125140 538340
rect 125060 538280 125140 538300
rect 125170 538340 125240 538440
rect 125170 538300 125190 538340
rect 125230 538300 125240 538340
rect 125170 538250 125240 538300
rect 124960 538200 125240 538250
rect 119330 537720 119400 537740
rect 119330 537670 119340 537720
rect 119380 537670 119400 537720
rect 119330 537650 119400 537670
rect 119430 537720 119500 537740
rect 119430 537670 119450 537720
rect 119490 537670 119500 537720
rect 119430 537650 119500 537670
rect 119690 537520 119760 537540
rect 119690 537360 119700 537520
rect 119740 537360 119760 537520
rect 119690 537340 119760 537360
rect 119790 537520 119860 537540
rect 119790 537360 119810 537520
rect 119850 537360 119860 537520
rect 119790 537340 119860 537360
rect 120070 537520 120140 537540
rect 120070 537360 120080 537520
rect 120120 537360 120140 537520
rect 120070 537340 120140 537360
rect 120170 537520 120240 537540
rect 120170 537360 120190 537520
rect 120230 537360 120240 537520
rect 120170 537340 120240 537360
rect 125450 536640 125730 536690
rect 125450 536590 125520 536640
rect 125450 536150 125460 536590
rect 125500 536150 125520 536590
rect 125450 536100 125520 536150
rect 125550 536590 125730 536610
rect 125550 536150 125570 536590
rect 125710 536150 125730 536590
rect 125550 536130 125730 536150
rect 125760 536590 125830 536690
rect 125760 536150 125780 536590
rect 125820 536150 125830 536590
rect 125760 536100 125830 536150
rect 125450 536050 125830 536100
rect 125890 536640 126170 536690
rect 125890 536590 125960 536640
rect 125890 536150 125900 536590
rect 125940 536150 125960 536590
rect 125890 536100 125960 536150
rect 125990 536590 126170 536610
rect 125990 536150 126010 536590
rect 126150 536150 126170 536590
rect 125990 536130 126170 536150
rect 126200 536590 126270 536690
rect 126200 536150 126220 536590
rect 126260 536150 126270 536590
rect 126200 536100 126270 536150
rect 125890 536050 126270 536100
rect 126330 536640 126610 536690
rect 126330 536590 126400 536640
rect 126330 536150 126340 536590
rect 126380 536150 126400 536590
rect 126330 536100 126400 536150
rect 126430 536590 126610 536610
rect 126430 536150 126450 536590
rect 126590 536150 126610 536590
rect 126430 536130 126610 536150
rect 126640 536590 126710 536690
rect 126640 536150 126660 536590
rect 126700 536150 126710 536590
rect 126640 536100 126710 536150
rect 126330 536050 126710 536100
rect 126770 536640 127050 536690
rect 126770 536590 126840 536640
rect 126770 536150 126780 536590
rect 126820 536150 126840 536590
rect 126770 536100 126840 536150
rect 126870 536590 127050 536610
rect 126870 536150 126890 536590
rect 127030 536150 127050 536590
rect 126870 536130 127050 536150
rect 127080 536590 127150 536690
rect 127080 536150 127100 536590
rect 127140 536150 127150 536590
rect 127080 536100 127150 536150
rect 126770 536050 127150 536100
rect 127210 536640 127490 536690
rect 127210 536590 127280 536640
rect 127210 536150 127220 536590
rect 127260 536150 127280 536590
rect 127210 536100 127280 536150
rect 127310 536590 127490 536610
rect 127310 536150 127330 536590
rect 127470 536150 127490 536590
rect 127310 536130 127490 536150
rect 127520 536590 127590 536690
rect 127520 536150 127540 536590
rect 127580 536150 127590 536590
rect 127520 536100 127590 536150
rect 127210 536050 127590 536100
rect 127650 536640 127930 536690
rect 127650 536590 127720 536640
rect 127650 536150 127660 536590
rect 127700 536150 127720 536590
rect 127650 536100 127720 536150
rect 127750 536590 127930 536610
rect 127750 536150 127770 536590
rect 127910 536150 127930 536590
rect 127750 536130 127930 536150
rect 127960 536590 128030 536690
rect 127960 536150 127980 536590
rect 128020 536150 128030 536590
rect 127960 536100 128030 536150
rect 127650 536050 128030 536100
rect 128090 536640 128370 536690
rect 128090 536590 128160 536640
rect 128090 536150 128100 536590
rect 128140 536150 128160 536590
rect 128090 536100 128160 536150
rect 128190 536590 128370 536610
rect 128190 536150 128210 536590
rect 128350 536150 128370 536590
rect 128190 536130 128370 536150
rect 128400 536590 128470 536690
rect 128400 536150 128420 536590
rect 128460 536150 128470 536590
rect 128400 536100 128470 536150
rect 128090 536050 128470 536100
rect 128530 536640 128810 536690
rect 128530 536590 128600 536640
rect 128530 536150 128540 536590
rect 128580 536150 128600 536590
rect 128530 536100 128600 536150
rect 128630 536590 128810 536610
rect 128630 536150 128650 536590
rect 128790 536150 128810 536590
rect 128630 536130 128810 536150
rect 128840 536590 128910 536690
rect 128840 536150 128860 536590
rect 128900 536150 128910 536590
rect 128840 536100 128910 536150
rect 128530 536050 128910 536100
rect 128970 536640 129250 536690
rect 128970 536590 129040 536640
rect 128970 536150 128980 536590
rect 129020 536150 129040 536590
rect 128970 536100 129040 536150
rect 129070 536590 129250 536610
rect 129070 536150 129090 536590
rect 129230 536150 129250 536590
rect 129070 536130 129250 536150
rect 129280 536590 129350 536690
rect 129280 536150 129300 536590
rect 129340 536150 129350 536590
rect 129280 536100 129350 536150
rect 128970 536050 129350 536100
rect 129410 536640 129690 536690
rect 129410 536590 129480 536640
rect 129410 536150 129420 536590
rect 129460 536150 129480 536590
rect 129410 536100 129480 536150
rect 129510 536590 129690 536610
rect 129510 536150 129530 536590
rect 129670 536150 129690 536590
rect 129510 536130 129690 536150
rect 129720 536590 129790 536690
rect 129720 536150 129740 536590
rect 129780 536150 129790 536590
rect 129720 536100 129790 536150
rect 129410 536050 129790 536100
rect 129850 536640 130130 536690
rect 129850 536590 129920 536640
rect 129850 536150 129860 536590
rect 129900 536150 129920 536590
rect 129850 536100 129920 536150
rect 129950 536590 130130 536610
rect 129950 536150 129970 536590
rect 130110 536150 130130 536590
rect 129950 536130 130130 536150
rect 130160 536590 130230 536690
rect 130160 536150 130180 536590
rect 130220 536150 130230 536590
rect 130160 536100 130230 536150
rect 129850 536050 130230 536100
rect 130290 536640 130570 536690
rect 130290 536590 130360 536640
rect 130290 536150 130300 536590
rect 130340 536150 130360 536590
rect 130290 536100 130360 536150
rect 130390 536590 130570 536610
rect 130390 536150 130410 536590
rect 130550 536150 130570 536590
rect 130390 536130 130570 536150
rect 130600 536590 130670 536690
rect 130600 536150 130620 536590
rect 130660 536150 130670 536590
rect 130600 536100 130670 536150
rect 130290 536050 130670 536100
rect 130730 536640 131010 536690
rect 130730 536590 130800 536640
rect 130730 536150 130740 536590
rect 130780 536150 130800 536590
rect 130730 536100 130800 536150
rect 130830 536590 131010 536610
rect 130830 536150 130850 536590
rect 130990 536150 131010 536590
rect 130830 536130 131010 536150
rect 131040 536590 131110 536690
rect 131040 536150 131060 536590
rect 131100 536150 131110 536590
rect 131040 536100 131110 536150
rect 130730 536050 131110 536100
rect 131170 536640 131450 536690
rect 131170 536590 131240 536640
rect 131170 536150 131180 536590
rect 131220 536150 131240 536590
rect 131170 536100 131240 536150
rect 131270 536590 131450 536610
rect 131270 536150 131290 536590
rect 131430 536150 131450 536590
rect 131270 536130 131450 536150
rect 131480 536590 131550 536690
rect 131480 536150 131500 536590
rect 131540 536150 131550 536590
rect 131480 536100 131550 536150
rect 131170 536050 131550 536100
rect 131610 536640 131890 536690
rect 131610 536590 131680 536640
rect 131610 536150 131620 536590
rect 131660 536150 131680 536590
rect 131610 536100 131680 536150
rect 131710 536590 131890 536610
rect 131710 536150 131730 536590
rect 131870 536150 131890 536590
rect 131710 536130 131890 536150
rect 131920 536590 131990 536690
rect 131920 536150 131940 536590
rect 131980 536150 131990 536590
rect 131920 536100 131990 536150
rect 131610 536050 131990 536100
rect 132050 536640 132330 536690
rect 132050 536590 132120 536640
rect 132050 536150 132060 536590
rect 132100 536150 132120 536590
rect 132050 536100 132120 536150
rect 132150 536590 132330 536610
rect 132150 536150 132170 536590
rect 132310 536150 132330 536590
rect 132150 536130 132330 536150
rect 132360 536590 132430 536690
rect 132360 536150 132380 536590
rect 132420 536150 132430 536590
rect 132360 536100 132430 536150
rect 132050 536050 132430 536100
rect 132490 536640 132770 536690
rect 132490 536590 132560 536640
rect 132490 536150 132500 536590
rect 132540 536150 132560 536590
rect 132490 536100 132560 536150
rect 132590 536590 132770 536610
rect 132590 536150 132610 536590
rect 132750 536150 132770 536590
rect 132590 536130 132770 536150
rect 132800 536590 132870 536690
rect 132800 536150 132820 536590
rect 132860 536150 132870 536590
rect 132800 536100 132870 536150
rect 132490 536050 132870 536100
rect 132930 536640 133210 536690
rect 132930 536590 133000 536640
rect 132930 536150 132940 536590
rect 132980 536150 133000 536590
rect 132930 536100 133000 536150
rect 133030 536590 133210 536610
rect 133030 536150 133050 536590
rect 133190 536150 133210 536590
rect 133030 536130 133210 536150
rect 133240 536590 133310 536690
rect 133240 536150 133260 536590
rect 133300 536150 133310 536590
rect 133240 536100 133310 536150
rect 132930 536050 133310 536100
rect 133370 536640 133650 536690
rect 133370 536590 133440 536640
rect 133370 536150 133380 536590
rect 133420 536150 133440 536590
rect 133370 536100 133440 536150
rect 133470 536590 133650 536610
rect 133470 536150 133490 536590
rect 133630 536150 133650 536590
rect 133470 536130 133650 536150
rect 133680 536590 133750 536690
rect 133680 536150 133700 536590
rect 133740 536150 133750 536590
rect 133680 536100 133750 536150
rect 133370 536050 133750 536100
<< pdiff >>
rect 119620 593260 119690 593280
rect 119260 593230 119330 593250
rect 119260 593180 119270 593230
rect 119310 593180 119330 593230
rect 119260 593160 119330 593180
rect 119360 593230 119430 593250
rect 119360 593180 119380 593230
rect 119420 593180 119430 593230
rect 119360 593160 119430 593180
rect 119620 593100 119630 593260
rect 119670 593100 119690 593260
rect 119620 593080 119690 593100
rect 119720 593260 119790 593280
rect 119720 593100 119740 593260
rect 119780 593100 119790 593260
rect 119720 593080 119790 593100
rect 120000 593260 120070 593280
rect 120000 593100 120010 593260
rect 120050 593100 120070 593260
rect 120000 593080 120070 593100
rect 120100 593260 120170 593280
rect 120100 593100 120120 593260
rect 120160 593100 120170 593260
rect 120100 593080 120170 593100
rect 119660 583720 119730 583740
rect 119300 583690 119370 583710
rect 119300 583640 119310 583690
rect 119350 583640 119370 583690
rect 119300 583620 119370 583640
rect 119400 583690 119470 583710
rect 119400 583640 119420 583690
rect 119460 583640 119470 583690
rect 119400 583620 119470 583640
rect 119660 583560 119670 583720
rect 119710 583560 119730 583720
rect 119660 583540 119730 583560
rect 119760 583720 119830 583740
rect 119760 583560 119780 583720
rect 119820 583560 119830 583720
rect 119760 583540 119830 583560
rect 120040 583720 120110 583740
rect 120040 583560 120050 583720
rect 120090 583560 120110 583720
rect 120040 583540 120110 583560
rect 120140 583720 120210 583740
rect 120140 583560 120160 583720
rect 120200 583560 120210 583720
rect 120140 583540 120210 583560
rect 119700 574700 119770 574720
rect 119340 574670 119410 574690
rect 119340 574620 119350 574670
rect 119390 574620 119410 574670
rect 119340 574600 119410 574620
rect 119440 574670 119510 574690
rect 119440 574620 119460 574670
rect 119500 574620 119510 574670
rect 119440 574600 119510 574620
rect 119700 574540 119710 574700
rect 119750 574540 119770 574700
rect 119700 574520 119770 574540
rect 119800 574700 119870 574720
rect 119800 574540 119820 574700
rect 119860 574540 119870 574700
rect 119800 574520 119870 574540
rect 120080 574700 120150 574720
rect 120080 574540 120090 574700
rect 120130 574540 120150 574700
rect 120080 574520 120150 574540
rect 120180 574700 120250 574720
rect 120180 574540 120200 574700
rect 120240 574540 120250 574700
rect 120180 574520 120250 574540
rect 119650 567030 119720 567050
rect 119290 567000 119360 567020
rect 119290 566950 119300 567000
rect 119340 566950 119360 567000
rect 119290 566930 119360 566950
rect 119390 567000 119460 567020
rect 119390 566950 119410 567000
rect 119450 566950 119460 567000
rect 119390 566930 119460 566950
rect 119650 566870 119660 567030
rect 119700 566870 119720 567030
rect 119650 566850 119720 566870
rect 119750 567030 119820 567050
rect 119750 566870 119770 567030
rect 119810 566870 119820 567030
rect 119750 566850 119820 566870
rect 120030 567030 120100 567050
rect 120030 566870 120040 567030
rect 120080 566870 120100 567030
rect 120030 566850 120100 566870
rect 120130 567030 120200 567050
rect 120130 566870 120150 567030
rect 120190 566870 120200 567030
rect 120130 566850 120200 566870
rect 119650 560490 119720 560510
rect 119290 560460 119360 560480
rect 119290 560410 119300 560460
rect 119340 560410 119360 560460
rect 119290 560390 119360 560410
rect 119390 560460 119460 560480
rect 119390 560410 119410 560460
rect 119450 560410 119460 560460
rect 119390 560390 119460 560410
rect 119650 560330 119660 560490
rect 119700 560330 119720 560490
rect 119650 560310 119720 560330
rect 119750 560490 119820 560510
rect 119750 560330 119770 560490
rect 119810 560330 119820 560490
rect 119750 560310 119820 560330
rect 120030 560490 120100 560510
rect 120030 560330 120040 560490
rect 120080 560330 120100 560490
rect 120030 560310 120100 560330
rect 120130 560490 120200 560510
rect 120130 560330 120150 560490
rect 120190 560330 120200 560490
rect 120130 560310 120200 560330
rect 119720 553660 119790 553680
rect 119360 553630 119430 553650
rect 119360 553580 119370 553630
rect 119410 553580 119430 553630
rect 119360 553560 119430 553580
rect 119460 553630 119530 553650
rect 119460 553580 119480 553630
rect 119520 553580 119530 553630
rect 119460 553560 119530 553580
rect 119720 553500 119730 553660
rect 119770 553500 119790 553660
rect 119720 553480 119790 553500
rect 119820 553660 119890 553680
rect 119820 553500 119840 553660
rect 119880 553500 119890 553660
rect 119820 553480 119890 553500
rect 120100 553660 120170 553680
rect 120100 553500 120110 553660
rect 120150 553500 120170 553660
rect 120100 553480 120170 553500
rect 120200 553660 120270 553680
rect 120200 553500 120220 553660
rect 120260 553500 120270 553660
rect 120200 553480 120270 553500
rect 119720 546090 119790 546110
rect 119360 546060 119430 546080
rect 119360 546010 119370 546060
rect 119410 546010 119430 546060
rect 119360 545990 119430 546010
rect 119460 546060 119530 546080
rect 119460 546010 119480 546060
rect 119520 546010 119530 546060
rect 119460 545990 119530 546010
rect 119720 545930 119730 546090
rect 119770 545930 119790 546090
rect 119720 545910 119790 545930
rect 119820 546090 119890 546110
rect 119820 545930 119840 546090
rect 119880 545930 119890 546090
rect 119820 545910 119890 545930
rect 120100 546090 120170 546110
rect 120100 545930 120110 546090
rect 120150 545930 120170 546090
rect 120100 545910 120170 545930
rect 120200 546090 120270 546110
rect 120200 545930 120220 546090
rect 120260 545930 120270 546090
rect 120200 545910 120270 545930
rect 119690 538030 119760 538050
rect 119330 538000 119400 538020
rect 119330 537950 119340 538000
rect 119380 537950 119400 538000
rect 119330 537930 119400 537950
rect 119430 538000 119500 538020
rect 119430 537950 119450 538000
rect 119490 537950 119500 538000
rect 119430 537930 119500 537950
rect 119690 537870 119700 538030
rect 119740 537870 119760 538030
rect 119690 537850 119760 537870
rect 119790 538030 119860 538050
rect 119790 537870 119810 538030
rect 119850 537870 119860 538030
rect 119790 537850 119860 537870
rect 120070 538030 120140 538050
rect 120070 537870 120080 538030
rect 120120 537870 120140 538030
rect 120070 537850 120140 537870
rect 120170 538030 120240 538050
rect 120170 537870 120190 538030
rect 120230 537870 120240 538030
rect 120170 537850 120240 537870
<< ndiffc >>
rect 124170 642360 124220 642400
rect 124350 642360 124400 642400
rect 124530 642360 124580 642400
rect 124710 642360 124760 642400
rect 124890 642360 124940 642400
rect 125070 642360 125120 642400
rect 125250 642360 125300 642400
rect 125430 642360 125480 642400
rect 125610 642360 125660 642400
rect 125790 642360 125840 642400
rect 125970 642360 126020 642400
rect 126150 642360 126200 642400
rect 126330 642360 126380 642400
rect 126510 642360 126560 642400
rect 126690 642360 126740 642400
rect 126870 642360 126920 642400
rect 127050 642360 127100 642400
rect 127230 642360 127280 642400
rect 127410 642360 127460 642400
rect 127590 642360 127640 642400
rect 127770 642360 127820 642400
rect 127950 642360 128000 642400
rect 128130 642360 128180 642400
rect 128310 642360 128360 642400
rect 128490 642360 128540 642400
rect 128670 642360 128720 642400
rect 128850 642360 128900 642400
rect 129030 642360 129080 642400
rect 129210 642360 129260 642400
rect 129390 642360 129440 642400
rect 129570 642360 129620 642400
rect 129750 642360 129800 642400
rect 129930 642360 129980 642400
rect 130110 642360 130160 642400
rect 130290 642360 130340 642400
rect 130470 642360 130520 642400
rect 130650 642360 130700 642400
rect 130830 642360 130880 642400
rect 131010 642360 131060 642400
rect 131190 642360 131240 642400
rect 124170 642250 124220 642290
rect 124350 642250 124400 642290
rect 124530 642250 124580 642290
rect 124710 642250 124760 642290
rect 124890 642250 124940 642290
rect 125070 642250 125120 642290
rect 125250 642250 125300 642290
rect 125430 642250 125480 642290
rect 125610 642250 125660 642290
rect 125790 642250 125840 642290
rect 125970 642250 126020 642290
rect 126150 642250 126200 642290
rect 126330 642250 126380 642290
rect 126510 642250 126560 642290
rect 126690 642250 126740 642290
rect 126870 642250 126920 642290
rect 127050 642250 127100 642290
rect 127230 642250 127280 642290
rect 127410 642250 127460 642290
rect 127590 642250 127640 642290
rect 127770 642250 127820 642290
rect 127950 642250 128000 642290
rect 128130 642250 128180 642290
rect 128310 642250 128360 642290
rect 128490 642250 128540 642290
rect 128670 642250 128720 642290
rect 128850 642250 128900 642290
rect 129030 642250 129080 642290
rect 129210 642250 129260 642290
rect 129390 642250 129440 642290
rect 129570 642250 129620 642290
rect 129750 642250 129800 642290
rect 129930 642250 129980 642290
rect 130110 642250 130160 642290
rect 130290 642250 130340 642290
rect 130470 642250 130520 642290
rect 130650 642250 130700 642290
rect 130830 642250 130880 642290
rect 131010 642250 131060 642290
rect 131190 642250 131240 642290
rect 124200 636190 124340 636230
rect 124440 636190 124580 636230
rect 124680 636190 124820 636230
rect 124920 636190 125060 636230
rect 125160 636190 125300 636230
rect 125400 636190 125540 636230
rect 125640 636190 125780 636230
rect 125880 636190 126020 636230
rect 126120 636190 126260 636230
rect 126360 636190 126500 636230
rect 126600 636190 126740 636230
rect 126840 636190 126980 636230
rect 127080 636190 127220 636230
rect 127320 636190 127460 636230
rect 127560 636190 127700 636230
rect 127800 636190 127940 636230
rect 128040 636190 128180 636230
rect 128280 636190 128420 636230
rect 128520 636190 128660 636230
rect 128760 636190 128900 636230
rect 124200 636080 124340 636120
rect 124440 636080 124580 636120
rect 124680 636080 124820 636120
rect 124920 636080 125060 636120
rect 125160 636080 125300 636120
rect 125400 636080 125540 636120
rect 125640 636080 125780 636120
rect 125880 636080 126020 636120
rect 126120 636080 126260 636120
rect 126360 636080 126500 636120
rect 126600 636080 126740 636120
rect 126840 636080 126980 636120
rect 127080 636080 127220 636120
rect 127320 636080 127460 636120
rect 127560 636080 127700 636120
rect 127800 636080 127940 636120
rect 128040 636080 128180 636120
rect 128280 636080 128420 636120
rect 128520 636080 128660 636120
rect 128760 636080 128900 636120
rect 124260 632600 124620 632640
rect 124260 632490 124620 632530
rect 124470 630160 124830 630200
rect 124930 630160 125290 630200
rect 125390 630160 125750 630200
rect 125850 630160 126210 630200
rect 126310 630160 126670 630200
rect 126770 630160 127130 630200
rect 127230 630160 127590 630200
rect 127690 630160 128050 630200
rect 128150 630160 128510 630200
rect 128610 630160 128970 630200
rect 124470 630050 124830 630090
rect 124930 630050 125290 630090
rect 125390 630050 125750 630090
rect 125850 630050 126210 630090
rect 126310 630050 126670 630090
rect 126770 630050 127130 630090
rect 127230 630050 127590 630090
rect 127690 630050 128050 630090
rect 128150 630050 128510 630090
rect 128610 630050 128970 630090
rect 124240 624930 124800 624970
rect 124240 624820 124800 624860
rect 124800 623640 125360 623680
rect 125460 623640 126020 623680
rect 126120 623640 126680 623680
rect 126780 623640 127340 623680
rect 127440 623640 128000 623680
rect 128100 623640 128660 623680
rect 124800 623530 125360 623570
rect 125460 623530 126020 623570
rect 126120 623530 126680 623570
rect 126780 623530 127340 623570
rect 127440 623530 128000 623570
rect 128100 623530 128660 623570
rect 125360 619310 125400 619350
rect 125470 619310 125510 619350
rect 125580 619310 125620 619350
rect 125430 618530 125470 618570
rect 125540 618530 125580 618570
rect 125650 618530 125690 618570
rect 125770 618530 125810 618570
rect 125880 618530 125920 618570
rect 125990 618530 126030 618570
rect 126110 618530 126150 618570
rect 126220 618530 126260 618570
rect 126330 618530 126370 618570
rect 126450 618530 126490 618570
rect 126560 618530 126600 618570
rect 126670 618530 126710 618570
rect 126790 618530 126830 618570
rect 126900 618530 126940 618570
rect 127010 618530 127050 618570
rect 127130 618530 127170 618570
rect 127240 618530 127280 618570
rect 127350 618530 127390 618570
rect 127470 618530 127510 618570
rect 127580 618530 127620 618570
rect 127690 618530 127730 618570
rect 127810 618530 127850 618570
rect 127920 618530 127960 618570
rect 128030 618530 128070 618570
rect 128150 618530 128190 618570
rect 128260 618530 128300 618570
rect 128370 618530 128410 618570
rect 128490 618530 128530 618570
rect 128600 618530 128640 618570
rect 128710 618530 128750 618570
rect 128830 618530 128870 618570
rect 128940 618530 128980 618570
rect 129050 618530 129090 618570
rect 129170 618530 129210 618570
rect 129280 618530 129320 618570
rect 129390 618530 129430 618570
rect 129510 618530 129550 618570
rect 129620 618530 129660 618570
rect 129730 618530 129770 618570
rect 129850 618530 129890 618570
rect 129960 618530 130000 618570
rect 130070 618530 130110 618570
rect 130190 618530 130230 618570
rect 130300 618530 130340 618570
rect 130410 618530 130450 618570
rect 130530 618530 130570 618570
rect 130640 618530 130680 618570
rect 130750 618530 130790 618570
rect 130870 618530 130910 618570
rect 130980 618530 131020 618570
rect 131090 618530 131130 618570
rect 131210 618530 131250 618570
rect 131320 618530 131360 618570
rect 131430 618530 131470 618570
rect 131550 618530 131590 618570
rect 131660 618530 131700 618570
rect 131770 618530 131810 618570
rect 125010 611860 125050 611900
rect 125120 611860 125160 611900
rect 125230 611860 125270 611900
rect 125080 610930 125120 611120
rect 125190 610930 125230 611120
rect 125300 610930 125340 611120
rect 125420 610930 125460 611120
rect 125530 610930 125570 611120
rect 125640 610930 125680 611120
rect 125760 610930 125800 611120
rect 125870 610930 125910 611120
rect 125980 610930 126020 611120
rect 126100 610930 126140 611120
rect 126210 610930 126250 611120
rect 126320 610930 126360 611120
rect 126440 610930 126480 611120
rect 126550 610930 126590 611120
rect 126660 610930 126700 611120
rect 126780 610930 126820 611120
rect 126890 610930 126930 611120
rect 127000 610930 127040 611120
rect 127120 610930 127160 611120
rect 127230 610930 127270 611120
rect 127340 610930 127380 611120
rect 127460 610930 127500 611120
rect 127570 610930 127610 611120
rect 127680 610930 127720 611120
rect 127800 610930 127840 611120
rect 127910 610930 127950 611120
rect 128020 610930 128060 611120
rect 128140 610930 128180 611120
rect 128250 610930 128290 611120
rect 128360 610930 128400 611120
rect 128480 610930 128520 611120
rect 128590 610930 128630 611120
rect 128700 610930 128740 611120
rect 128820 610930 128860 611120
rect 128930 610930 128970 611120
rect 129040 610930 129080 611120
rect 129160 610930 129200 611120
rect 129270 610930 129310 611120
rect 129380 610930 129420 611120
rect 129500 610930 129540 611120
rect 129610 610930 129650 611120
rect 129720 610930 129760 611120
rect 129840 610930 129880 611120
rect 129950 610930 129990 611120
rect 130060 610930 130100 611120
rect 130180 610930 130220 611120
rect 130290 610930 130330 611120
rect 130400 610930 130440 611120
rect 130520 610930 130560 611120
rect 130630 610930 130670 611120
rect 130740 610930 130780 611120
rect 130860 610930 130900 611120
rect 130970 610930 131010 611120
rect 131080 610930 131120 611120
rect 131200 610930 131240 611120
rect 131310 610930 131350 611120
rect 131420 610930 131460 611120
rect 125140 605810 125180 605850
rect 125250 605810 125290 605850
rect 125360 605810 125400 605850
rect 125210 604780 125250 605070
rect 125320 604780 125360 605070
rect 125430 604780 125470 605070
rect 125550 604780 125590 605070
rect 125660 604780 125700 605070
rect 125770 604780 125810 605070
rect 125890 604780 125930 605070
rect 126000 604780 126040 605070
rect 126110 604780 126150 605070
rect 126230 604780 126270 605070
rect 126340 604780 126380 605070
rect 126450 604780 126490 605070
rect 126570 604780 126610 605070
rect 126680 604780 126720 605070
rect 126790 604780 126830 605070
rect 126910 604780 126950 605070
rect 127020 604780 127060 605070
rect 127130 604780 127170 605070
rect 127250 604780 127290 605070
rect 127360 604780 127400 605070
rect 127470 604780 127510 605070
rect 127590 604780 127630 605070
rect 127700 604780 127740 605070
rect 127810 604780 127850 605070
rect 127930 604780 127970 605070
rect 128040 604780 128080 605070
rect 128150 604780 128190 605070
rect 128270 604780 128310 605070
rect 128380 604780 128420 605070
rect 128490 604780 128530 605070
rect 128610 604780 128650 605070
rect 128720 604780 128760 605070
rect 128830 604780 128870 605070
rect 128950 604780 128990 605070
rect 129060 604780 129100 605070
rect 129170 604780 129210 605070
rect 129290 604780 129330 605070
rect 129400 604780 129440 605070
rect 129510 604780 129550 605070
rect 129630 604780 129670 605070
rect 129740 604780 129780 605070
rect 129850 604780 129890 605070
rect 129970 604780 130010 605070
rect 130080 604780 130120 605070
rect 130190 604780 130230 605070
rect 130310 604780 130350 605070
rect 130420 604780 130460 605070
rect 130530 604780 130570 605070
rect 130650 604780 130690 605070
rect 130760 604780 130800 605070
rect 130870 604780 130910 605070
rect 130990 604780 131030 605070
rect 131100 604780 131140 605070
rect 131210 604780 131250 605070
rect 131330 604780 131370 605070
rect 131440 604780 131480 605070
rect 131550 604780 131590 605070
rect 124940 599550 124980 599590
rect 125050 599550 125090 599590
rect 125160 599550 125200 599590
rect 125010 598420 125050 598810
rect 125120 598420 125160 598810
rect 125230 598420 125270 598810
rect 125350 598420 125390 598810
rect 125460 598420 125500 598810
rect 125570 598420 125610 598810
rect 125690 598420 125730 598810
rect 125800 598420 125840 598810
rect 125910 598420 125950 598810
rect 126030 598420 126070 598810
rect 126140 598420 126180 598810
rect 126250 598420 126290 598810
rect 126370 598420 126410 598810
rect 126480 598420 126520 598810
rect 126590 598420 126630 598810
rect 126710 598420 126750 598810
rect 126820 598420 126860 598810
rect 126930 598420 126970 598810
rect 127050 598420 127090 598810
rect 127160 598420 127200 598810
rect 127270 598420 127310 598810
rect 127390 598420 127430 598810
rect 127500 598420 127540 598810
rect 127610 598420 127650 598810
rect 127730 598420 127770 598810
rect 127840 598420 127880 598810
rect 127950 598420 127990 598810
rect 128070 598420 128110 598810
rect 128180 598420 128220 598810
rect 128290 598420 128330 598810
rect 128410 598420 128450 598810
rect 128520 598420 128560 598810
rect 128630 598420 128670 598810
rect 128750 598420 128790 598810
rect 128860 598420 128900 598810
rect 128970 598420 129010 598810
rect 129090 598420 129130 598810
rect 129200 598420 129240 598810
rect 129310 598420 129350 598810
rect 129430 598420 129470 598810
rect 129540 598420 129580 598810
rect 129650 598420 129690 598810
rect 129770 598420 129810 598810
rect 129880 598420 129920 598810
rect 129990 598420 130030 598810
rect 130110 598420 130150 598810
rect 130220 598420 130260 598810
rect 130330 598420 130370 598810
rect 130450 598420 130490 598810
rect 130560 598420 130600 598810
rect 130670 598420 130710 598810
rect 130790 598420 130830 598810
rect 130900 598420 130940 598810
rect 131010 598420 131050 598810
rect 131130 598420 131170 598810
rect 131240 598420 131280 598810
rect 131350 598420 131390 598810
rect 119270 592900 119310 592950
rect 119380 592900 119420 592950
rect 119630 592590 119670 592750
rect 119740 592590 119780 592750
rect 120010 592590 120050 592750
rect 120120 592590 120160 592750
rect 124900 592000 124940 592040
rect 125010 592000 125050 592040
rect 125120 592000 125160 592040
rect 124970 590770 125010 591260
rect 125080 590770 125120 591260
rect 125190 590770 125230 591260
rect 125310 590770 125350 591260
rect 125420 590770 125460 591260
rect 125530 590770 125570 591260
rect 125650 590770 125690 591260
rect 125760 590770 125800 591260
rect 125870 590770 125910 591260
rect 125990 590770 126030 591260
rect 126100 590770 126140 591260
rect 126210 590770 126250 591260
rect 126330 590770 126370 591260
rect 126440 590770 126480 591260
rect 126550 590770 126590 591260
rect 126670 590770 126710 591260
rect 126780 590770 126820 591260
rect 126890 590770 126930 591260
rect 127010 590770 127050 591260
rect 127120 590770 127160 591260
rect 127230 590770 127270 591260
rect 127350 590770 127390 591260
rect 127460 590770 127500 591260
rect 127570 590770 127610 591260
rect 127690 590770 127730 591260
rect 127800 590770 127840 591260
rect 127910 590770 127950 591260
rect 128030 590770 128070 591260
rect 128140 590770 128180 591260
rect 128250 590770 128290 591260
rect 128370 590770 128410 591260
rect 128480 590770 128520 591260
rect 128590 590770 128630 591260
rect 128710 590770 128750 591260
rect 128820 590770 128860 591260
rect 128930 590770 128970 591260
rect 129050 590770 129090 591260
rect 129160 590770 129200 591260
rect 129270 590770 129310 591260
rect 129390 590770 129430 591260
rect 129500 590770 129540 591260
rect 129610 590770 129650 591260
rect 129730 590770 129770 591260
rect 129840 590770 129880 591260
rect 129950 590770 129990 591260
rect 130070 590770 130110 591260
rect 130180 590770 130220 591260
rect 130290 590770 130330 591260
rect 130410 590770 130450 591260
rect 130520 590770 130560 591260
rect 130630 590770 130670 591260
rect 130750 590770 130790 591260
rect 130860 590770 130900 591260
rect 130970 590770 131010 591260
rect 131090 590770 131130 591260
rect 131200 590770 131240 591260
rect 131310 590770 131350 591260
rect 119310 583360 119350 583410
rect 119420 583360 119460 583410
rect 119670 583050 119710 583210
rect 119780 583050 119820 583210
rect 120050 583050 120090 583210
rect 120160 583050 120200 583210
rect 125360 583020 125400 583060
rect 125470 583020 125510 583060
rect 125580 583020 125620 583060
rect 125430 582240 125470 582280
rect 125540 582240 125630 582280
rect 125700 582240 125740 582280
rect 125820 582240 125860 582280
rect 125930 582240 126020 582280
rect 126090 582240 126130 582280
rect 126210 582240 126250 582280
rect 126320 582240 126410 582280
rect 126480 582240 126520 582280
rect 126600 582240 126640 582280
rect 126710 582240 126800 582280
rect 126870 582240 126910 582280
rect 126990 582240 127030 582280
rect 127100 582240 127190 582280
rect 127260 582240 127300 582280
rect 127380 582240 127420 582280
rect 127490 582240 127580 582280
rect 127650 582240 127690 582280
rect 127770 582240 127810 582280
rect 127880 582240 127970 582280
rect 128040 582240 128080 582280
rect 128160 582240 128200 582280
rect 128270 582240 128360 582280
rect 128430 582240 128470 582280
rect 128550 582240 128590 582280
rect 128660 582240 128750 582280
rect 128820 582240 128860 582280
rect 128940 582240 128980 582280
rect 129050 582240 129140 582280
rect 129210 582240 129250 582280
rect 129330 582240 129370 582280
rect 129440 582240 129530 582280
rect 129600 582240 129640 582280
rect 129720 582240 129760 582280
rect 129830 582240 129920 582280
rect 129990 582240 130030 582280
rect 130110 582240 130150 582280
rect 130220 582240 130310 582280
rect 130380 582240 130420 582280
rect 130500 582240 130540 582280
rect 130610 582240 130700 582280
rect 130770 582240 130810 582280
rect 130890 582240 130930 582280
rect 131000 582240 131090 582280
rect 131160 582240 131200 582280
rect 131280 582240 131320 582280
rect 131390 582240 131480 582280
rect 131550 582240 131590 582280
rect 131670 582240 131710 582280
rect 131780 582240 131870 582280
rect 131940 582240 131980 582280
rect 132060 582240 132100 582280
rect 132170 582240 132260 582280
rect 132330 582240 132370 582280
rect 132450 582240 132490 582280
rect 132560 582240 132650 582280
rect 132720 582240 132760 582280
rect 119350 574340 119390 574390
rect 119460 574340 119500 574390
rect 119710 574030 119750 574190
rect 119820 574030 119860 574190
rect 120090 574030 120130 574190
rect 120200 574030 120240 574190
rect 125400 574000 125440 574040
rect 125510 574000 125550 574040
rect 125620 574000 125660 574040
rect 125470 573120 125510 573260
rect 125580 573120 125670 573260
rect 125740 573120 125780 573260
rect 125860 573120 125900 573260
rect 125970 573120 126060 573260
rect 126130 573120 126170 573260
rect 126250 573120 126290 573260
rect 126360 573120 126450 573260
rect 126520 573120 126560 573260
rect 126640 573120 126680 573260
rect 126750 573120 126840 573260
rect 126910 573120 126950 573260
rect 127030 573120 127070 573260
rect 127140 573120 127230 573260
rect 127300 573120 127340 573260
rect 127420 573120 127460 573260
rect 127530 573120 127620 573260
rect 127690 573120 127730 573260
rect 127810 573120 127850 573260
rect 127920 573120 128010 573260
rect 128080 573120 128120 573260
rect 128200 573120 128240 573260
rect 128310 573120 128400 573260
rect 128470 573120 128510 573260
rect 128590 573120 128630 573260
rect 128700 573120 128790 573260
rect 128860 573120 128900 573260
rect 128980 573120 129020 573260
rect 129090 573120 129180 573260
rect 129250 573120 129290 573260
rect 129370 573120 129410 573260
rect 129480 573120 129570 573260
rect 129640 573120 129680 573260
rect 129760 573120 129800 573260
rect 129870 573120 129960 573260
rect 130030 573120 130070 573260
rect 130150 573120 130190 573260
rect 130260 573120 130350 573260
rect 130420 573120 130460 573260
rect 130540 573120 130580 573260
rect 130650 573120 130740 573260
rect 130810 573120 130850 573260
rect 130930 573120 130970 573260
rect 131040 573120 131130 573260
rect 131200 573120 131240 573260
rect 131320 573120 131360 573260
rect 131430 573120 131520 573260
rect 131590 573120 131630 573260
rect 131710 573120 131750 573260
rect 131820 573120 131910 573260
rect 131980 573120 132020 573260
rect 132100 573120 132140 573260
rect 132210 573120 132300 573260
rect 132370 573120 132410 573260
rect 132490 573120 132530 573260
rect 132600 573120 132690 573260
rect 132760 573120 132800 573260
rect 119300 566670 119340 566720
rect 119410 566670 119450 566720
rect 119660 566360 119700 566520
rect 119770 566360 119810 566520
rect 120040 566360 120080 566520
rect 120150 566360 120190 566520
rect 125350 566330 125390 566370
rect 125460 566330 125500 566370
rect 125570 566330 125610 566370
rect 125420 565350 125460 565590
rect 125530 565350 125620 565590
rect 125690 565350 125730 565590
rect 125810 565350 125850 565590
rect 125920 565350 126010 565590
rect 126080 565350 126120 565590
rect 126200 565350 126240 565590
rect 126310 565350 126400 565590
rect 126470 565350 126510 565590
rect 126590 565350 126630 565590
rect 126700 565350 126790 565590
rect 126860 565350 126900 565590
rect 126980 565350 127020 565590
rect 127090 565350 127180 565590
rect 127250 565350 127290 565590
rect 127370 565350 127410 565590
rect 127480 565350 127570 565590
rect 127640 565350 127680 565590
rect 127760 565350 127800 565590
rect 127870 565350 127960 565590
rect 128030 565350 128070 565590
rect 128150 565350 128190 565590
rect 128260 565350 128350 565590
rect 128420 565350 128460 565590
rect 128540 565350 128580 565590
rect 128650 565350 128740 565590
rect 128810 565350 128850 565590
rect 128930 565350 128970 565590
rect 129040 565350 129130 565590
rect 129200 565350 129240 565590
rect 129320 565350 129360 565590
rect 129430 565350 129520 565590
rect 129590 565350 129630 565590
rect 129710 565350 129750 565590
rect 129820 565350 129910 565590
rect 129980 565350 130020 565590
rect 130100 565350 130140 565590
rect 130210 565350 130300 565590
rect 130370 565350 130410 565590
rect 130490 565350 130530 565590
rect 130600 565350 130690 565590
rect 130760 565350 130800 565590
rect 130880 565350 130920 565590
rect 130990 565350 131080 565590
rect 131150 565350 131190 565590
rect 131270 565350 131310 565590
rect 131380 565350 131470 565590
rect 131540 565350 131580 565590
rect 131660 565350 131700 565590
rect 131770 565350 131860 565590
rect 131930 565350 131970 565590
rect 132050 565350 132090 565590
rect 132160 565350 132250 565590
rect 132320 565350 132360 565590
rect 132440 565350 132480 565590
rect 132550 565350 132640 565590
rect 132710 565350 132750 565590
rect 119300 560130 119340 560180
rect 119410 560130 119450 560180
rect 119660 559820 119700 559980
rect 119770 559820 119810 559980
rect 120040 559820 120080 559980
rect 120150 559820 120190 559980
rect 125350 559790 125390 559830
rect 125460 559790 125500 559830
rect 125570 559790 125610 559830
rect 125420 558710 125460 559050
rect 125530 558710 125620 559050
rect 125690 558710 125730 559050
rect 125810 558710 125850 559050
rect 125920 558710 126010 559050
rect 126080 558710 126120 559050
rect 126200 558710 126240 559050
rect 126310 558710 126400 559050
rect 126470 558710 126510 559050
rect 126590 558710 126630 559050
rect 126700 558710 126790 559050
rect 126860 558710 126900 559050
rect 126980 558710 127020 559050
rect 127090 558710 127180 559050
rect 127250 558710 127290 559050
rect 127370 558710 127410 559050
rect 127480 558710 127570 559050
rect 127640 558710 127680 559050
rect 127760 558710 127800 559050
rect 127870 558710 127960 559050
rect 128030 558710 128070 559050
rect 128150 558710 128190 559050
rect 128260 558710 128350 559050
rect 128420 558710 128460 559050
rect 128540 558710 128580 559050
rect 128650 558710 128740 559050
rect 128810 558710 128850 559050
rect 128930 558710 128970 559050
rect 129040 558710 129130 559050
rect 129200 558710 129240 559050
rect 129320 558710 129360 559050
rect 129430 558710 129520 559050
rect 129590 558710 129630 559050
rect 129710 558710 129750 559050
rect 129820 558710 129910 559050
rect 129980 558710 130020 559050
rect 130100 558710 130140 559050
rect 130210 558710 130300 559050
rect 130370 558710 130410 559050
rect 130490 558710 130530 559050
rect 130600 558710 130690 559050
rect 130760 558710 130800 559050
rect 130880 558710 130920 559050
rect 130990 558710 131080 559050
rect 131150 558710 131190 559050
rect 131270 558710 131310 559050
rect 131380 558710 131470 559050
rect 131540 558710 131580 559050
rect 131660 558710 131700 559050
rect 131770 558710 131860 559050
rect 131930 558710 131970 559050
rect 132050 558710 132090 559050
rect 132160 558710 132250 559050
rect 132320 558710 132360 559050
rect 132440 558710 132480 559050
rect 132550 558710 132640 559050
rect 132710 558710 132750 559050
rect 125000 553930 125040 553970
rect 125110 553930 125150 553970
rect 125220 553930 125260 553970
rect 119370 553300 119410 553350
rect 119480 553300 119520 553350
rect 119730 552990 119770 553150
rect 119840 552990 119880 553150
rect 120110 552990 120150 553150
rect 120220 552990 120260 553150
rect 125490 552180 125530 552220
rect 125600 552180 125740 552220
rect 125810 552180 125850 552220
rect 125930 552180 125970 552220
rect 126040 552180 126180 552220
rect 126250 552180 126290 552220
rect 126370 552180 126410 552220
rect 126480 552180 126620 552220
rect 126690 552180 126730 552220
rect 126810 552180 126850 552220
rect 126920 552180 127060 552220
rect 127130 552180 127170 552220
rect 127250 552180 127290 552220
rect 127360 552180 127500 552220
rect 127570 552180 127610 552220
rect 127690 552180 127730 552220
rect 127800 552180 127940 552220
rect 128010 552180 128050 552220
rect 128130 552180 128170 552220
rect 128240 552180 128380 552220
rect 128450 552180 128490 552220
rect 128570 552180 128610 552220
rect 128680 552180 128820 552220
rect 128890 552180 128930 552220
rect 129010 552180 129050 552220
rect 129120 552180 129260 552220
rect 129330 552180 129370 552220
rect 129450 552180 129490 552220
rect 129560 552180 129700 552220
rect 129770 552180 129810 552220
rect 129890 552180 129930 552220
rect 130000 552180 130140 552220
rect 130210 552180 130250 552220
rect 130330 552180 130370 552220
rect 130440 552180 130580 552220
rect 130650 552180 130690 552220
rect 130770 552180 130810 552220
rect 130880 552180 131020 552220
rect 131090 552180 131130 552220
rect 131210 552180 131250 552220
rect 131320 552180 131460 552220
rect 131530 552180 131570 552220
rect 131650 552180 131690 552220
rect 131760 552180 131900 552220
rect 131970 552180 132010 552220
rect 132090 552180 132130 552220
rect 132200 552180 132340 552220
rect 132410 552180 132450 552220
rect 132530 552180 132570 552220
rect 132640 552180 132780 552220
rect 132850 552180 132890 552220
rect 132970 552180 133010 552220
rect 133080 552180 133220 552220
rect 133290 552180 133330 552220
rect 133410 552180 133450 552220
rect 133520 552180 133660 552220
rect 133730 552180 133770 552220
rect 125000 546360 125040 546400
rect 125110 546360 125150 546400
rect 125220 546360 125260 546400
rect 119370 545730 119410 545780
rect 119480 545730 119520 545780
rect 119730 545420 119770 545580
rect 119840 545420 119880 545580
rect 120110 545420 120150 545580
rect 120220 545420 120260 545580
rect 125490 544410 125530 544650
rect 125600 544410 125740 544650
rect 125810 544410 125850 544650
rect 125930 544410 125970 544650
rect 126040 544410 126180 544650
rect 126250 544410 126290 544650
rect 126370 544410 126410 544650
rect 126480 544410 126620 544650
rect 126690 544410 126730 544650
rect 126810 544410 126850 544650
rect 126920 544410 127060 544650
rect 127130 544410 127170 544650
rect 127250 544410 127290 544650
rect 127360 544410 127500 544650
rect 127570 544410 127610 544650
rect 127690 544410 127730 544650
rect 127800 544410 127940 544650
rect 128010 544410 128050 544650
rect 128130 544410 128170 544650
rect 128240 544410 128380 544650
rect 128450 544410 128490 544650
rect 128570 544410 128610 544650
rect 128680 544410 128820 544650
rect 128890 544410 128930 544650
rect 129010 544410 129050 544650
rect 129120 544410 129260 544650
rect 129330 544410 129370 544650
rect 129450 544410 129490 544650
rect 129560 544410 129700 544650
rect 129770 544410 129810 544650
rect 129890 544410 129930 544650
rect 130000 544410 130140 544650
rect 130210 544410 130250 544650
rect 130330 544410 130370 544650
rect 130440 544410 130580 544650
rect 130650 544410 130690 544650
rect 130770 544410 130810 544650
rect 130880 544410 131020 544650
rect 131090 544410 131130 544650
rect 131210 544410 131250 544650
rect 131320 544410 131460 544650
rect 131530 544410 131570 544650
rect 131650 544410 131690 544650
rect 131760 544410 131900 544650
rect 131970 544410 132010 544650
rect 132090 544410 132130 544650
rect 132200 544410 132340 544650
rect 132410 544410 132450 544650
rect 132530 544410 132570 544650
rect 132640 544410 132780 544650
rect 132850 544410 132890 544650
rect 132970 544410 133010 544650
rect 133080 544410 133220 544650
rect 133290 544410 133330 544650
rect 133410 544410 133450 544650
rect 133520 544410 133660 544650
rect 133730 544410 133770 544650
rect 124970 538300 125010 538340
rect 125080 538300 125120 538340
rect 125190 538300 125230 538340
rect 119340 537670 119380 537720
rect 119450 537670 119490 537720
rect 119700 537360 119740 537520
rect 119810 537360 119850 537520
rect 120080 537360 120120 537520
rect 120190 537360 120230 537520
rect 125460 536150 125500 536590
rect 125570 536150 125710 536590
rect 125780 536150 125820 536590
rect 125900 536150 125940 536590
rect 126010 536150 126150 536590
rect 126220 536150 126260 536590
rect 126340 536150 126380 536590
rect 126450 536150 126590 536590
rect 126660 536150 126700 536590
rect 126780 536150 126820 536590
rect 126890 536150 127030 536590
rect 127100 536150 127140 536590
rect 127220 536150 127260 536590
rect 127330 536150 127470 536590
rect 127540 536150 127580 536590
rect 127660 536150 127700 536590
rect 127770 536150 127910 536590
rect 127980 536150 128020 536590
rect 128100 536150 128140 536590
rect 128210 536150 128350 536590
rect 128420 536150 128460 536590
rect 128540 536150 128580 536590
rect 128650 536150 128790 536590
rect 128860 536150 128900 536590
rect 128980 536150 129020 536590
rect 129090 536150 129230 536590
rect 129300 536150 129340 536590
rect 129420 536150 129460 536590
rect 129530 536150 129670 536590
rect 129740 536150 129780 536590
rect 129860 536150 129900 536590
rect 129970 536150 130110 536590
rect 130180 536150 130220 536590
rect 130300 536150 130340 536590
rect 130410 536150 130550 536590
rect 130620 536150 130660 536590
rect 130740 536150 130780 536590
rect 130850 536150 130990 536590
rect 131060 536150 131100 536590
rect 131180 536150 131220 536590
rect 131290 536150 131430 536590
rect 131500 536150 131540 536590
rect 131620 536150 131660 536590
rect 131730 536150 131870 536590
rect 131940 536150 131980 536590
rect 132060 536150 132100 536590
rect 132170 536150 132310 536590
rect 132380 536150 132420 536590
rect 132500 536150 132540 536590
rect 132610 536150 132750 536590
rect 132820 536150 132860 536590
rect 132940 536150 132980 536590
rect 133050 536150 133190 536590
rect 133260 536150 133300 536590
rect 133380 536150 133420 536590
rect 133490 536150 133630 536590
rect 133700 536150 133740 536590
<< pdiffc >>
rect 119270 593180 119310 593230
rect 119380 593180 119420 593230
rect 119630 593100 119670 593260
rect 119740 593100 119780 593260
rect 120010 593100 120050 593260
rect 120120 593100 120160 593260
rect 119310 583640 119350 583690
rect 119420 583640 119460 583690
rect 119670 583560 119710 583720
rect 119780 583560 119820 583720
rect 120050 583560 120090 583720
rect 120160 583560 120200 583720
rect 119350 574620 119390 574670
rect 119460 574620 119500 574670
rect 119710 574540 119750 574700
rect 119820 574540 119860 574700
rect 120090 574540 120130 574700
rect 120200 574540 120240 574700
rect 119300 566950 119340 567000
rect 119410 566950 119450 567000
rect 119660 566870 119700 567030
rect 119770 566870 119810 567030
rect 120040 566870 120080 567030
rect 120150 566870 120190 567030
rect 119300 560410 119340 560460
rect 119410 560410 119450 560460
rect 119660 560330 119700 560490
rect 119770 560330 119810 560490
rect 120040 560330 120080 560490
rect 120150 560330 120190 560490
rect 119370 553580 119410 553630
rect 119480 553580 119520 553630
rect 119730 553500 119770 553660
rect 119840 553500 119880 553660
rect 120110 553500 120150 553660
rect 120220 553500 120260 553660
rect 119370 546010 119410 546060
rect 119480 546010 119520 546060
rect 119730 545930 119770 546090
rect 119840 545930 119880 546090
rect 120110 545930 120150 546090
rect 120220 545930 120260 546090
rect 119340 537950 119380 538000
rect 119450 537950 119490 538000
rect 119700 537870 119740 538030
rect 119810 537870 119850 538030
rect 120080 537870 120120 538030
rect 120190 537870 120230 538030
<< psubdiff >>
rect 123830 643020 131630 643040
rect 123830 642900 123870 643020
rect 124000 642900 124110 643020
rect 124240 642900 124410 643020
rect 124540 642900 124710 643020
rect 124840 642900 125010 643020
rect 125140 642900 125310 643020
rect 125440 642900 125610 643020
rect 125740 642900 125910 643020
rect 126040 642900 126210 643020
rect 126340 642900 126510 643020
rect 126640 642900 126810 643020
rect 126940 642900 127110 643020
rect 127240 642900 127410 643020
rect 127540 642900 127710 643020
rect 127840 642900 128010 643020
rect 128140 642900 128310 643020
rect 128440 642900 128610 643020
rect 128740 642900 128910 643020
rect 129040 642900 129210 643020
rect 129340 642900 129510 643020
rect 129640 642900 129810 643020
rect 129940 642900 130110 643020
rect 130240 642900 130410 643020
rect 130540 642900 130710 643020
rect 130840 642900 131010 643020
rect 131140 642900 131310 643020
rect 131440 642900 131630 643020
rect 123830 642820 123960 642900
rect 131500 642810 131630 642900
rect 123830 642610 123960 642700
rect 131500 642630 131630 642690
rect 123830 641930 123960 642040
rect 123830 641760 123960 641810
rect 131500 641760 131630 642060
rect 123830 641640 123980 641760
rect 124110 641640 124280 641760
rect 124410 641640 124580 641760
rect 124710 641640 124880 641760
rect 125010 641640 125180 641760
rect 125310 641640 125480 641760
rect 125610 641640 125780 641760
rect 125910 641640 126080 641760
rect 126210 641640 126380 641760
rect 126510 641640 126680 641760
rect 126810 641640 126980 641760
rect 127110 641640 127280 641760
rect 127410 641640 127580 641760
rect 127710 641640 127880 641760
rect 128010 641640 128180 641760
rect 128310 641640 128480 641760
rect 128610 641640 128780 641760
rect 128910 641640 129080 641760
rect 129210 641640 129380 641760
rect 129510 641640 129680 641760
rect 129810 641640 129980 641760
rect 130110 641640 130280 641760
rect 130410 641640 130580 641760
rect 130710 641640 130880 641760
rect 131010 641640 131180 641760
rect 131310 641640 131470 641760
rect 131600 641640 131630 641760
rect 123830 641620 131630 641640
rect 123880 636810 129230 636820
rect 123880 636690 124020 636810
rect 124150 636690 124320 636810
rect 124450 636690 124620 636810
rect 124750 636690 124920 636810
rect 125050 636690 125220 636810
rect 125350 636690 125520 636810
rect 125650 636690 125820 636810
rect 125950 636690 126120 636810
rect 126250 636690 126420 636810
rect 126550 636690 126720 636810
rect 126850 636690 127020 636810
rect 127150 636690 127320 636810
rect 127450 636690 127620 636810
rect 127750 636690 127920 636810
rect 128050 636690 128220 636810
rect 128350 636690 128520 636810
rect 128650 636690 128820 636810
rect 128950 636700 129230 636810
rect 128950 636690 129100 636700
rect 123880 636680 129100 636690
rect 123880 636610 124010 636680
rect 123880 636360 124010 636490
rect 129100 636470 129230 636580
rect 123880 636100 124010 636240
rect 123880 635820 124010 635980
rect 123880 635660 124010 635700
rect 129100 635820 129230 635900
rect 129100 635660 129230 635700
rect 123880 635540 124020 635660
rect 124150 635540 124320 635660
rect 124450 635540 124620 635660
rect 124750 635540 124920 635660
rect 125050 635540 125220 635660
rect 125350 635540 125520 635660
rect 125650 635540 125820 635660
rect 125950 635540 126120 635660
rect 126250 635540 126420 635660
rect 126550 635540 126720 635660
rect 126850 635540 127020 635660
rect 127150 635540 127320 635660
rect 127450 635540 127620 635660
rect 127750 635540 127920 635660
rect 128050 635540 128220 635660
rect 128350 635540 128520 635660
rect 128650 635540 128820 635660
rect 128950 635540 129230 635660
rect 124160 630720 129300 630740
rect 124160 630600 124390 630720
rect 124520 630600 124690 630720
rect 124820 630600 124990 630720
rect 125120 630600 125290 630720
rect 125420 630600 125590 630720
rect 125720 630600 125890 630720
rect 126020 630600 126190 630720
rect 126320 630600 126490 630720
rect 126620 630600 126790 630720
rect 126920 630600 127090 630720
rect 127220 630600 127390 630720
rect 127520 630600 127690 630720
rect 127820 630600 127990 630720
rect 128120 630600 128290 630720
rect 128420 630600 128590 630720
rect 128720 630600 128890 630720
rect 129020 630620 129300 630720
rect 129020 630600 129170 630620
rect 124160 630590 129170 630600
rect 124160 630240 124290 630470
rect 129170 630410 129300 630500
rect 124160 629860 124290 630120
rect 124160 629690 124290 629740
rect 129170 629690 129300 629840
rect 124160 629680 129300 629690
rect 124160 629560 124390 629680
rect 124520 629560 124690 629680
rect 124820 629560 124990 629680
rect 125120 629560 125290 629680
rect 125420 629560 125590 629680
rect 125720 629560 125890 629680
rect 126020 629560 126190 629680
rect 126320 629560 126490 629680
rect 126620 629560 126790 629680
rect 126920 629560 127090 629680
rect 127220 629560 127390 629680
rect 127520 629560 127690 629680
rect 127820 629560 127990 629680
rect 128120 629560 128290 629680
rect 128420 629560 128590 629680
rect 128720 629560 128890 629680
rect 129020 629560 129300 629680
rect 124160 629540 129300 629560
rect 124410 624210 128950 624220
rect 124410 624140 124630 624210
rect 124540 624090 124630 624140
rect 124760 624090 124930 624210
rect 125060 624090 125230 624210
rect 125360 624090 125530 624210
rect 125660 624090 125830 624210
rect 125960 624090 126130 624210
rect 126260 624090 126430 624210
rect 126560 624090 126730 624210
rect 126860 624090 127030 624210
rect 127160 624090 127330 624210
rect 127460 624090 127630 624210
rect 127760 624090 127930 624210
rect 128060 624090 128230 624210
rect 128360 624090 128530 624210
rect 128660 624150 128950 624210
rect 128660 624090 128820 624150
rect 124540 624070 128820 624090
rect 124410 623840 124540 624020
rect 124410 623540 124540 623720
rect 128820 623890 128950 624030
rect 124410 623240 124540 623420
rect 128820 623170 128950 623320
rect 124540 623160 128950 623170
rect 124540 623120 124670 623160
rect 124410 623040 124670 623120
rect 124800 623040 124970 623160
rect 125100 623040 125270 623160
rect 125400 623040 125570 623160
rect 125700 623040 125870 623160
rect 126000 623040 126170 623160
rect 126300 623040 126470 623160
rect 126600 623040 126770 623160
rect 126900 623040 127070 623160
rect 127200 623040 127370 623160
rect 127500 623040 127670 623160
rect 127800 623040 127970 623160
rect 128100 623040 128270 623160
rect 128400 623040 128570 623160
rect 128700 623040 128950 623160
rect 124410 623020 128950 623040
rect 125040 618860 125230 618990
rect 125370 618860 125730 618990
rect 125870 618860 126230 618990
rect 126370 618860 126730 618990
rect 126870 618860 127230 618990
rect 127370 618860 127730 618990
rect 127870 618860 128230 618990
rect 128370 618860 128730 618990
rect 128870 618860 129230 618990
rect 129370 618860 129730 618990
rect 129870 618860 130230 618990
rect 130370 618860 130730 618990
rect 130870 618860 131230 618990
rect 131370 618860 131730 618990
rect 131870 618860 132080 618990
rect 125040 618770 125180 618860
rect 131940 618790 132080 618860
rect 125040 618410 125180 618640
rect 125040 618190 125180 618280
rect 131940 618420 132080 618660
rect 131940 618190 132080 618290
rect 125040 618060 125230 618190
rect 125370 618060 125730 618190
rect 125870 618060 126230 618190
rect 126370 618060 126730 618190
rect 126870 618060 127230 618190
rect 127370 618060 127730 618190
rect 127870 618060 128230 618190
rect 128370 618060 128730 618190
rect 128870 618060 129230 618190
rect 129370 618060 129730 618190
rect 129870 618060 130230 618190
rect 130370 618060 130730 618190
rect 130870 618060 131230 618190
rect 131370 618060 131730 618190
rect 131870 618060 132080 618190
rect 124690 611410 124880 611540
rect 125020 611410 125380 611540
rect 125520 611410 125880 611540
rect 126020 611410 126380 611540
rect 126520 611410 126880 611540
rect 127020 611410 127380 611540
rect 127520 611410 127880 611540
rect 128020 611410 128380 611540
rect 128520 611410 128880 611540
rect 129020 611410 129380 611540
rect 129520 611410 129880 611540
rect 130020 611410 130380 611540
rect 130520 611410 130880 611540
rect 131020 611410 131380 611540
rect 131520 611410 131730 611540
rect 124690 611320 124830 611410
rect 131590 611340 131730 611410
rect 124690 610960 124830 611190
rect 131590 610970 131730 611210
rect 124690 610740 124830 610830
rect 131590 610740 131730 610840
rect 124690 610610 124880 610740
rect 125020 610610 125380 610740
rect 125520 610610 125880 610740
rect 126020 610610 126380 610740
rect 126520 610610 126880 610740
rect 127020 610610 127380 610740
rect 127520 610610 127880 610740
rect 128020 610610 128380 610740
rect 128520 610610 128880 610740
rect 129020 610610 129380 610740
rect 129520 610610 129880 610740
rect 130020 610610 130380 610740
rect 130520 610610 130880 610740
rect 131020 610610 131380 610740
rect 131520 610610 131730 610740
rect 124820 605360 125010 605490
rect 125150 605360 125510 605490
rect 125650 605360 126010 605490
rect 126150 605360 126510 605490
rect 126650 605360 127010 605490
rect 127150 605360 127510 605490
rect 127650 605360 128010 605490
rect 128150 605360 128510 605490
rect 128650 605360 129010 605490
rect 129150 605360 129510 605490
rect 129650 605360 130010 605490
rect 130150 605360 130510 605490
rect 130650 605360 131010 605490
rect 131150 605360 131510 605490
rect 131650 605360 131860 605490
rect 124820 605270 124960 605360
rect 131720 605290 131860 605360
rect 124820 604810 124960 605140
rect 131720 604820 131860 605160
rect 124820 604590 124960 604680
rect 131720 604590 131860 604690
rect 124820 604460 125010 604590
rect 125150 604460 125510 604590
rect 125650 604460 126010 604590
rect 126150 604460 126510 604590
rect 126650 604460 127010 604590
rect 127150 604460 127510 604590
rect 127650 604460 128010 604590
rect 128150 604460 128510 604590
rect 128650 604460 129010 604590
rect 129150 604460 129510 604590
rect 129650 604460 130010 604590
rect 130150 604460 130510 604590
rect 130650 604460 131010 604590
rect 131150 604460 131510 604590
rect 131650 604460 131860 604590
rect 124620 599100 124810 599230
rect 124950 599100 125310 599230
rect 125450 599100 125810 599230
rect 125950 599100 126310 599230
rect 126450 599100 126810 599230
rect 126950 599100 127310 599230
rect 127450 599100 127810 599230
rect 127950 599100 128310 599230
rect 128450 599100 128810 599230
rect 128950 599100 129310 599230
rect 129450 599100 129810 599230
rect 129950 599100 130310 599230
rect 130450 599100 130810 599230
rect 130950 599100 131310 599230
rect 131450 599100 131660 599230
rect 124620 599010 124760 599100
rect 131520 599030 131660 599100
rect 124620 598450 124760 598880
rect 131520 598460 131660 598900
rect 124620 598230 124760 598320
rect 131520 598230 131660 598330
rect 124620 598100 124810 598230
rect 124950 598100 125310 598230
rect 125450 598100 125810 598230
rect 125950 598100 126310 598230
rect 126450 598100 126810 598230
rect 126950 598100 127310 598230
rect 127450 598100 127810 598230
rect 127950 598100 128310 598230
rect 128450 598100 128810 598230
rect 128950 598100 129310 598230
rect 129450 598100 129810 598230
rect 129950 598100 130310 598230
rect 130450 598100 130810 598230
rect 130950 598100 131310 598230
rect 131450 598100 131660 598230
rect 119510 592750 119620 592770
rect 119510 592590 119540 592750
rect 119580 592590 119620 592750
rect 119510 592570 119620 592590
rect 120170 592750 120280 592770
rect 120170 592590 120210 592750
rect 120250 592590 120280 592750
rect 120170 592570 120280 592590
rect 124580 591550 124770 591680
rect 124910 591550 125270 591680
rect 125410 591550 125770 591680
rect 125910 591550 126270 591680
rect 126410 591550 126770 591680
rect 126910 591550 127270 591680
rect 127410 591550 127770 591680
rect 127910 591550 128270 591680
rect 128410 591550 128770 591680
rect 128910 591550 129270 591680
rect 129410 591550 129770 591680
rect 129910 591550 130270 591680
rect 130410 591550 130770 591680
rect 130910 591550 131270 591680
rect 131410 591550 131620 591680
rect 124580 591460 124720 591550
rect 131480 591480 131620 591550
rect 124580 590800 124720 591330
rect 131480 590810 131620 591350
rect 124580 590580 124720 590670
rect 131480 590580 131620 590680
rect 124580 590450 124770 590580
rect 124910 590450 125270 590580
rect 125410 590450 125770 590580
rect 125910 590450 126270 590580
rect 126410 590450 126770 590580
rect 126910 590450 127270 590580
rect 127410 590450 127770 590580
rect 127910 590450 128270 590580
rect 128410 590450 128770 590580
rect 128910 590450 129270 590580
rect 129410 590450 129770 590580
rect 129910 590450 130270 590580
rect 130410 590450 130770 590580
rect 130910 590450 131270 590580
rect 131410 590450 131620 590580
rect 119550 583210 119660 583230
rect 119550 583050 119580 583210
rect 119620 583050 119660 583210
rect 119550 583030 119660 583050
rect 120210 583210 120320 583230
rect 120210 583050 120250 583210
rect 120290 583050 120320 583210
rect 120210 583030 120320 583050
rect 125040 582570 125230 582700
rect 125370 582570 125780 582700
rect 125920 582570 126330 582700
rect 126520 582570 126930 582700
rect 127070 582570 127480 582700
rect 127670 582570 128080 582700
rect 128220 582570 128630 582700
rect 128820 582570 129230 582700
rect 129370 582570 129780 582700
rect 129970 582570 130380 582700
rect 130520 582570 130930 582700
rect 131120 582570 131530 582700
rect 131670 582570 132080 582700
rect 132270 582570 132680 582700
rect 132820 582570 133030 582700
rect 125040 582480 125180 582570
rect 132890 582500 133030 582570
rect 125040 582120 125180 582350
rect 125040 581900 125180 581990
rect 132890 582130 133030 582370
rect 132890 581900 133030 582000
rect 125040 581770 125230 581900
rect 125370 581770 125780 581900
rect 125920 581770 126330 581900
rect 126520 581770 126930 581900
rect 127070 581770 127480 581900
rect 127670 581770 128080 581900
rect 128220 581770 128630 581900
rect 128820 581770 129230 581900
rect 129370 581770 129780 581900
rect 129970 581770 130380 581900
rect 130520 581770 130930 581900
rect 131120 581770 131530 581900
rect 131670 581770 132080 581900
rect 132270 581770 132680 581900
rect 132820 581770 133030 581900
rect 119590 574190 119700 574210
rect 119590 574030 119620 574190
rect 119660 574030 119700 574190
rect 119590 574010 119700 574030
rect 120250 574190 120360 574210
rect 120250 574030 120290 574190
rect 120330 574030 120360 574190
rect 120250 574010 120360 574030
rect 125080 573550 125270 573680
rect 125410 573550 125820 573680
rect 125960 573550 126370 573680
rect 126560 573550 126970 573680
rect 127110 573550 127520 573680
rect 127710 573550 128120 573680
rect 128260 573550 128670 573680
rect 128860 573550 129270 573680
rect 129410 573550 129820 573680
rect 130010 573550 130420 573680
rect 130560 573550 130970 573680
rect 131160 573550 131570 573680
rect 131710 573550 132120 573680
rect 132310 573550 132720 573680
rect 132860 573550 133070 573680
rect 125080 573460 125220 573550
rect 132930 573480 133070 573550
rect 125080 573000 125220 573330
rect 125080 572780 125220 572870
rect 132930 573010 133070 573350
rect 132930 572780 133070 572880
rect 125080 572650 125270 572780
rect 125410 572650 125820 572780
rect 125960 572650 126370 572780
rect 126560 572650 126970 572780
rect 127110 572650 127520 572780
rect 127710 572650 128120 572780
rect 128260 572650 128670 572780
rect 128860 572650 129270 572780
rect 129410 572650 129820 572780
rect 130010 572650 130420 572780
rect 130560 572650 130970 572780
rect 131160 572650 131570 572780
rect 131710 572650 132120 572780
rect 132310 572650 132720 572780
rect 132860 572650 133070 572780
rect 119540 566520 119650 566540
rect 119540 566360 119570 566520
rect 119610 566360 119650 566520
rect 119540 566340 119650 566360
rect 120200 566520 120310 566540
rect 120200 566360 120240 566520
rect 120280 566360 120310 566520
rect 120200 566340 120310 566360
rect 125030 565880 125220 566010
rect 125360 565880 125770 566010
rect 125910 565880 126320 566010
rect 126510 565880 126920 566010
rect 127060 565880 127470 566010
rect 127660 565880 128070 566010
rect 128210 565880 128620 566010
rect 128810 565880 129220 566010
rect 129360 565880 129770 566010
rect 129960 565880 130370 566010
rect 130510 565880 130920 566010
rect 131110 565880 131520 566010
rect 131660 565880 132070 566010
rect 132260 565880 132670 566010
rect 132810 565880 133020 566010
rect 125030 565790 125170 565880
rect 132880 565810 133020 565880
rect 125030 565230 125170 565660
rect 125030 565010 125170 565100
rect 132880 565240 133020 565680
rect 132880 565010 133020 565110
rect 125030 564880 125220 565010
rect 125360 564880 125770 565010
rect 125910 564880 126320 565010
rect 126510 564880 126920 565010
rect 127060 564880 127470 565010
rect 127660 564880 128070 565010
rect 128210 564880 128620 565010
rect 128810 564880 129220 565010
rect 129360 564880 129770 565010
rect 129960 564880 130370 565010
rect 130510 564880 130920 565010
rect 131110 564880 131520 565010
rect 131660 564880 132070 565010
rect 132260 564880 132670 565010
rect 132810 564880 133020 565010
rect 119540 559980 119650 560000
rect 119540 559820 119570 559980
rect 119610 559820 119650 559980
rect 119540 559800 119650 559820
rect 120200 559980 120310 560000
rect 120200 559820 120240 559980
rect 120280 559820 120310 559980
rect 120200 559800 120310 559820
rect 125030 559340 125220 559470
rect 125360 559340 125770 559470
rect 125910 559340 126320 559470
rect 126510 559340 126920 559470
rect 127060 559340 127470 559470
rect 127660 559340 128070 559470
rect 128210 559340 128620 559470
rect 128810 559340 129220 559470
rect 129360 559340 129770 559470
rect 129960 559340 130370 559470
rect 130510 559340 130920 559470
rect 131110 559340 131520 559470
rect 131660 559340 132070 559470
rect 132260 559340 132670 559470
rect 132810 559340 133020 559470
rect 125030 559250 125170 559340
rect 132880 559270 133020 559340
rect 125030 558590 125170 559120
rect 125030 558370 125170 558460
rect 132880 558600 133020 559140
rect 132880 558370 133020 558470
rect 125030 558240 125220 558370
rect 125360 558240 125770 558370
rect 125910 558240 126320 558370
rect 126510 558240 126920 558370
rect 127060 558240 127470 558370
rect 127660 558240 128070 558370
rect 128210 558240 128620 558370
rect 128810 558240 129220 558370
rect 129360 558240 129770 558370
rect 129960 558240 130370 558370
rect 130510 558240 130920 558370
rect 131110 558240 131520 558370
rect 131660 558240 132070 558370
rect 132260 558240 132670 558370
rect 132810 558240 133020 558370
rect 119610 553150 119720 553170
rect 119610 552990 119640 553150
rect 119680 552990 119720 553150
rect 119610 552970 119720 552990
rect 120270 553150 120380 553170
rect 120270 552990 120310 553150
rect 120350 552990 120380 553150
rect 120270 552970 120380 552990
rect 125100 552510 125290 552640
rect 125430 552510 125890 552640
rect 126030 552510 126490 552640
rect 126730 552510 127190 552640
rect 127330 552510 127790 552640
rect 128030 552510 128490 552640
rect 128630 552510 129090 552640
rect 129330 552510 129790 552640
rect 129930 552510 130390 552640
rect 130630 552510 131090 552640
rect 131230 552510 131690 552640
rect 131930 552510 132390 552640
rect 132530 552510 132990 552640
rect 133230 552510 133690 552640
rect 133830 552510 134040 552640
rect 125100 552420 125240 552510
rect 133900 552440 134040 552510
rect 125100 552060 125240 552290
rect 125100 551840 125240 551930
rect 133900 552070 134040 552310
rect 133900 551840 134040 551940
rect 125100 551710 125290 551840
rect 125430 551710 125890 551840
rect 126030 551710 126490 551840
rect 126730 551710 127190 551840
rect 127330 551710 127790 551840
rect 128030 551710 128490 551840
rect 128630 551710 129090 551840
rect 129330 551710 129790 551840
rect 129930 551710 130390 551840
rect 130630 551710 131090 551840
rect 131230 551710 131690 551840
rect 131930 551710 132390 551840
rect 132530 551710 132990 551840
rect 133230 551710 133690 551840
rect 133830 551710 134040 551840
rect 119610 545580 119720 545600
rect 119610 545420 119640 545580
rect 119680 545420 119720 545580
rect 119610 545400 119720 545420
rect 120270 545580 120380 545600
rect 120270 545420 120310 545580
rect 120350 545420 120380 545580
rect 120270 545400 120380 545420
rect 125100 544940 125290 545070
rect 125430 544940 125890 545070
rect 126030 544940 126490 545070
rect 126730 544940 127190 545070
rect 127330 544940 127790 545070
rect 128030 544940 128490 545070
rect 128630 544940 129090 545070
rect 129330 544940 129790 545070
rect 129930 544940 130390 545070
rect 130630 544940 131090 545070
rect 131230 544940 131690 545070
rect 131930 544940 132390 545070
rect 132530 544940 132990 545070
rect 133230 544940 133690 545070
rect 133830 544940 134040 545070
rect 125100 544850 125240 544940
rect 133900 544870 134040 544940
rect 125100 544290 125240 544720
rect 125100 544070 125240 544160
rect 133900 544300 134040 544740
rect 133900 544070 134040 544170
rect 125100 543940 125290 544070
rect 125430 543940 125890 544070
rect 126030 543940 126490 544070
rect 126730 543940 127190 544070
rect 127330 543940 127790 544070
rect 128030 543940 128490 544070
rect 128630 543940 129090 544070
rect 129330 543940 129790 544070
rect 129930 543940 130390 544070
rect 130630 543940 131090 544070
rect 131230 543940 131690 544070
rect 131930 543940 132390 544070
rect 132530 543940 132990 544070
rect 133230 543940 133690 544070
rect 133830 543940 134040 544070
rect 119580 537520 119690 537540
rect 119580 537360 119610 537520
rect 119650 537360 119690 537520
rect 119580 537340 119690 537360
rect 120240 537520 120350 537540
rect 120240 537360 120280 537520
rect 120320 537360 120350 537520
rect 120240 537340 120350 537360
rect 125070 536880 125260 537010
rect 125400 536880 125860 537010
rect 126000 536880 126460 537010
rect 126700 536880 127160 537010
rect 127300 536880 127760 537010
rect 128000 536880 128460 537010
rect 128600 536880 129060 537010
rect 129300 536880 129760 537010
rect 129900 536880 130360 537010
rect 130600 536880 131060 537010
rect 131200 536880 131660 537010
rect 131900 536880 132360 537010
rect 132500 536880 132960 537010
rect 133200 536880 133660 537010
rect 133800 536880 134010 537010
rect 125070 536790 125210 536880
rect 133870 536810 134010 536880
rect 125070 536030 125210 536660
rect 125070 535810 125210 535900
rect 133870 536040 134010 536680
rect 133870 535810 134010 535910
rect 125070 535680 125260 535810
rect 125400 535680 125860 535810
rect 126000 535680 126460 535810
rect 126700 535680 127160 535810
rect 127300 535680 127760 535810
rect 128000 535680 128460 535810
rect 128600 535680 129060 535810
rect 129300 535680 129760 535810
rect 129900 535680 130360 535810
rect 130600 535680 131060 535810
rect 131200 535680 131660 535810
rect 131900 535680 132360 535810
rect 132500 535680 132960 535810
rect 133200 535680 133660 535810
rect 133800 535680 134010 535810
<< nsubdiff >>
rect 119510 593260 119620 593280
rect 119510 593100 119540 593260
rect 119580 593100 119620 593260
rect 119510 593080 119620 593100
rect 120170 593260 120280 593280
rect 120170 593100 120210 593260
rect 120250 593100 120280 593260
rect 120170 593080 120280 593100
rect 119550 583720 119660 583740
rect 119550 583560 119580 583720
rect 119620 583560 119660 583720
rect 119550 583540 119660 583560
rect 120210 583720 120320 583740
rect 120210 583560 120250 583720
rect 120290 583560 120320 583720
rect 120210 583540 120320 583560
rect 119590 574700 119700 574720
rect 119590 574540 119620 574700
rect 119660 574540 119700 574700
rect 119590 574520 119700 574540
rect 120250 574700 120360 574720
rect 120250 574540 120290 574700
rect 120330 574540 120360 574700
rect 120250 574520 120360 574540
rect 119540 567030 119650 567050
rect 119540 566870 119570 567030
rect 119610 566870 119650 567030
rect 119540 566850 119650 566870
rect 120200 567030 120310 567050
rect 120200 566870 120240 567030
rect 120280 566870 120310 567030
rect 120200 566850 120310 566870
rect 119540 560490 119650 560510
rect 119540 560330 119570 560490
rect 119610 560330 119650 560490
rect 119540 560310 119650 560330
rect 120200 560490 120310 560510
rect 120200 560330 120240 560490
rect 120280 560330 120310 560490
rect 120200 560310 120310 560330
rect 119610 553660 119720 553680
rect 119610 553500 119640 553660
rect 119680 553500 119720 553660
rect 119610 553480 119720 553500
rect 120270 553660 120380 553680
rect 120270 553500 120310 553660
rect 120350 553500 120380 553660
rect 120270 553480 120380 553500
rect 119610 546090 119720 546110
rect 119610 545930 119640 546090
rect 119680 545930 119720 546090
rect 119610 545910 119720 545930
rect 120270 546090 120380 546110
rect 120270 545930 120310 546090
rect 120350 545930 120380 546090
rect 120270 545910 120380 545930
rect 119580 538030 119690 538050
rect 119580 537870 119610 538030
rect 119650 537870 119690 538030
rect 119580 537850 119690 537870
rect 120240 538030 120350 538050
rect 120240 537870 120280 538030
rect 120320 537870 120350 538030
rect 120240 537850 120350 537870
<< psubdiffcont >>
rect 123870 642900 124000 643020
rect 124110 642900 124240 643020
rect 124410 642900 124540 643020
rect 124710 642900 124840 643020
rect 125010 642900 125140 643020
rect 125310 642900 125440 643020
rect 125610 642900 125740 643020
rect 125910 642900 126040 643020
rect 126210 642900 126340 643020
rect 126510 642900 126640 643020
rect 126810 642900 126940 643020
rect 127110 642900 127240 643020
rect 127410 642900 127540 643020
rect 127710 642900 127840 643020
rect 128010 642900 128140 643020
rect 128310 642900 128440 643020
rect 128610 642900 128740 643020
rect 128910 642900 129040 643020
rect 129210 642900 129340 643020
rect 129510 642900 129640 643020
rect 129810 642900 129940 643020
rect 130110 642900 130240 643020
rect 130410 642900 130540 643020
rect 130710 642900 130840 643020
rect 131010 642900 131140 643020
rect 131310 642900 131440 643020
rect 123830 642700 123960 642820
rect 123830 642040 123960 642610
rect 131500 642690 131630 642810
rect 123830 641810 123960 641930
rect 131500 642060 131630 642630
rect 123980 641640 124110 641760
rect 124280 641640 124410 641760
rect 124580 641640 124710 641760
rect 124880 641640 125010 641760
rect 125180 641640 125310 641760
rect 125480 641640 125610 641760
rect 125780 641640 125910 641760
rect 126080 641640 126210 641760
rect 126380 641640 126510 641760
rect 126680 641640 126810 641760
rect 126980 641640 127110 641760
rect 127280 641640 127410 641760
rect 127580 641640 127710 641760
rect 127880 641640 128010 641760
rect 128180 641640 128310 641760
rect 128480 641640 128610 641760
rect 128780 641640 128910 641760
rect 129080 641640 129210 641760
rect 129380 641640 129510 641760
rect 129680 641640 129810 641760
rect 129980 641640 130110 641760
rect 130280 641640 130410 641760
rect 130580 641640 130710 641760
rect 130880 641640 131010 641760
rect 131180 641640 131310 641760
rect 131470 641640 131600 641760
rect 124020 636690 124150 636810
rect 124320 636690 124450 636810
rect 124620 636690 124750 636810
rect 124920 636690 125050 636810
rect 125220 636690 125350 636810
rect 125520 636690 125650 636810
rect 125820 636690 125950 636810
rect 126120 636690 126250 636810
rect 126420 636690 126550 636810
rect 126720 636690 126850 636810
rect 127020 636690 127150 636810
rect 127320 636690 127450 636810
rect 127620 636690 127750 636810
rect 127920 636690 128050 636810
rect 128220 636690 128350 636810
rect 128520 636690 128650 636810
rect 128820 636690 128950 636810
rect 123880 636490 124010 636610
rect 123880 636240 124010 636360
rect 129100 636580 129230 636700
rect 123880 635980 124010 636100
rect 123880 635700 124010 635820
rect 129100 635900 129230 636470
rect 129100 635700 129230 635820
rect 124020 635540 124150 635660
rect 124320 635540 124450 635660
rect 124620 635540 124750 635660
rect 124920 635540 125050 635660
rect 125220 635540 125350 635660
rect 125520 635540 125650 635660
rect 125820 635540 125950 635660
rect 126120 635540 126250 635660
rect 126420 635540 126550 635660
rect 126720 635540 126850 635660
rect 127020 635540 127150 635660
rect 127320 635540 127450 635660
rect 127620 635540 127750 635660
rect 127920 635540 128050 635660
rect 128220 635540 128350 635660
rect 128520 635540 128650 635660
rect 128820 635540 128950 635660
rect 124390 630600 124520 630720
rect 124690 630600 124820 630720
rect 124990 630600 125120 630720
rect 125290 630600 125420 630720
rect 125590 630600 125720 630720
rect 125890 630600 126020 630720
rect 126190 630600 126320 630720
rect 126490 630600 126620 630720
rect 126790 630600 126920 630720
rect 127090 630600 127220 630720
rect 127390 630600 127520 630720
rect 127690 630600 127820 630720
rect 127990 630600 128120 630720
rect 128290 630600 128420 630720
rect 128590 630600 128720 630720
rect 128890 630600 129020 630720
rect 124160 630470 124290 630590
rect 124160 630120 124290 630240
rect 129170 630500 129300 630620
rect 124160 629740 124290 629860
rect 129170 629840 129300 630410
rect 124390 629560 124520 629680
rect 124690 629560 124820 629680
rect 124990 629560 125120 629680
rect 125290 629560 125420 629680
rect 125590 629560 125720 629680
rect 125890 629560 126020 629680
rect 126190 629560 126320 629680
rect 126490 629560 126620 629680
rect 126790 629560 126920 629680
rect 127090 629560 127220 629680
rect 127390 629560 127520 629680
rect 127690 629560 127820 629680
rect 127990 629560 128120 629680
rect 128290 629560 128420 629680
rect 128590 629560 128720 629680
rect 128890 629560 129020 629680
rect 124410 624020 124540 624140
rect 124630 624090 124760 624210
rect 124930 624090 125060 624210
rect 125230 624090 125360 624210
rect 125530 624090 125660 624210
rect 125830 624090 125960 624210
rect 126130 624090 126260 624210
rect 126430 624090 126560 624210
rect 126730 624090 126860 624210
rect 127030 624090 127160 624210
rect 127330 624090 127460 624210
rect 127630 624090 127760 624210
rect 127930 624090 128060 624210
rect 128230 624090 128360 624210
rect 128530 624090 128660 624210
rect 128820 624030 128950 624150
rect 124410 623720 124540 623840
rect 124410 623420 124540 623540
rect 124410 623120 124540 623240
rect 128820 623320 128950 623890
rect 124670 623040 124800 623160
rect 124970 623040 125100 623160
rect 125270 623040 125400 623160
rect 125570 623040 125700 623160
rect 125870 623040 126000 623160
rect 126170 623040 126300 623160
rect 126470 623040 126600 623160
rect 126770 623040 126900 623160
rect 127070 623040 127200 623160
rect 127370 623040 127500 623160
rect 127670 623040 127800 623160
rect 127970 623040 128100 623160
rect 128270 623040 128400 623160
rect 128570 623040 128700 623160
rect 125230 618860 125370 618990
rect 125730 618860 125870 618990
rect 126230 618860 126370 618990
rect 126730 618860 126870 618990
rect 127230 618860 127370 618990
rect 127730 618860 127870 618990
rect 128230 618860 128370 618990
rect 128730 618860 128870 618990
rect 129230 618860 129370 618990
rect 129730 618860 129870 618990
rect 130230 618860 130370 618990
rect 130730 618860 130870 618990
rect 131230 618860 131370 618990
rect 131730 618860 131870 618990
rect 125040 618640 125180 618770
rect 131940 618660 132080 618790
rect 125040 618280 125180 618410
rect 131940 618290 132080 618420
rect 125230 618060 125370 618190
rect 125730 618060 125870 618190
rect 126230 618060 126370 618190
rect 126730 618060 126870 618190
rect 127230 618060 127370 618190
rect 127730 618060 127870 618190
rect 128230 618060 128370 618190
rect 128730 618060 128870 618190
rect 129230 618060 129370 618190
rect 129730 618060 129870 618190
rect 130230 618060 130370 618190
rect 130730 618060 130870 618190
rect 131230 618060 131370 618190
rect 131730 618060 131870 618190
rect 124880 611410 125020 611540
rect 125380 611410 125520 611540
rect 125880 611410 126020 611540
rect 126380 611410 126520 611540
rect 126880 611410 127020 611540
rect 127380 611410 127520 611540
rect 127880 611410 128020 611540
rect 128380 611410 128520 611540
rect 128880 611410 129020 611540
rect 129380 611410 129520 611540
rect 129880 611410 130020 611540
rect 130380 611410 130520 611540
rect 130880 611410 131020 611540
rect 131380 611410 131520 611540
rect 124690 611190 124830 611320
rect 124690 610830 124830 610960
rect 131590 611210 131730 611340
rect 131590 610840 131730 610970
rect 124880 610610 125020 610740
rect 125380 610610 125520 610740
rect 125880 610610 126020 610740
rect 126380 610610 126520 610740
rect 126880 610610 127020 610740
rect 127380 610610 127520 610740
rect 127880 610610 128020 610740
rect 128380 610610 128520 610740
rect 128880 610610 129020 610740
rect 129380 610610 129520 610740
rect 129880 610610 130020 610740
rect 130380 610610 130520 610740
rect 130880 610610 131020 610740
rect 131380 610610 131520 610740
rect 125010 605360 125150 605490
rect 125510 605360 125650 605490
rect 126010 605360 126150 605490
rect 126510 605360 126650 605490
rect 127010 605360 127150 605490
rect 127510 605360 127650 605490
rect 128010 605360 128150 605490
rect 128510 605360 128650 605490
rect 129010 605360 129150 605490
rect 129510 605360 129650 605490
rect 130010 605360 130150 605490
rect 130510 605360 130650 605490
rect 131010 605360 131150 605490
rect 131510 605360 131650 605490
rect 124820 605140 124960 605270
rect 124820 604680 124960 604810
rect 131720 605160 131860 605290
rect 131720 604690 131860 604820
rect 125010 604460 125150 604590
rect 125510 604460 125650 604590
rect 126010 604460 126150 604590
rect 126510 604460 126650 604590
rect 127010 604460 127150 604590
rect 127510 604460 127650 604590
rect 128010 604460 128150 604590
rect 128510 604460 128650 604590
rect 129010 604460 129150 604590
rect 129510 604460 129650 604590
rect 130010 604460 130150 604590
rect 130510 604460 130650 604590
rect 131010 604460 131150 604590
rect 131510 604460 131650 604590
rect 124810 599100 124950 599230
rect 125310 599100 125450 599230
rect 125810 599100 125950 599230
rect 126310 599100 126450 599230
rect 126810 599100 126950 599230
rect 127310 599100 127450 599230
rect 127810 599100 127950 599230
rect 128310 599100 128450 599230
rect 128810 599100 128950 599230
rect 129310 599100 129450 599230
rect 129810 599100 129950 599230
rect 130310 599100 130450 599230
rect 130810 599100 130950 599230
rect 131310 599100 131450 599230
rect 124620 598880 124760 599010
rect 124620 598320 124760 598450
rect 131520 598900 131660 599030
rect 131520 598330 131660 598460
rect 124810 598100 124950 598230
rect 125310 598100 125450 598230
rect 125810 598100 125950 598230
rect 126310 598100 126450 598230
rect 126810 598100 126950 598230
rect 127310 598100 127450 598230
rect 127810 598100 127950 598230
rect 128310 598100 128450 598230
rect 128810 598100 128950 598230
rect 129310 598100 129450 598230
rect 129810 598100 129950 598230
rect 130310 598100 130450 598230
rect 130810 598100 130950 598230
rect 131310 598100 131450 598230
rect 119540 592590 119580 592750
rect 120210 592590 120250 592750
rect 124770 591550 124910 591680
rect 125270 591550 125410 591680
rect 125770 591550 125910 591680
rect 126270 591550 126410 591680
rect 126770 591550 126910 591680
rect 127270 591550 127410 591680
rect 127770 591550 127910 591680
rect 128270 591550 128410 591680
rect 128770 591550 128910 591680
rect 129270 591550 129410 591680
rect 129770 591550 129910 591680
rect 130270 591550 130410 591680
rect 130770 591550 130910 591680
rect 131270 591550 131410 591680
rect 124580 591330 124720 591460
rect 124580 590670 124720 590800
rect 131480 591350 131620 591480
rect 131480 590680 131620 590810
rect 124770 590450 124910 590580
rect 125270 590450 125410 590580
rect 125770 590450 125910 590580
rect 126270 590450 126410 590580
rect 126770 590450 126910 590580
rect 127270 590450 127410 590580
rect 127770 590450 127910 590580
rect 128270 590450 128410 590580
rect 128770 590450 128910 590580
rect 129270 590450 129410 590580
rect 129770 590450 129910 590580
rect 130270 590450 130410 590580
rect 130770 590450 130910 590580
rect 131270 590450 131410 590580
rect 119580 583050 119620 583210
rect 120250 583050 120290 583210
rect 125230 582570 125370 582700
rect 125780 582570 125920 582700
rect 126330 582570 126520 582700
rect 126930 582570 127070 582700
rect 127480 582570 127670 582700
rect 128080 582570 128220 582700
rect 128630 582570 128820 582700
rect 129230 582570 129370 582700
rect 129780 582570 129970 582700
rect 130380 582570 130520 582700
rect 130930 582570 131120 582700
rect 131530 582570 131670 582700
rect 132080 582570 132270 582700
rect 132680 582570 132820 582700
rect 125040 582350 125180 582480
rect 132890 582370 133030 582500
rect 125040 581990 125180 582120
rect 132890 582000 133030 582130
rect 125230 581770 125370 581900
rect 125780 581770 125920 581900
rect 126330 581770 126520 581900
rect 126930 581770 127070 581900
rect 127480 581770 127670 581900
rect 128080 581770 128220 581900
rect 128630 581770 128820 581900
rect 129230 581770 129370 581900
rect 129780 581770 129970 581900
rect 130380 581770 130520 581900
rect 130930 581770 131120 581900
rect 131530 581770 131670 581900
rect 132080 581770 132270 581900
rect 132680 581770 132820 581900
rect 119620 574030 119660 574190
rect 120290 574030 120330 574190
rect 125270 573550 125410 573680
rect 125820 573550 125960 573680
rect 126370 573550 126560 573680
rect 126970 573550 127110 573680
rect 127520 573550 127710 573680
rect 128120 573550 128260 573680
rect 128670 573550 128860 573680
rect 129270 573550 129410 573680
rect 129820 573550 130010 573680
rect 130420 573550 130560 573680
rect 130970 573550 131160 573680
rect 131570 573550 131710 573680
rect 132120 573550 132310 573680
rect 132720 573550 132860 573680
rect 125080 573330 125220 573460
rect 132930 573350 133070 573480
rect 125080 572870 125220 573000
rect 132930 572880 133070 573010
rect 125270 572650 125410 572780
rect 125820 572650 125960 572780
rect 126370 572650 126560 572780
rect 126970 572650 127110 572780
rect 127520 572650 127710 572780
rect 128120 572650 128260 572780
rect 128670 572650 128860 572780
rect 129270 572650 129410 572780
rect 129820 572650 130010 572780
rect 130420 572650 130560 572780
rect 130970 572650 131160 572780
rect 131570 572650 131710 572780
rect 132120 572650 132310 572780
rect 132720 572650 132860 572780
rect 119570 566360 119610 566520
rect 120240 566360 120280 566520
rect 125220 565880 125360 566010
rect 125770 565880 125910 566010
rect 126320 565880 126510 566010
rect 126920 565880 127060 566010
rect 127470 565880 127660 566010
rect 128070 565880 128210 566010
rect 128620 565880 128810 566010
rect 129220 565880 129360 566010
rect 129770 565880 129960 566010
rect 130370 565880 130510 566010
rect 130920 565880 131110 566010
rect 131520 565880 131660 566010
rect 132070 565880 132260 566010
rect 132670 565880 132810 566010
rect 125030 565660 125170 565790
rect 132880 565680 133020 565810
rect 125030 565100 125170 565230
rect 132880 565110 133020 565240
rect 125220 564880 125360 565010
rect 125770 564880 125910 565010
rect 126320 564880 126510 565010
rect 126920 564880 127060 565010
rect 127470 564880 127660 565010
rect 128070 564880 128210 565010
rect 128620 564880 128810 565010
rect 129220 564880 129360 565010
rect 129770 564880 129960 565010
rect 130370 564880 130510 565010
rect 130920 564880 131110 565010
rect 131520 564880 131660 565010
rect 132070 564880 132260 565010
rect 132670 564880 132810 565010
rect 119570 559820 119610 559980
rect 120240 559820 120280 559980
rect 125220 559340 125360 559470
rect 125770 559340 125910 559470
rect 126320 559340 126510 559470
rect 126920 559340 127060 559470
rect 127470 559340 127660 559470
rect 128070 559340 128210 559470
rect 128620 559340 128810 559470
rect 129220 559340 129360 559470
rect 129770 559340 129960 559470
rect 130370 559340 130510 559470
rect 130920 559340 131110 559470
rect 131520 559340 131660 559470
rect 132070 559340 132260 559470
rect 132670 559340 132810 559470
rect 125030 559120 125170 559250
rect 132880 559140 133020 559270
rect 125030 558460 125170 558590
rect 132880 558470 133020 558600
rect 125220 558240 125360 558370
rect 125770 558240 125910 558370
rect 126320 558240 126510 558370
rect 126920 558240 127060 558370
rect 127470 558240 127660 558370
rect 128070 558240 128210 558370
rect 128620 558240 128810 558370
rect 129220 558240 129360 558370
rect 129770 558240 129960 558370
rect 130370 558240 130510 558370
rect 130920 558240 131110 558370
rect 131520 558240 131660 558370
rect 132070 558240 132260 558370
rect 132670 558240 132810 558370
rect 119640 552990 119680 553150
rect 120310 552990 120350 553150
rect 125290 552510 125430 552640
rect 125890 552510 126030 552640
rect 126490 552510 126730 552640
rect 127190 552510 127330 552640
rect 127790 552510 128030 552640
rect 128490 552510 128630 552640
rect 129090 552510 129330 552640
rect 129790 552510 129930 552640
rect 130390 552510 130630 552640
rect 131090 552510 131230 552640
rect 131690 552510 131930 552640
rect 132390 552510 132530 552640
rect 132990 552510 133230 552640
rect 133690 552510 133830 552640
rect 125100 552290 125240 552420
rect 133900 552310 134040 552440
rect 125100 551930 125240 552060
rect 133900 551940 134040 552070
rect 125290 551710 125430 551840
rect 125890 551710 126030 551840
rect 126490 551710 126730 551840
rect 127190 551710 127330 551840
rect 127790 551710 128030 551840
rect 128490 551710 128630 551840
rect 129090 551710 129330 551840
rect 129790 551710 129930 551840
rect 130390 551710 130630 551840
rect 131090 551710 131230 551840
rect 131690 551710 131930 551840
rect 132390 551710 132530 551840
rect 132990 551710 133230 551840
rect 133690 551710 133830 551840
rect 119640 545420 119680 545580
rect 120310 545420 120350 545580
rect 125290 544940 125430 545070
rect 125890 544940 126030 545070
rect 126490 544940 126730 545070
rect 127190 544940 127330 545070
rect 127790 544940 128030 545070
rect 128490 544940 128630 545070
rect 129090 544940 129330 545070
rect 129790 544940 129930 545070
rect 130390 544940 130630 545070
rect 131090 544940 131230 545070
rect 131690 544940 131930 545070
rect 132390 544940 132530 545070
rect 132990 544940 133230 545070
rect 133690 544940 133830 545070
rect 125100 544720 125240 544850
rect 133900 544740 134040 544870
rect 125100 544160 125240 544290
rect 133900 544170 134040 544300
rect 125290 543940 125430 544070
rect 125890 543940 126030 544070
rect 126490 543940 126730 544070
rect 127190 543940 127330 544070
rect 127790 543940 128030 544070
rect 128490 543940 128630 544070
rect 129090 543940 129330 544070
rect 129790 543940 129930 544070
rect 130390 543940 130630 544070
rect 131090 543940 131230 544070
rect 131690 543940 131930 544070
rect 132390 543940 132530 544070
rect 132990 543940 133230 544070
rect 133690 543940 133830 544070
rect 119610 537360 119650 537520
rect 120280 537360 120320 537520
rect 125260 536880 125400 537010
rect 125860 536880 126000 537010
rect 126460 536880 126700 537010
rect 127160 536880 127300 537010
rect 127760 536880 128000 537010
rect 128460 536880 128600 537010
rect 129060 536880 129300 537010
rect 129760 536880 129900 537010
rect 130360 536880 130600 537010
rect 131060 536880 131200 537010
rect 131660 536880 131900 537010
rect 132360 536880 132500 537010
rect 132960 536880 133200 537010
rect 133660 536880 133800 537010
rect 125070 536660 125210 536790
rect 133870 536680 134010 536810
rect 125070 535900 125210 536030
rect 133870 535910 134010 536040
rect 125260 535680 125400 535810
rect 125860 535680 126000 535810
rect 126460 535680 126700 535810
rect 127160 535680 127300 535810
rect 127760 535680 128000 535810
rect 128460 535680 128600 535810
rect 129060 535680 129300 535810
rect 129760 535680 129900 535810
rect 130360 535680 130600 535810
rect 131060 535680 131200 535810
rect 131660 535680 131900 535810
rect 132360 535680 132500 535810
rect 132960 535680 133200 535810
rect 133660 535680 133800 535810
<< nsubdiffcont >>
rect 119540 593100 119580 593260
rect 120210 593100 120250 593260
rect 119580 583560 119620 583720
rect 120250 583560 120290 583720
rect 119620 574540 119660 574700
rect 120290 574540 120330 574700
rect 119570 566870 119610 567030
rect 120240 566870 120280 567030
rect 119570 560330 119610 560490
rect 120240 560330 120280 560490
rect 119640 553500 119680 553660
rect 120310 553500 120350 553660
rect 119640 545930 119680 546090
rect 120310 545930 120350 546090
rect 119610 537870 119650 538030
rect 120280 537870 120320 538030
<< poly >>
rect 124020 642750 124100 642770
rect 124020 642710 124040 642750
rect 124080 642740 124100 642750
rect 124080 642710 124130 642740
rect 124020 642690 124130 642710
rect 124100 642340 124130 642690
rect 124100 642310 124150 642340
rect 124240 642310 124330 642340
rect 124420 642310 124510 642340
rect 124600 642310 124690 642340
rect 124780 642310 124870 642340
rect 124960 642310 125050 642340
rect 125140 642310 125230 642340
rect 125320 642310 125410 642340
rect 125500 642310 125590 642340
rect 125680 642310 125770 642340
rect 125860 642310 125950 642340
rect 126040 642310 126130 642340
rect 126220 642310 126310 642340
rect 126400 642310 126490 642340
rect 126580 642310 126670 642340
rect 126760 642310 126850 642340
rect 126940 642310 127030 642340
rect 127120 642310 127210 642340
rect 127300 642310 127390 642340
rect 127480 642310 127570 642340
rect 127660 642310 127750 642340
rect 127840 642310 127930 642340
rect 128020 642310 128110 642340
rect 128200 642310 128290 642340
rect 128380 642310 128470 642340
rect 128560 642310 128650 642340
rect 128740 642310 128830 642340
rect 128920 642310 129010 642340
rect 129100 642310 129190 642340
rect 129280 642310 129370 642340
rect 129460 642310 129550 642340
rect 129640 642310 129730 642340
rect 129820 642310 129910 642340
rect 130000 642310 130090 642340
rect 130180 642310 130270 642340
rect 130360 642310 130450 642340
rect 130540 642310 130630 642340
rect 130720 642310 130810 642340
rect 130900 642310 130990 642340
rect 131080 642310 131170 642340
rect 131260 642310 131350 642340
rect 124050 636170 124130 636190
rect 124050 636130 124070 636170
rect 124110 636140 124180 636170
rect 124360 636140 124420 636170
rect 124600 636140 124660 636170
rect 124840 636140 124900 636170
rect 125080 636140 125140 636170
rect 125320 636140 125380 636170
rect 125560 636140 125620 636170
rect 125800 636140 125860 636170
rect 126040 636140 126100 636170
rect 126280 636140 126340 636170
rect 126520 636140 126580 636170
rect 126760 636140 126820 636170
rect 127000 636140 127060 636170
rect 127240 636140 127300 636170
rect 127480 636140 127540 636170
rect 127720 636140 127780 636170
rect 127960 636140 128020 636170
rect 128200 636140 128260 636170
rect 128440 636140 128500 636170
rect 128680 636140 128740 636170
rect 128920 636140 128980 636170
rect 124110 636130 124130 636140
rect 124050 636110 124130 636130
rect 124180 632550 124240 632580
rect 124640 632550 124700 632580
rect 124330 630140 124410 630160
rect 124330 630100 124350 630140
rect 124390 630110 124450 630140
rect 124850 630110 124910 630140
rect 125310 630110 125370 630140
rect 125770 630110 125830 630140
rect 126230 630110 126290 630140
rect 126690 630110 126750 630140
rect 127150 630110 127210 630140
rect 127610 630110 127670 630140
rect 128070 630110 128130 630140
rect 128530 630110 128590 630140
rect 128990 630110 129050 630140
rect 124390 630100 124410 630110
rect 124330 630080 124410 630100
rect 124160 624880 124220 624910
rect 124820 624880 124880 624910
rect 124580 624010 124660 624030
rect 124580 623970 124600 624010
rect 124640 623970 124690 624010
rect 124580 623950 124690 623970
rect 124660 623620 124690 623950
rect 124660 623590 124780 623620
rect 125380 623590 125440 623620
rect 126040 623590 126100 623620
rect 126700 623590 126760 623620
rect 127360 623590 127420 623620
rect 128020 623590 128080 623620
rect 128680 623590 128740 623620
rect 125510 619550 125570 619570
rect 125510 619510 125520 619550
rect 125560 619510 125570 619550
rect 125510 619490 125570 619510
rect 125530 619450 125560 619490
rect 125580 618770 125640 618790
rect 125580 618730 125590 618770
rect 125630 618730 125640 618770
rect 125580 618710 125640 618730
rect 125920 618770 125980 618790
rect 125920 618730 125930 618770
rect 125970 618730 125980 618770
rect 125920 618710 125980 618730
rect 126260 618770 126320 618790
rect 126260 618730 126270 618770
rect 126310 618730 126320 618770
rect 126260 618710 126320 618730
rect 126600 618770 126660 618790
rect 126600 618730 126610 618770
rect 126650 618730 126660 618770
rect 126600 618710 126660 618730
rect 126940 618770 127000 618790
rect 126940 618730 126950 618770
rect 126990 618730 127000 618770
rect 126940 618710 127000 618730
rect 127280 618770 127340 618790
rect 127280 618730 127290 618770
rect 127330 618730 127340 618770
rect 127280 618710 127340 618730
rect 127620 618770 127680 618790
rect 127620 618730 127630 618770
rect 127670 618730 127680 618770
rect 127620 618710 127680 618730
rect 127960 618770 128020 618790
rect 127960 618730 127970 618770
rect 128010 618730 128020 618770
rect 127960 618710 128020 618730
rect 128300 618770 128360 618790
rect 128300 618730 128310 618770
rect 128350 618730 128360 618770
rect 128300 618710 128360 618730
rect 128640 618770 128700 618790
rect 128640 618730 128650 618770
rect 128690 618730 128700 618770
rect 128640 618710 128700 618730
rect 128980 618770 129040 618790
rect 128980 618730 128990 618770
rect 129030 618730 129040 618770
rect 128980 618710 129040 618730
rect 129320 618770 129380 618790
rect 129320 618730 129330 618770
rect 129370 618730 129380 618770
rect 129320 618710 129380 618730
rect 129660 618770 129720 618790
rect 129660 618730 129670 618770
rect 129710 618730 129720 618770
rect 129660 618710 129720 618730
rect 130000 618770 130060 618790
rect 130000 618730 130010 618770
rect 130050 618730 130060 618770
rect 130000 618710 130060 618730
rect 130340 618770 130400 618790
rect 130340 618730 130350 618770
rect 130390 618730 130400 618770
rect 130340 618710 130400 618730
rect 130680 618770 130740 618790
rect 130680 618730 130690 618770
rect 130730 618730 130740 618770
rect 130680 618710 130740 618730
rect 131020 618770 131080 618790
rect 131020 618730 131030 618770
rect 131070 618730 131080 618770
rect 131020 618710 131080 618730
rect 131360 618770 131420 618790
rect 131360 618730 131370 618770
rect 131410 618730 131420 618770
rect 131360 618710 131420 618730
rect 131700 618770 131760 618790
rect 131700 618730 131710 618770
rect 131750 618730 131760 618770
rect 131700 618710 131760 618730
rect 125600 618670 125630 618710
rect 125940 618670 125970 618710
rect 126280 618670 126310 618710
rect 126620 618670 126650 618710
rect 126960 618670 126990 618710
rect 127300 618670 127330 618710
rect 127640 618670 127670 618710
rect 127980 618670 128010 618710
rect 128320 618670 128350 618710
rect 128660 618670 128690 618710
rect 129000 618670 129030 618710
rect 129340 618670 129370 618710
rect 129680 618670 129710 618710
rect 130020 618670 130050 618710
rect 130360 618670 130390 618710
rect 130700 618670 130730 618710
rect 131040 618670 131070 618710
rect 131380 618670 131410 618710
rect 131720 618670 131750 618710
rect 125160 612100 125220 612120
rect 125160 612060 125170 612100
rect 125210 612060 125220 612100
rect 125160 612040 125220 612060
rect 125180 612000 125210 612040
rect 125230 611320 125290 611340
rect 125230 611280 125240 611320
rect 125280 611280 125290 611320
rect 125230 611260 125290 611280
rect 125570 611320 125630 611340
rect 125570 611280 125580 611320
rect 125620 611280 125630 611320
rect 125570 611260 125630 611280
rect 125910 611320 125970 611340
rect 125910 611280 125920 611320
rect 125960 611280 125970 611320
rect 125910 611260 125970 611280
rect 126250 611320 126310 611340
rect 126250 611280 126260 611320
rect 126300 611280 126310 611320
rect 126250 611260 126310 611280
rect 126590 611320 126650 611340
rect 126590 611280 126600 611320
rect 126640 611280 126650 611320
rect 126590 611260 126650 611280
rect 126930 611320 126990 611340
rect 126930 611280 126940 611320
rect 126980 611280 126990 611320
rect 126930 611260 126990 611280
rect 127270 611320 127330 611340
rect 127270 611280 127280 611320
rect 127320 611280 127330 611320
rect 127270 611260 127330 611280
rect 127610 611320 127670 611340
rect 127610 611280 127620 611320
rect 127660 611280 127670 611320
rect 127610 611260 127670 611280
rect 127950 611320 128010 611340
rect 127950 611280 127960 611320
rect 128000 611280 128010 611320
rect 127950 611260 128010 611280
rect 128290 611320 128350 611340
rect 128290 611280 128300 611320
rect 128340 611280 128350 611320
rect 128290 611260 128350 611280
rect 128630 611320 128690 611340
rect 128630 611280 128640 611320
rect 128680 611280 128690 611320
rect 128630 611260 128690 611280
rect 128970 611320 129030 611340
rect 128970 611280 128980 611320
rect 129020 611280 129030 611320
rect 128970 611260 129030 611280
rect 129310 611320 129370 611340
rect 129310 611280 129320 611320
rect 129360 611280 129370 611320
rect 129310 611260 129370 611280
rect 129650 611320 129710 611340
rect 129650 611280 129660 611320
rect 129700 611280 129710 611320
rect 129650 611260 129710 611280
rect 129990 611320 130050 611340
rect 129990 611280 130000 611320
rect 130040 611280 130050 611320
rect 129990 611260 130050 611280
rect 130330 611320 130390 611340
rect 130330 611280 130340 611320
rect 130380 611280 130390 611320
rect 130330 611260 130390 611280
rect 130670 611320 130730 611340
rect 130670 611280 130680 611320
rect 130720 611280 130730 611320
rect 130670 611260 130730 611280
rect 131010 611320 131070 611340
rect 131010 611280 131020 611320
rect 131060 611280 131070 611320
rect 131010 611260 131070 611280
rect 131350 611320 131410 611340
rect 131350 611280 131360 611320
rect 131400 611280 131410 611320
rect 131350 611260 131410 611280
rect 125250 611220 125280 611260
rect 125590 611220 125620 611260
rect 125930 611220 125960 611260
rect 126270 611220 126300 611260
rect 126610 611220 126640 611260
rect 126950 611220 126980 611260
rect 127290 611220 127320 611260
rect 127630 611220 127660 611260
rect 127970 611220 128000 611260
rect 128310 611220 128340 611260
rect 128650 611220 128680 611260
rect 128990 611220 129020 611260
rect 129330 611220 129360 611260
rect 129670 611220 129700 611260
rect 130010 611220 130040 611260
rect 130350 611220 130380 611260
rect 130690 611220 130720 611260
rect 131030 611220 131060 611260
rect 131370 611220 131400 611260
rect 125290 606050 125350 606070
rect 125290 606010 125300 606050
rect 125340 606010 125350 606050
rect 125290 605990 125350 606010
rect 125310 605950 125340 605990
rect 125360 605270 125420 605290
rect 125360 605230 125370 605270
rect 125410 605230 125420 605270
rect 125360 605210 125420 605230
rect 125700 605270 125760 605290
rect 125700 605230 125710 605270
rect 125750 605230 125760 605270
rect 125700 605210 125760 605230
rect 126040 605270 126100 605290
rect 126040 605230 126050 605270
rect 126090 605230 126100 605270
rect 126040 605210 126100 605230
rect 126380 605270 126440 605290
rect 126380 605230 126390 605270
rect 126430 605230 126440 605270
rect 126380 605210 126440 605230
rect 126720 605270 126780 605290
rect 126720 605230 126730 605270
rect 126770 605230 126780 605270
rect 126720 605210 126780 605230
rect 127060 605270 127120 605290
rect 127060 605230 127070 605270
rect 127110 605230 127120 605270
rect 127060 605210 127120 605230
rect 127400 605270 127460 605290
rect 127400 605230 127410 605270
rect 127450 605230 127460 605270
rect 127400 605210 127460 605230
rect 127740 605270 127800 605290
rect 127740 605230 127750 605270
rect 127790 605230 127800 605270
rect 127740 605210 127800 605230
rect 128080 605270 128140 605290
rect 128080 605230 128090 605270
rect 128130 605230 128140 605270
rect 128080 605210 128140 605230
rect 128420 605270 128480 605290
rect 128420 605230 128430 605270
rect 128470 605230 128480 605270
rect 128420 605210 128480 605230
rect 128760 605270 128820 605290
rect 128760 605230 128770 605270
rect 128810 605230 128820 605270
rect 128760 605210 128820 605230
rect 129100 605270 129160 605290
rect 129100 605230 129110 605270
rect 129150 605230 129160 605270
rect 129100 605210 129160 605230
rect 129440 605270 129500 605290
rect 129440 605230 129450 605270
rect 129490 605230 129500 605270
rect 129440 605210 129500 605230
rect 129780 605270 129840 605290
rect 129780 605230 129790 605270
rect 129830 605230 129840 605270
rect 129780 605210 129840 605230
rect 130120 605270 130180 605290
rect 130120 605230 130130 605270
rect 130170 605230 130180 605270
rect 130120 605210 130180 605230
rect 130460 605270 130520 605290
rect 130460 605230 130470 605270
rect 130510 605230 130520 605270
rect 130460 605210 130520 605230
rect 130800 605270 130860 605290
rect 130800 605230 130810 605270
rect 130850 605230 130860 605270
rect 130800 605210 130860 605230
rect 131140 605270 131200 605290
rect 131140 605230 131150 605270
rect 131190 605230 131200 605270
rect 131140 605210 131200 605230
rect 131480 605270 131540 605290
rect 131480 605230 131490 605270
rect 131530 605230 131540 605270
rect 131480 605210 131540 605230
rect 125380 605170 125410 605210
rect 125720 605170 125750 605210
rect 126060 605170 126090 605210
rect 126400 605170 126430 605210
rect 126740 605170 126770 605210
rect 127080 605170 127110 605210
rect 127420 605170 127450 605210
rect 127760 605170 127790 605210
rect 128100 605170 128130 605210
rect 128440 605170 128470 605210
rect 128780 605170 128810 605210
rect 129120 605170 129150 605210
rect 129460 605170 129490 605210
rect 129800 605170 129830 605210
rect 130140 605170 130170 605210
rect 130480 605170 130510 605210
rect 130820 605170 130850 605210
rect 131160 605170 131190 605210
rect 131500 605170 131530 605210
rect 125090 599790 125150 599810
rect 125090 599750 125100 599790
rect 125140 599750 125150 599790
rect 125090 599730 125150 599750
rect 125110 599690 125140 599730
rect 125160 599010 125220 599030
rect 125160 598970 125170 599010
rect 125210 598970 125220 599010
rect 125160 598950 125220 598970
rect 125500 599010 125560 599030
rect 125500 598970 125510 599010
rect 125550 598970 125560 599010
rect 125500 598950 125560 598970
rect 125840 599010 125900 599030
rect 125840 598970 125850 599010
rect 125890 598970 125900 599010
rect 125840 598950 125900 598970
rect 126180 599010 126240 599030
rect 126180 598970 126190 599010
rect 126230 598970 126240 599010
rect 126180 598950 126240 598970
rect 126520 599010 126580 599030
rect 126520 598970 126530 599010
rect 126570 598970 126580 599010
rect 126520 598950 126580 598970
rect 126860 599010 126920 599030
rect 126860 598970 126870 599010
rect 126910 598970 126920 599010
rect 126860 598950 126920 598970
rect 127200 599010 127260 599030
rect 127200 598970 127210 599010
rect 127250 598970 127260 599010
rect 127200 598950 127260 598970
rect 127540 599010 127600 599030
rect 127540 598970 127550 599010
rect 127590 598970 127600 599010
rect 127540 598950 127600 598970
rect 127880 599010 127940 599030
rect 127880 598970 127890 599010
rect 127930 598970 127940 599010
rect 127880 598950 127940 598970
rect 128220 599010 128280 599030
rect 128220 598970 128230 599010
rect 128270 598970 128280 599010
rect 128220 598950 128280 598970
rect 128560 599010 128620 599030
rect 128560 598970 128570 599010
rect 128610 598970 128620 599010
rect 128560 598950 128620 598970
rect 128900 599010 128960 599030
rect 128900 598970 128910 599010
rect 128950 598970 128960 599010
rect 128900 598950 128960 598970
rect 129240 599010 129300 599030
rect 129240 598970 129250 599010
rect 129290 598970 129300 599010
rect 129240 598950 129300 598970
rect 129580 599010 129640 599030
rect 129580 598970 129590 599010
rect 129630 598970 129640 599010
rect 129580 598950 129640 598970
rect 129920 599010 129980 599030
rect 129920 598970 129930 599010
rect 129970 598970 129980 599010
rect 129920 598950 129980 598970
rect 130260 599010 130320 599030
rect 130260 598970 130270 599010
rect 130310 598970 130320 599010
rect 130260 598950 130320 598970
rect 130600 599010 130660 599030
rect 130600 598970 130610 599010
rect 130650 598970 130660 599010
rect 130600 598950 130660 598970
rect 130940 599010 131000 599030
rect 130940 598970 130950 599010
rect 130990 598970 131000 599010
rect 130940 598950 131000 598970
rect 131280 599010 131340 599030
rect 131280 598970 131290 599010
rect 131330 598970 131340 599010
rect 131280 598950 131340 598970
rect 125180 598910 125210 598950
rect 125520 598910 125550 598950
rect 125860 598910 125890 598950
rect 126200 598910 126230 598950
rect 126540 598910 126570 598950
rect 126880 598910 126910 598950
rect 127220 598910 127250 598950
rect 127560 598910 127590 598950
rect 127900 598910 127930 598950
rect 128240 598910 128270 598950
rect 128580 598910 128610 598950
rect 128920 598910 128950 598950
rect 129260 598910 129290 598950
rect 129600 598910 129630 598950
rect 129940 598910 129970 598950
rect 130280 598910 130310 598950
rect 130620 598910 130650 598950
rect 130960 598910 130990 598950
rect 131300 598910 131330 598950
rect 119100 593420 119180 593440
rect 119100 593380 119120 593420
rect 119160 593410 119180 593420
rect 119160 593380 120100 593410
rect 119100 593360 119180 593380
rect 119330 593250 119360 593380
rect 119690 593280 119720 593310
rect 120070 593280 120100 593380
rect 119330 592970 119360 593160
rect 119470 593020 119550 593040
rect 119690 593020 119720 593080
rect 119850 593030 119930 593050
rect 119850 593020 119870 593030
rect 119470 592980 119490 593020
rect 119530 592990 119870 593020
rect 119910 592990 119930 593030
rect 119530 592980 119550 592990
rect 119470 592960 119550 592980
rect 119850 592970 119930 592990
rect 120070 592920 120100 593080
rect 120220 593020 120300 593040
rect 120220 592980 120240 593020
rect 120280 592980 120300 593020
rect 120220 592960 120300 592980
rect 119690 592890 120100 592920
rect 119330 592850 119360 592880
rect 119690 592770 119720 592890
rect 120240 592840 120270 592960
rect 120070 592810 120270 592840
rect 120070 592770 120100 592810
rect 119690 592540 119720 592570
rect 120070 592540 120100 592570
rect 125050 592240 125110 592260
rect 125050 592200 125060 592240
rect 125100 592200 125110 592240
rect 125050 592180 125110 592200
rect 125070 592140 125100 592180
rect 125120 591460 125180 591480
rect 125120 591420 125130 591460
rect 125170 591420 125180 591460
rect 125120 591400 125180 591420
rect 125460 591460 125520 591480
rect 125460 591420 125470 591460
rect 125510 591420 125520 591460
rect 125460 591400 125520 591420
rect 125800 591460 125860 591480
rect 125800 591420 125810 591460
rect 125850 591420 125860 591460
rect 125800 591400 125860 591420
rect 126140 591460 126200 591480
rect 126140 591420 126150 591460
rect 126190 591420 126200 591460
rect 126140 591400 126200 591420
rect 126480 591460 126540 591480
rect 126480 591420 126490 591460
rect 126530 591420 126540 591460
rect 126480 591400 126540 591420
rect 126820 591460 126880 591480
rect 126820 591420 126830 591460
rect 126870 591420 126880 591460
rect 126820 591400 126880 591420
rect 127160 591460 127220 591480
rect 127160 591420 127170 591460
rect 127210 591420 127220 591460
rect 127160 591400 127220 591420
rect 127500 591460 127560 591480
rect 127500 591420 127510 591460
rect 127550 591420 127560 591460
rect 127500 591400 127560 591420
rect 127840 591460 127900 591480
rect 127840 591420 127850 591460
rect 127890 591420 127900 591460
rect 127840 591400 127900 591420
rect 128180 591460 128240 591480
rect 128180 591420 128190 591460
rect 128230 591420 128240 591460
rect 128180 591400 128240 591420
rect 128520 591460 128580 591480
rect 128520 591420 128530 591460
rect 128570 591420 128580 591460
rect 128520 591400 128580 591420
rect 128860 591460 128920 591480
rect 128860 591420 128870 591460
rect 128910 591420 128920 591460
rect 128860 591400 128920 591420
rect 129200 591460 129260 591480
rect 129200 591420 129210 591460
rect 129250 591420 129260 591460
rect 129200 591400 129260 591420
rect 129540 591460 129600 591480
rect 129540 591420 129550 591460
rect 129590 591420 129600 591460
rect 129540 591400 129600 591420
rect 129880 591460 129940 591480
rect 129880 591420 129890 591460
rect 129930 591420 129940 591460
rect 129880 591400 129940 591420
rect 130220 591460 130280 591480
rect 130220 591420 130230 591460
rect 130270 591420 130280 591460
rect 130220 591400 130280 591420
rect 130560 591460 130620 591480
rect 130560 591420 130570 591460
rect 130610 591420 130620 591460
rect 130560 591400 130620 591420
rect 130900 591460 130960 591480
rect 130900 591420 130910 591460
rect 130950 591420 130960 591460
rect 130900 591400 130960 591420
rect 131240 591460 131300 591480
rect 131240 591420 131250 591460
rect 131290 591420 131300 591460
rect 131240 591400 131300 591420
rect 125140 591360 125170 591400
rect 125480 591360 125510 591400
rect 125820 591360 125850 591400
rect 126160 591360 126190 591400
rect 126500 591360 126530 591400
rect 126840 591360 126870 591400
rect 127180 591360 127210 591400
rect 127520 591360 127550 591400
rect 127860 591360 127890 591400
rect 128200 591360 128230 591400
rect 128540 591360 128570 591400
rect 128880 591360 128910 591400
rect 129220 591360 129250 591400
rect 129560 591360 129590 591400
rect 129900 591360 129930 591400
rect 130240 591360 130270 591400
rect 130580 591360 130610 591400
rect 130920 591360 130950 591400
rect 131260 591360 131290 591400
rect 119140 583880 119220 583900
rect 119140 583840 119160 583880
rect 119200 583870 119220 583880
rect 119200 583840 120140 583870
rect 119140 583820 119220 583840
rect 119370 583710 119400 583840
rect 119730 583740 119760 583770
rect 120110 583740 120140 583840
rect 119370 583430 119400 583620
rect 119510 583480 119590 583500
rect 119730 583480 119760 583540
rect 119890 583490 119970 583510
rect 119890 583480 119910 583490
rect 119510 583440 119530 583480
rect 119570 583450 119910 583480
rect 119950 583450 119970 583490
rect 119570 583440 119590 583450
rect 119510 583420 119590 583440
rect 119890 583430 119970 583450
rect 120110 583380 120140 583540
rect 120260 583480 120340 583500
rect 120260 583440 120280 583480
rect 120320 583440 120340 583480
rect 120260 583420 120340 583440
rect 119730 583350 120140 583380
rect 119370 583310 119400 583340
rect 119730 583230 119760 583350
rect 120280 583300 120310 583420
rect 120110 583270 120310 583300
rect 120110 583230 120140 583270
rect 125510 583260 125570 583280
rect 125510 583220 125520 583260
rect 125560 583220 125570 583260
rect 125510 583200 125570 583220
rect 125530 583160 125560 583200
rect 119730 583000 119760 583030
rect 120110 583000 120140 583030
rect 125630 582480 125690 582500
rect 125630 582440 125640 582480
rect 125680 582440 125690 582480
rect 125630 582420 125690 582440
rect 126020 582480 126080 582500
rect 126020 582440 126030 582480
rect 126070 582440 126080 582480
rect 126020 582420 126080 582440
rect 126410 582480 126470 582500
rect 126410 582440 126420 582480
rect 126460 582440 126470 582480
rect 126410 582420 126470 582440
rect 126800 582480 126860 582500
rect 126800 582440 126810 582480
rect 126850 582440 126860 582480
rect 126800 582420 126860 582440
rect 127190 582480 127250 582500
rect 127190 582440 127200 582480
rect 127240 582440 127250 582480
rect 127190 582420 127250 582440
rect 127580 582480 127640 582500
rect 127580 582440 127590 582480
rect 127630 582440 127640 582480
rect 127580 582420 127640 582440
rect 127970 582480 128030 582500
rect 127970 582440 127980 582480
rect 128020 582440 128030 582480
rect 127970 582420 128030 582440
rect 128360 582480 128420 582500
rect 128360 582440 128370 582480
rect 128410 582440 128420 582480
rect 128360 582420 128420 582440
rect 128750 582480 128810 582500
rect 128750 582440 128760 582480
rect 128800 582440 128810 582480
rect 128750 582420 128810 582440
rect 129140 582480 129200 582500
rect 129140 582440 129150 582480
rect 129190 582440 129200 582480
rect 129140 582420 129200 582440
rect 129530 582480 129590 582500
rect 129530 582440 129540 582480
rect 129580 582440 129590 582480
rect 129530 582420 129590 582440
rect 129920 582480 129980 582500
rect 129920 582440 129930 582480
rect 129970 582440 129980 582480
rect 129920 582420 129980 582440
rect 130310 582480 130370 582500
rect 130310 582440 130320 582480
rect 130360 582440 130370 582480
rect 130310 582420 130370 582440
rect 130700 582480 130760 582500
rect 130700 582440 130710 582480
rect 130750 582440 130760 582480
rect 130700 582420 130760 582440
rect 131090 582480 131150 582500
rect 131090 582440 131100 582480
rect 131140 582440 131150 582480
rect 131090 582420 131150 582440
rect 131480 582480 131540 582500
rect 131480 582440 131490 582480
rect 131530 582440 131540 582480
rect 131480 582420 131540 582440
rect 131870 582480 131930 582500
rect 131870 582440 131880 582480
rect 131920 582440 131930 582480
rect 131870 582420 131930 582440
rect 132260 582480 132320 582500
rect 132260 582440 132270 582480
rect 132310 582440 132320 582480
rect 132260 582420 132320 582440
rect 132650 582480 132710 582500
rect 132650 582440 132660 582480
rect 132700 582440 132710 582480
rect 132650 582420 132710 582440
rect 125650 582380 125680 582420
rect 126040 582380 126070 582420
rect 126430 582380 126460 582420
rect 126820 582380 126850 582420
rect 127210 582380 127240 582420
rect 127600 582380 127630 582420
rect 127990 582380 128020 582420
rect 128380 582380 128410 582420
rect 128770 582380 128800 582420
rect 129160 582380 129190 582420
rect 129550 582380 129580 582420
rect 129940 582380 129970 582420
rect 130330 582380 130360 582420
rect 130720 582380 130750 582420
rect 131110 582380 131140 582420
rect 131500 582380 131530 582420
rect 131890 582380 131920 582420
rect 132280 582380 132310 582420
rect 132670 582380 132700 582420
rect 119180 574860 119260 574880
rect 119180 574820 119200 574860
rect 119240 574850 119260 574860
rect 119240 574820 120180 574850
rect 119180 574800 119260 574820
rect 119410 574690 119440 574820
rect 119770 574720 119800 574750
rect 120150 574720 120180 574820
rect 119410 574410 119440 574600
rect 119550 574460 119630 574480
rect 119770 574460 119800 574520
rect 119930 574470 120010 574490
rect 119930 574460 119950 574470
rect 119550 574420 119570 574460
rect 119610 574430 119950 574460
rect 119990 574430 120010 574470
rect 119610 574420 119630 574430
rect 119550 574400 119630 574420
rect 119930 574410 120010 574430
rect 120150 574360 120180 574520
rect 120300 574460 120380 574480
rect 120300 574420 120320 574460
rect 120360 574420 120380 574460
rect 120300 574400 120380 574420
rect 119770 574330 120180 574360
rect 119410 574290 119440 574320
rect 119770 574210 119800 574330
rect 120320 574280 120350 574400
rect 120150 574250 120350 574280
rect 120150 574210 120180 574250
rect 125550 574240 125610 574260
rect 125550 574200 125560 574240
rect 125600 574200 125610 574240
rect 125550 574180 125610 574200
rect 125570 574140 125600 574180
rect 119770 573980 119800 574010
rect 120150 573980 120180 574010
rect 125670 573460 125730 573480
rect 125670 573420 125680 573460
rect 125720 573420 125730 573460
rect 125670 573400 125730 573420
rect 126060 573460 126120 573480
rect 126060 573420 126070 573460
rect 126110 573420 126120 573460
rect 126060 573400 126120 573420
rect 126450 573460 126510 573480
rect 126450 573420 126460 573460
rect 126500 573420 126510 573460
rect 126450 573400 126510 573420
rect 126840 573460 126900 573480
rect 126840 573420 126850 573460
rect 126890 573420 126900 573460
rect 126840 573400 126900 573420
rect 127230 573460 127290 573480
rect 127230 573420 127240 573460
rect 127280 573420 127290 573460
rect 127230 573400 127290 573420
rect 127620 573460 127680 573480
rect 127620 573420 127630 573460
rect 127670 573420 127680 573460
rect 127620 573400 127680 573420
rect 128010 573460 128070 573480
rect 128010 573420 128020 573460
rect 128060 573420 128070 573460
rect 128010 573400 128070 573420
rect 128400 573460 128460 573480
rect 128400 573420 128410 573460
rect 128450 573420 128460 573460
rect 128400 573400 128460 573420
rect 128790 573460 128850 573480
rect 128790 573420 128800 573460
rect 128840 573420 128850 573460
rect 128790 573400 128850 573420
rect 129180 573460 129240 573480
rect 129180 573420 129190 573460
rect 129230 573420 129240 573460
rect 129180 573400 129240 573420
rect 129570 573460 129630 573480
rect 129570 573420 129580 573460
rect 129620 573420 129630 573460
rect 129570 573400 129630 573420
rect 129960 573460 130020 573480
rect 129960 573420 129970 573460
rect 130010 573420 130020 573460
rect 129960 573400 130020 573420
rect 130350 573460 130410 573480
rect 130350 573420 130360 573460
rect 130400 573420 130410 573460
rect 130350 573400 130410 573420
rect 130740 573460 130800 573480
rect 130740 573420 130750 573460
rect 130790 573420 130800 573460
rect 130740 573400 130800 573420
rect 131130 573460 131190 573480
rect 131130 573420 131140 573460
rect 131180 573420 131190 573460
rect 131130 573400 131190 573420
rect 131520 573460 131580 573480
rect 131520 573420 131530 573460
rect 131570 573420 131580 573460
rect 131520 573400 131580 573420
rect 131910 573460 131970 573480
rect 131910 573420 131920 573460
rect 131960 573420 131970 573460
rect 131910 573400 131970 573420
rect 132300 573460 132360 573480
rect 132300 573420 132310 573460
rect 132350 573420 132360 573460
rect 132300 573400 132360 573420
rect 132690 573460 132750 573480
rect 132690 573420 132700 573460
rect 132740 573420 132750 573460
rect 132690 573400 132750 573420
rect 125690 573360 125720 573400
rect 126080 573360 126110 573400
rect 126470 573360 126500 573400
rect 126860 573360 126890 573400
rect 127250 573360 127280 573400
rect 127640 573360 127670 573400
rect 128030 573360 128060 573400
rect 128420 573360 128450 573400
rect 128810 573360 128840 573400
rect 129200 573360 129230 573400
rect 129590 573360 129620 573400
rect 129980 573360 130010 573400
rect 130370 573360 130400 573400
rect 130760 573360 130790 573400
rect 131150 573360 131180 573400
rect 131540 573360 131570 573400
rect 131930 573360 131960 573400
rect 132320 573360 132350 573400
rect 132710 573360 132740 573400
rect 119130 567190 119210 567210
rect 119130 567150 119150 567190
rect 119190 567180 119210 567190
rect 119190 567150 120130 567180
rect 119130 567130 119210 567150
rect 119360 567020 119390 567150
rect 119720 567050 119750 567080
rect 120100 567050 120130 567150
rect 119360 566740 119390 566930
rect 119500 566790 119580 566810
rect 119720 566790 119750 566850
rect 119880 566800 119960 566820
rect 119880 566790 119900 566800
rect 119500 566750 119520 566790
rect 119560 566760 119900 566790
rect 119940 566760 119960 566800
rect 119560 566750 119580 566760
rect 119500 566730 119580 566750
rect 119880 566740 119960 566760
rect 120100 566690 120130 566850
rect 120250 566790 120330 566810
rect 120250 566750 120270 566790
rect 120310 566750 120330 566790
rect 120250 566730 120330 566750
rect 119720 566660 120130 566690
rect 119360 566620 119390 566650
rect 119720 566540 119750 566660
rect 120270 566610 120300 566730
rect 120100 566580 120300 566610
rect 120100 566540 120130 566580
rect 125500 566570 125560 566590
rect 125500 566530 125510 566570
rect 125550 566530 125560 566570
rect 125500 566510 125560 566530
rect 125520 566470 125550 566510
rect 119720 566310 119750 566340
rect 120100 566310 120130 566340
rect 125620 565790 125680 565810
rect 125620 565750 125630 565790
rect 125670 565750 125680 565790
rect 125620 565730 125680 565750
rect 126010 565790 126070 565810
rect 126010 565750 126020 565790
rect 126060 565750 126070 565790
rect 126010 565730 126070 565750
rect 126400 565790 126460 565810
rect 126400 565750 126410 565790
rect 126450 565750 126460 565790
rect 126400 565730 126460 565750
rect 126790 565790 126850 565810
rect 126790 565750 126800 565790
rect 126840 565750 126850 565790
rect 126790 565730 126850 565750
rect 127180 565790 127240 565810
rect 127180 565750 127190 565790
rect 127230 565750 127240 565790
rect 127180 565730 127240 565750
rect 127570 565790 127630 565810
rect 127570 565750 127580 565790
rect 127620 565750 127630 565790
rect 127570 565730 127630 565750
rect 127960 565790 128020 565810
rect 127960 565750 127970 565790
rect 128010 565750 128020 565790
rect 127960 565730 128020 565750
rect 128350 565790 128410 565810
rect 128350 565750 128360 565790
rect 128400 565750 128410 565790
rect 128350 565730 128410 565750
rect 128740 565790 128800 565810
rect 128740 565750 128750 565790
rect 128790 565750 128800 565790
rect 128740 565730 128800 565750
rect 129130 565790 129190 565810
rect 129130 565750 129140 565790
rect 129180 565750 129190 565790
rect 129130 565730 129190 565750
rect 129520 565790 129580 565810
rect 129520 565750 129530 565790
rect 129570 565750 129580 565790
rect 129520 565730 129580 565750
rect 129910 565790 129970 565810
rect 129910 565750 129920 565790
rect 129960 565750 129970 565790
rect 129910 565730 129970 565750
rect 130300 565790 130360 565810
rect 130300 565750 130310 565790
rect 130350 565750 130360 565790
rect 130300 565730 130360 565750
rect 130690 565790 130750 565810
rect 130690 565750 130700 565790
rect 130740 565750 130750 565790
rect 130690 565730 130750 565750
rect 131080 565790 131140 565810
rect 131080 565750 131090 565790
rect 131130 565750 131140 565790
rect 131080 565730 131140 565750
rect 131470 565790 131530 565810
rect 131470 565750 131480 565790
rect 131520 565750 131530 565790
rect 131470 565730 131530 565750
rect 131860 565790 131920 565810
rect 131860 565750 131870 565790
rect 131910 565750 131920 565790
rect 131860 565730 131920 565750
rect 132250 565790 132310 565810
rect 132250 565750 132260 565790
rect 132300 565750 132310 565790
rect 132250 565730 132310 565750
rect 132640 565790 132700 565810
rect 132640 565750 132650 565790
rect 132690 565750 132700 565790
rect 132640 565730 132700 565750
rect 125640 565690 125670 565730
rect 126030 565690 126060 565730
rect 126420 565690 126450 565730
rect 126810 565690 126840 565730
rect 127200 565690 127230 565730
rect 127590 565690 127620 565730
rect 127980 565690 128010 565730
rect 128370 565690 128400 565730
rect 128760 565690 128790 565730
rect 129150 565690 129180 565730
rect 129540 565690 129570 565730
rect 129930 565690 129960 565730
rect 130320 565690 130350 565730
rect 130710 565690 130740 565730
rect 131100 565690 131130 565730
rect 131490 565690 131520 565730
rect 131880 565690 131910 565730
rect 132270 565690 132300 565730
rect 132660 565690 132690 565730
rect 119130 560650 119210 560670
rect 119130 560610 119150 560650
rect 119190 560640 119210 560650
rect 119190 560610 120130 560640
rect 119130 560590 119210 560610
rect 119360 560480 119390 560610
rect 119720 560510 119750 560540
rect 120100 560510 120130 560610
rect 119360 560200 119390 560390
rect 119500 560250 119580 560270
rect 119720 560250 119750 560310
rect 119880 560260 119960 560280
rect 119880 560250 119900 560260
rect 119500 560210 119520 560250
rect 119560 560220 119900 560250
rect 119940 560220 119960 560260
rect 119560 560210 119580 560220
rect 119500 560190 119580 560210
rect 119880 560200 119960 560220
rect 120100 560150 120130 560310
rect 120250 560250 120330 560270
rect 120250 560210 120270 560250
rect 120310 560210 120330 560250
rect 120250 560190 120330 560210
rect 119720 560120 120130 560150
rect 119360 560080 119390 560110
rect 119720 560000 119750 560120
rect 120270 560070 120300 560190
rect 120100 560040 120300 560070
rect 120100 560000 120130 560040
rect 125500 560030 125560 560050
rect 125500 559990 125510 560030
rect 125550 559990 125560 560030
rect 125500 559970 125560 559990
rect 125520 559930 125550 559970
rect 119720 559770 119750 559800
rect 120100 559770 120130 559800
rect 125620 559250 125680 559270
rect 125620 559210 125630 559250
rect 125670 559210 125680 559250
rect 125620 559190 125680 559210
rect 126010 559250 126070 559270
rect 126010 559210 126020 559250
rect 126060 559210 126070 559250
rect 126010 559190 126070 559210
rect 126400 559250 126460 559270
rect 126400 559210 126410 559250
rect 126450 559210 126460 559250
rect 126400 559190 126460 559210
rect 126790 559250 126850 559270
rect 126790 559210 126800 559250
rect 126840 559210 126850 559250
rect 126790 559190 126850 559210
rect 127180 559250 127240 559270
rect 127180 559210 127190 559250
rect 127230 559210 127240 559250
rect 127180 559190 127240 559210
rect 127570 559250 127630 559270
rect 127570 559210 127580 559250
rect 127620 559210 127630 559250
rect 127570 559190 127630 559210
rect 127960 559250 128020 559270
rect 127960 559210 127970 559250
rect 128010 559210 128020 559250
rect 127960 559190 128020 559210
rect 128350 559250 128410 559270
rect 128350 559210 128360 559250
rect 128400 559210 128410 559250
rect 128350 559190 128410 559210
rect 128740 559250 128800 559270
rect 128740 559210 128750 559250
rect 128790 559210 128800 559250
rect 128740 559190 128800 559210
rect 129130 559250 129190 559270
rect 129130 559210 129140 559250
rect 129180 559210 129190 559250
rect 129130 559190 129190 559210
rect 129520 559250 129580 559270
rect 129520 559210 129530 559250
rect 129570 559210 129580 559250
rect 129520 559190 129580 559210
rect 129910 559250 129970 559270
rect 129910 559210 129920 559250
rect 129960 559210 129970 559250
rect 129910 559190 129970 559210
rect 130300 559250 130360 559270
rect 130300 559210 130310 559250
rect 130350 559210 130360 559250
rect 130300 559190 130360 559210
rect 130690 559250 130750 559270
rect 130690 559210 130700 559250
rect 130740 559210 130750 559250
rect 130690 559190 130750 559210
rect 131080 559250 131140 559270
rect 131080 559210 131090 559250
rect 131130 559210 131140 559250
rect 131080 559190 131140 559210
rect 131470 559250 131530 559270
rect 131470 559210 131480 559250
rect 131520 559210 131530 559250
rect 131470 559190 131530 559210
rect 131860 559250 131920 559270
rect 131860 559210 131870 559250
rect 131910 559210 131920 559250
rect 131860 559190 131920 559210
rect 132250 559250 132310 559270
rect 132250 559210 132260 559250
rect 132300 559210 132310 559250
rect 132250 559190 132310 559210
rect 132640 559250 132700 559270
rect 132640 559210 132650 559250
rect 132690 559210 132700 559250
rect 132640 559190 132700 559210
rect 125640 559150 125670 559190
rect 126030 559150 126060 559190
rect 126420 559150 126450 559190
rect 126810 559150 126840 559190
rect 127200 559150 127230 559190
rect 127590 559150 127620 559190
rect 127980 559150 128010 559190
rect 128370 559150 128400 559190
rect 128760 559150 128790 559190
rect 129150 559150 129180 559190
rect 129540 559150 129570 559190
rect 129930 559150 129960 559190
rect 130320 559150 130350 559190
rect 130710 559150 130740 559190
rect 131100 559150 131130 559190
rect 131490 559150 131520 559190
rect 131880 559150 131910 559190
rect 132270 559150 132300 559190
rect 132660 559150 132690 559190
rect 125150 554170 125210 554190
rect 125150 554130 125160 554170
rect 125200 554130 125210 554170
rect 125150 554110 125210 554130
rect 125170 554070 125200 554110
rect 119200 553820 119280 553840
rect 119200 553780 119220 553820
rect 119260 553810 119280 553820
rect 119260 553780 120200 553810
rect 119200 553760 119280 553780
rect 119430 553650 119460 553780
rect 119790 553680 119820 553710
rect 120170 553680 120200 553780
rect 119430 553370 119460 553560
rect 119570 553420 119650 553440
rect 119790 553420 119820 553480
rect 119950 553430 120030 553450
rect 119950 553420 119970 553430
rect 119570 553380 119590 553420
rect 119630 553390 119970 553420
rect 120010 553390 120030 553430
rect 119630 553380 119650 553390
rect 119570 553360 119650 553380
rect 119950 553370 120030 553390
rect 120170 553320 120200 553480
rect 120320 553420 120400 553440
rect 120320 553380 120340 553420
rect 120380 553380 120400 553420
rect 120320 553360 120400 553380
rect 119790 553290 120200 553320
rect 119430 553250 119460 553280
rect 119790 553170 119820 553290
rect 120340 553240 120370 553360
rect 120170 553210 120370 553240
rect 120170 553170 120200 553210
rect 119790 552940 119820 552970
rect 120170 552940 120200 552970
rect 125740 552420 125800 552440
rect 125740 552380 125750 552420
rect 125790 552380 125800 552420
rect 125740 552360 125800 552380
rect 126180 552420 126240 552440
rect 126180 552380 126190 552420
rect 126230 552380 126240 552420
rect 126180 552360 126240 552380
rect 126620 552420 126680 552440
rect 126620 552380 126630 552420
rect 126670 552380 126680 552420
rect 126620 552360 126680 552380
rect 127060 552420 127120 552440
rect 127060 552380 127070 552420
rect 127110 552380 127120 552420
rect 127060 552360 127120 552380
rect 127500 552420 127560 552440
rect 127500 552380 127510 552420
rect 127550 552380 127560 552420
rect 127500 552360 127560 552380
rect 127940 552420 128000 552440
rect 127940 552380 127950 552420
rect 127990 552380 128000 552420
rect 127940 552360 128000 552380
rect 128380 552420 128440 552440
rect 128380 552380 128390 552420
rect 128430 552380 128440 552420
rect 128380 552360 128440 552380
rect 128820 552420 128880 552440
rect 128820 552380 128830 552420
rect 128870 552380 128880 552420
rect 128820 552360 128880 552380
rect 129260 552420 129320 552440
rect 129260 552380 129270 552420
rect 129310 552380 129320 552420
rect 129260 552360 129320 552380
rect 129700 552420 129760 552440
rect 129700 552380 129710 552420
rect 129750 552380 129760 552420
rect 129700 552360 129760 552380
rect 130140 552420 130200 552440
rect 130140 552380 130150 552420
rect 130190 552380 130200 552420
rect 130140 552360 130200 552380
rect 130580 552420 130640 552440
rect 130580 552380 130590 552420
rect 130630 552380 130640 552420
rect 130580 552360 130640 552380
rect 131020 552420 131080 552440
rect 131020 552380 131030 552420
rect 131070 552380 131080 552420
rect 131020 552360 131080 552380
rect 131460 552420 131520 552440
rect 131460 552380 131470 552420
rect 131510 552380 131520 552420
rect 131460 552360 131520 552380
rect 131900 552420 131960 552440
rect 131900 552380 131910 552420
rect 131950 552380 131960 552420
rect 131900 552360 131960 552380
rect 132340 552420 132400 552440
rect 132340 552380 132350 552420
rect 132390 552380 132400 552420
rect 132340 552360 132400 552380
rect 132780 552420 132840 552440
rect 132780 552380 132790 552420
rect 132830 552380 132840 552420
rect 132780 552360 132840 552380
rect 133220 552420 133280 552440
rect 133220 552380 133230 552420
rect 133270 552380 133280 552420
rect 133220 552360 133280 552380
rect 133660 552420 133720 552440
rect 133660 552380 133670 552420
rect 133710 552380 133720 552420
rect 133660 552360 133720 552380
rect 125760 552320 125790 552360
rect 126200 552320 126230 552360
rect 126640 552320 126670 552360
rect 127080 552320 127110 552360
rect 127520 552320 127550 552360
rect 127960 552320 127990 552360
rect 128400 552320 128430 552360
rect 128840 552320 128870 552360
rect 129280 552320 129310 552360
rect 129720 552320 129750 552360
rect 130160 552320 130190 552360
rect 130600 552320 130630 552360
rect 131040 552320 131070 552360
rect 131480 552320 131510 552360
rect 131920 552320 131950 552360
rect 132360 552320 132390 552360
rect 132800 552320 132830 552360
rect 133240 552320 133270 552360
rect 133680 552320 133710 552360
rect 125150 546600 125210 546620
rect 125150 546560 125160 546600
rect 125200 546560 125210 546600
rect 125150 546540 125210 546560
rect 125170 546500 125200 546540
rect 119200 546250 119280 546270
rect 119200 546210 119220 546250
rect 119260 546240 119280 546250
rect 119260 546210 120200 546240
rect 119200 546190 119280 546210
rect 119430 546080 119460 546210
rect 119790 546110 119820 546140
rect 120170 546110 120200 546210
rect 119430 545800 119460 545990
rect 119570 545850 119650 545870
rect 119790 545850 119820 545910
rect 119950 545860 120030 545880
rect 119950 545850 119970 545860
rect 119570 545810 119590 545850
rect 119630 545820 119970 545850
rect 120010 545820 120030 545860
rect 119630 545810 119650 545820
rect 119570 545790 119650 545810
rect 119950 545800 120030 545820
rect 120170 545750 120200 545910
rect 120320 545850 120400 545870
rect 120320 545810 120340 545850
rect 120380 545810 120400 545850
rect 120320 545790 120400 545810
rect 119790 545720 120200 545750
rect 119430 545680 119460 545710
rect 119790 545600 119820 545720
rect 120340 545670 120370 545790
rect 120170 545640 120370 545670
rect 120170 545600 120200 545640
rect 119790 545370 119820 545400
rect 120170 545370 120200 545400
rect 125740 544850 125800 544870
rect 125740 544810 125750 544850
rect 125790 544810 125800 544850
rect 125740 544790 125800 544810
rect 126180 544850 126240 544870
rect 126180 544810 126190 544850
rect 126230 544810 126240 544850
rect 126180 544790 126240 544810
rect 126620 544850 126680 544870
rect 126620 544810 126630 544850
rect 126670 544810 126680 544850
rect 126620 544790 126680 544810
rect 127060 544850 127120 544870
rect 127060 544810 127070 544850
rect 127110 544810 127120 544850
rect 127060 544790 127120 544810
rect 127500 544850 127560 544870
rect 127500 544810 127510 544850
rect 127550 544810 127560 544850
rect 127500 544790 127560 544810
rect 127940 544850 128000 544870
rect 127940 544810 127950 544850
rect 127990 544810 128000 544850
rect 127940 544790 128000 544810
rect 128380 544850 128440 544870
rect 128380 544810 128390 544850
rect 128430 544810 128440 544850
rect 128380 544790 128440 544810
rect 128820 544850 128880 544870
rect 128820 544810 128830 544850
rect 128870 544810 128880 544850
rect 128820 544790 128880 544810
rect 129260 544850 129320 544870
rect 129260 544810 129270 544850
rect 129310 544810 129320 544850
rect 129260 544790 129320 544810
rect 129700 544850 129760 544870
rect 129700 544810 129710 544850
rect 129750 544810 129760 544850
rect 129700 544790 129760 544810
rect 130140 544850 130200 544870
rect 130140 544810 130150 544850
rect 130190 544810 130200 544850
rect 130140 544790 130200 544810
rect 130580 544850 130640 544870
rect 130580 544810 130590 544850
rect 130630 544810 130640 544850
rect 130580 544790 130640 544810
rect 131020 544850 131080 544870
rect 131020 544810 131030 544850
rect 131070 544810 131080 544850
rect 131020 544790 131080 544810
rect 131460 544850 131520 544870
rect 131460 544810 131470 544850
rect 131510 544810 131520 544850
rect 131460 544790 131520 544810
rect 131900 544850 131960 544870
rect 131900 544810 131910 544850
rect 131950 544810 131960 544850
rect 131900 544790 131960 544810
rect 132340 544850 132400 544870
rect 132340 544810 132350 544850
rect 132390 544810 132400 544850
rect 132340 544790 132400 544810
rect 132780 544850 132840 544870
rect 132780 544810 132790 544850
rect 132830 544810 132840 544850
rect 132780 544790 132840 544810
rect 133220 544850 133280 544870
rect 133220 544810 133230 544850
rect 133270 544810 133280 544850
rect 133220 544790 133280 544810
rect 133660 544850 133720 544870
rect 133660 544810 133670 544850
rect 133710 544810 133720 544850
rect 133660 544790 133720 544810
rect 125760 544750 125790 544790
rect 126200 544750 126230 544790
rect 126640 544750 126670 544790
rect 127080 544750 127110 544790
rect 127520 544750 127550 544790
rect 127960 544750 127990 544790
rect 128400 544750 128430 544790
rect 128840 544750 128870 544790
rect 129280 544750 129310 544790
rect 129720 544750 129750 544790
rect 130160 544750 130190 544790
rect 130600 544750 130630 544790
rect 131040 544750 131070 544790
rect 131480 544750 131510 544790
rect 131920 544750 131950 544790
rect 132360 544750 132390 544790
rect 132800 544750 132830 544790
rect 133240 544750 133270 544790
rect 133680 544750 133710 544790
rect 125120 538540 125180 538560
rect 125120 538500 125130 538540
rect 125170 538500 125180 538540
rect 125120 538480 125180 538500
rect 125140 538440 125170 538480
rect 119170 538190 119250 538210
rect 119170 538150 119190 538190
rect 119230 538180 119250 538190
rect 119230 538150 120170 538180
rect 119170 538130 119250 538150
rect 119400 538020 119430 538150
rect 119760 538050 119790 538080
rect 120140 538050 120170 538150
rect 119400 537740 119430 537930
rect 119540 537790 119620 537810
rect 119760 537790 119790 537850
rect 119920 537800 120000 537820
rect 119920 537790 119940 537800
rect 119540 537750 119560 537790
rect 119600 537760 119940 537790
rect 119980 537760 120000 537800
rect 119600 537750 119620 537760
rect 119540 537730 119620 537750
rect 119920 537740 120000 537760
rect 120140 537690 120170 537850
rect 120290 537790 120370 537810
rect 120290 537750 120310 537790
rect 120350 537750 120370 537790
rect 120290 537730 120370 537750
rect 119760 537660 120170 537690
rect 119400 537620 119430 537650
rect 119760 537540 119790 537660
rect 120310 537610 120340 537730
rect 120140 537580 120340 537610
rect 120140 537540 120170 537580
rect 119760 537310 119790 537340
rect 120140 537310 120170 537340
rect 125710 536790 125770 536810
rect 125710 536750 125720 536790
rect 125760 536750 125770 536790
rect 125710 536730 125770 536750
rect 126150 536790 126210 536810
rect 126150 536750 126160 536790
rect 126200 536750 126210 536790
rect 126150 536730 126210 536750
rect 126590 536790 126650 536810
rect 126590 536750 126600 536790
rect 126640 536750 126650 536790
rect 126590 536730 126650 536750
rect 127030 536790 127090 536810
rect 127030 536750 127040 536790
rect 127080 536750 127090 536790
rect 127030 536730 127090 536750
rect 127470 536790 127530 536810
rect 127470 536750 127480 536790
rect 127520 536750 127530 536790
rect 127470 536730 127530 536750
rect 127910 536790 127970 536810
rect 127910 536750 127920 536790
rect 127960 536750 127970 536790
rect 127910 536730 127970 536750
rect 128350 536790 128410 536810
rect 128350 536750 128360 536790
rect 128400 536750 128410 536790
rect 128350 536730 128410 536750
rect 128790 536790 128850 536810
rect 128790 536750 128800 536790
rect 128840 536750 128850 536790
rect 128790 536730 128850 536750
rect 129230 536790 129290 536810
rect 129230 536750 129240 536790
rect 129280 536750 129290 536790
rect 129230 536730 129290 536750
rect 129670 536790 129730 536810
rect 129670 536750 129680 536790
rect 129720 536750 129730 536790
rect 129670 536730 129730 536750
rect 130110 536790 130170 536810
rect 130110 536750 130120 536790
rect 130160 536750 130170 536790
rect 130110 536730 130170 536750
rect 130550 536790 130610 536810
rect 130550 536750 130560 536790
rect 130600 536750 130610 536790
rect 130550 536730 130610 536750
rect 130990 536790 131050 536810
rect 130990 536750 131000 536790
rect 131040 536750 131050 536790
rect 130990 536730 131050 536750
rect 131430 536790 131490 536810
rect 131430 536750 131440 536790
rect 131480 536750 131490 536790
rect 131430 536730 131490 536750
rect 131870 536790 131930 536810
rect 131870 536750 131880 536790
rect 131920 536750 131930 536790
rect 131870 536730 131930 536750
rect 132310 536790 132370 536810
rect 132310 536750 132320 536790
rect 132360 536750 132370 536790
rect 132310 536730 132370 536750
rect 132750 536790 132810 536810
rect 132750 536750 132760 536790
rect 132800 536750 132810 536790
rect 132750 536730 132810 536750
rect 133190 536790 133250 536810
rect 133190 536750 133200 536790
rect 133240 536750 133250 536790
rect 133190 536730 133250 536750
rect 133630 536790 133690 536810
rect 133630 536750 133640 536790
rect 133680 536750 133690 536790
rect 133630 536730 133690 536750
rect 125730 536690 125760 536730
rect 126170 536690 126200 536730
rect 126610 536690 126640 536730
rect 127050 536690 127080 536730
rect 127490 536690 127520 536730
rect 127930 536690 127960 536730
rect 128370 536690 128400 536730
rect 128810 536690 128840 536730
rect 129250 536690 129280 536730
rect 129690 536690 129720 536730
rect 130130 536690 130160 536730
rect 130570 536690 130600 536730
rect 131010 536690 131040 536730
rect 131450 536690 131480 536730
rect 131890 536690 131920 536730
rect 132330 536690 132360 536730
rect 132770 536690 132800 536730
rect 133210 536690 133240 536730
rect 133650 536690 133680 536730
<< polycont >>
rect 124040 642710 124080 642750
rect 124070 636130 124110 636170
rect 124350 630100 124390 630140
rect 124600 623970 124640 624010
rect 125520 619510 125560 619550
rect 125590 618730 125630 618770
rect 125930 618730 125970 618770
rect 126270 618730 126310 618770
rect 126610 618730 126650 618770
rect 126950 618730 126990 618770
rect 127290 618730 127330 618770
rect 127630 618730 127670 618770
rect 127970 618730 128010 618770
rect 128310 618730 128350 618770
rect 128650 618730 128690 618770
rect 128990 618730 129030 618770
rect 129330 618730 129370 618770
rect 129670 618730 129710 618770
rect 130010 618730 130050 618770
rect 130350 618730 130390 618770
rect 130690 618730 130730 618770
rect 131030 618730 131070 618770
rect 131370 618730 131410 618770
rect 131710 618730 131750 618770
rect 125170 612060 125210 612100
rect 125240 611280 125280 611320
rect 125580 611280 125620 611320
rect 125920 611280 125960 611320
rect 126260 611280 126300 611320
rect 126600 611280 126640 611320
rect 126940 611280 126980 611320
rect 127280 611280 127320 611320
rect 127620 611280 127660 611320
rect 127960 611280 128000 611320
rect 128300 611280 128340 611320
rect 128640 611280 128680 611320
rect 128980 611280 129020 611320
rect 129320 611280 129360 611320
rect 129660 611280 129700 611320
rect 130000 611280 130040 611320
rect 130340 611280 130380 611320
rect 130680 611280 130720 611320
rect 131020 611280 131060 611320
rect 131360 611280 131400 611320
rect 125300 606010 125340 606050
rect 125370 605230 125410 605270
rect 125710 605230 125750 605270
rect 126050 605230 126090 605270
rect 126390 605230 126430 605270
rect 126730 605230 126770 605270
rect 127070 605230 127110 605270
rect 127410 605230 127450 605270
rect 127750 605230 127790 605270
rect 128090 605230 128130 605270
rect 128430 605230 128470 605270
rect 128770 605230 128810 605270
rect 129110 605230 129150 605270
rect 129450 605230 129490 605270
rect 129790 605230 129830 605270
rect 130130 605230 130170 605270
rect 130470 605230 130510 605270
rect 130810 605230 130850 605270
rect 131150 605230 131190 605270
rect 131490 605230 131530 605270
rect 125100 599750 125140 599790
rect 125170 598970 125210 599010
rect 125510 598970 125550 599010
rect 125850 598970 125890 599010
rect 126190 598970 126230 599010
rect 126530 598970 126570 599010
rect 126870 598970 126910 599010
rect 127210 598970 127250 599010
rect 127550 598970 127590 599010
rect 127890 598970 127930 599010
rect 128230 598970 128270 599010
rect 128570 598970 128610 599010
rect 128910 598970 128950 599010
rect 129250 598970 129290 599010
rect 129590 598970 129630 599010
rect 129930 598970 129970 599010
rect 130270 598970 130310 599010
rect 130610 598970 130650 599010
rect 130950 598970 130990 599010
rect 131290 598970 131330 599010
rect 119120 593380 119160 593420
rect 119490 592980 119530 593020
rect 119870 592990 119910 593030
rect 120240 592980 120280 593020
rect 125060 592200 125100 592240
rect 125130 591420 125170 591460
rect 125470 591420 125510 591460
rect 125810 591420 125850 591460
rect 126150 591420 126190 591460
rect 126490 591420 126530 591460
rect 126830 591420 126870 591460
rect 127170 591420 127210 591460
rect 127510 591420 127550 591460
rect 127850 591420 127890 591460
rect 128190 591420 128230 591460
rect 128530 591420 128570 591460
rect 128870 591420 128910 591460
rect 129210 591420 129250 591460
rect 129550 591420 129590 591460
rect 129890 591420 129930 591460
rect 130230 591420 130270 591460
rect 130570 591420 130610 591460
rect 130910 591420 130950 591460
rect 131250 591420 131290 591460
rect 119160 583840 119200 583880
rect 119530 583440 119570 583480
rect 119910 583450 119950 583490
rect 120280 583440 120320 583480
rect 125520 583220 125560 583260
rect 125640 582440 125680 582480
rect 126030 582440 126070 582480
rect 126420 582440 126460 582480
rect 126810 582440 126850 582480
rect 127200 582440 127240 582480
rect 127590 582440 127630 582480
rect 127980 582440 128020 582480
rect 128370 582440 128410 582480
rect 128760 582440 128800 582480
rect 129150 582440 129190 582480
rect 129540 582440 129580 582480
rect 129930 582440 129970 582480
rect 130320 582440 130360 582480
rect 130710 582440 130750 582480
rect 131100 582440 131140 582480
rect 131490 582440 131530 582480
rect 131880 582440 131920 582480
rect 132270 582440 132310 582480
rect 132660 582440 132700 582480
rect 119200 574820 119240 574860
rect 119570 574420 119610 574460
rect 119950 574430 119990 574470
rect 120320 574420 120360 574460
rect 125560 574200 125600 574240
rect 125680 573420 125720 573460
rect 126070 573420 126110 573460
rect 126460 573420 126500 573460
rect 126850 573420 126890 573460
rect 127240 573420 127280 573460
rect 127630 573420 127670 573460
rect 128020 573420 128060 573460
rect 128410 573420 128450 573460
rect 128800 573420 128840 573460
rect 129190 573420 129230 573460
rect 129580 573420 129620 573460
rect 129970 573420 130010 573460
rect 130360 573420 130400 573460
rect 130750 573420 130790 573460
rect 131140 573420 131180 573460
rect 131530 573420 131570 573460
rect 131920 573420 131960 573460
rect 132310 573420 132350 573460
rect 132700 573420 132740 573460
rect 119150 567150 119190 567190
rect 119520 566750 119560 566790
rect 119900 566760 119940 566800
rect 120270 566750 120310 566790
rect 125510 566530 125550 566570
rect 125630 565750 125670 565790
rect 126020 565750 126060 565790
rect 126410 565750 126450 565790
rect 126800 565750 126840 565790
rect 127190 565750 127230 565790
rect 127580 565750 127620 565790
rect 127970 565750 128010 565790
rect 128360 565750 128400 565790
rect 128750 565750 128790 565790
rect 129140 565750 129180 565790
rect 129530 565750 129570 565790
rect 129920 565750 129960 565790
rect 130310 565750 130350 565790
rect 130700 565750 130740 565790
rect 131090 565750 131130 565790
rect 131480 565750 131520 565790
rect 131870 565750 131910 565790
rect 132260 565750 132300 565790
rect 132650 565750 132690 565790
rect 119150 560610 119190 560650
rect 119520 560210 119560 560250
rect 119900 560220 119940 560260
rect 120270 560210 120310 560250
rect 125510 559990 125550 560030
rect 125630 559210 125670 559250
rect 126020 559210 126060 559250
rect 126410 559210 126450 559250
rect 126800 559210 126840 559250
rect 127190 559210 127230 559250
rect 127580 559210 127620 559250
rect 127970 559210 128010 559250
rect 128360 559210 128400 559250
rect 128750 559210 128790 559250
rect 129140 559210 129180 559250
rect 129530 559210 129570 559250
rect 129920 559210 129960 559250
rect 130310 559210 130350 559250
rect 130700 559210 130740 559250
rect 131090 559210 131130 559250
rect 131480 559210 131520 559250
rect 131870 559210 131910 559250
rect 132260 559210 132300 559250
rect 132650 559210 132690 559250
rect 125160 554130 125200 554170
rect 119220 553780 119260 553820
rect 119590 553380 119630 553420
rect 119970 553390 120010 553430
rect 120340 553380 120380 553420
rect 125750 552380 125790 552420
rect 126190 552380 126230 552420
rect 126630 552380 126670 552420
rect 127070 552380 127110 552420
rect 127510 552380 127550 552420
rect 127950 552380 127990 552420
rect 128390 552380 128430 552420
rect 128830 552380 128870 552420
rect 129270 552380 129310 552420
rect 129710 552380 129750 552420
rect 130150 552380 130190 552420
rect 130590 552380 130630 552420
rect 131030 552380 131070 552420
rect 131470 552380 131510 552420
rect 131910 552380 131950 552420
rect 132350 552380 132390 552420
rect 132790 552380 132830 552420
rect 133230 552380 133270 552420
rect 133670 552380 133710 552420
rect 125160 546560 125200 546600
rect 119220 546210 119260 546250
rect 119590 545810 119630 545850
rect 119970 545820 120010 545860
rect 120340 545810 120380 545850
rect 125750 544810 125790 544850
rect 126190 544810 126230 544850
rect 126630 544810 126670 544850
rect 127070 544810 127110 544850
rect 127510 544810 127550 544850
rect 127950 544810 127990 544850
rect 128390 544810 128430 544850
rect 128830 544810 128870 544850
rect 129270 544810 129310 544850
rect 129710 544810 129750 544850
rect 130150 544810 130190 544850
rect 130590 544810 130630 544850
rect 131030 544810 131070 544850
rect 131470 544810 131510 544850
rect 131910 544810 131950 544850
rect 132350 544810 132390 544850
rect 132790 544810 132830 544850
rect 133230 544810 133270 544850
rect 133670 544810 133710 544850
rect 125130 538500 125170 538540
rect 119190 538150 119230 538190
rect 119560 537750 119600 537790
rect 119940 537760 119980 537800
rect 120310 537750 120350 537790
rect 125720 536750 125760 536790
rect 126160 536750 126200 536790
rect 126600 536750 126640 536790
rect 127040 536750 127080 536790
rect 127480 536750 127520 536790
rect 127920 536750 127960 536790
rect 128360 536750 128400 536790
rect 128800 536750 128840 536790
rect 129240 536750 129280 536790
rect 129680 536750 129720 536790
rect 130120 536750 130160 536790
rect 130560 536750 130600 536790
rect 131000 536750 131040 536790
rect 131440 536750 131480 536790
rect 131880 536750 131920 536790
rect 132320 536750 132360 536790
rect 132760 536750 132800 536790
rect 133200 536750 133240 536790
rect 133640 536750 133680 536790
<< locali >>
rect 82712 687217 85064 687251
rect 82622 686909 82889 686955
rect 82946 686909 83149 686955
rect 83526 686902 83626 686952
rect 82727 686673 85079 686707
rect 123830 643020 131630 643040
rect 123830 642900 123870 643020
rect 124000 642900 124110 643020
rect 124240 642900 124410 643020
rect 124540 642900 124710 643020
rect 124840 642900 125010 643020
rect 125140 642900 125310 643020
rect 125440 642900 125610 643020
rect 125740 642900 125910 643020
rect 126040 642900 126210 643020
rect 126340 642900 126510 643020
rect 126640 642900 126810 643020
rect 126940 642900 127110 643020
rect 127240 642900 127410 643020
rect 127540 642900 127710 643020
rect 127840 642900 128010 643020
rect 128140 642900 128310 643020
rect 128440 642900 128610 643020
rect 128740 642900 128910 643020
rect 129040 642900 129210 643020
rect 129340 642900 129510 643020
rect 129640 642900 129810 643020
rect 129940 642900 130110 643020
rect 130240 642900 130410 643020
rect 130540 642900 130710 643020
rect 130840 642900 131010 643020
rect 131140 642900 131310 643020
rect 131440 642900 131630 643020
rect 123830 642820 123960 642900
rect 131500 642810 131630 642900
rect 123830 642610 123960 642700
rect 124020 642750 124100 642770
rect 124020 642710 124040 642750
rect 124080 642710 124100 642750
rect 124020 642690 124100 642710
rect 131500 642630 131630 642690
rect 124150 642500 124240 642520
rect 124150 642450 124170 642500
rect 124220 642450 124240 642500
rect 124150 642400 124240 642450
rect 124150 642360 124170 642400
rect 124220 642360 124240 642400
rect 124150 642350 124240 642360
rect 124330 642500 124420 642520
rect 124330 642450 124350 642500
rect 124400 642450 124420 642500
rect 124330 642400 124420 642450
rect 124330 642360 124350 642400
rect 124400 642360 124420 642400
rect 124330 642350 124420 642360
rect 124510 642500 124600 642520
rect 124510 642450 124530 642500
rect 124580 642450 124600 642500
rect 124510 642400 124600 642450
rect 124510 642360 124530 642400
rect 124580 642360 124600 642400
rect 124510 642350 124600 642360
rect 124690 642500 124780 642520
rect 124690 642450 124710 642500
rect 124760 642450 124780 642500
rect 124690 642400 124780 642450
rect 124690 642360 124710 642400
rect 124760 642360 124780 642400
rect 124690 642350 124780 642360
rect 124870 642500 124960 642520
rect 124870 642450 124890 642500
rect 124940 642450 124960 642500
rect 124870 642400 124960 642450
rect 124870 642360 124890 642400
rect 124940 642360 124960 642400
rect 124870 642350 124960 642360
rect 125050 642500 125140 642520
rect 125050 642450 125070 642500
rect 125120 642450 125140 642500
rect 125050 642400 125140 642450
rect 125050 642360 125070 642400
rect 125120 642360 125140 642400
rect 125050 642350 125140 642360
rect 125230 642500 125320 642520
rect 125230 642450 125250 642500
rect 125300 642450 125320 642500
rect 125230 642400 125320 642450
rect 125230 642360 125250 642400
rect 125300 642360 125320 642400
rect 125230 642350 125320 642360
rect 125410 642500 125500 642520
rect 125410 642450 125430 642500
rect 125480 642450 125500 642500
rect 125410 642400 125500 642450
rect 125410 642360 125430 642400
rect 125480 642360 125500 642400
rect 125410 642350 125500 642360
rect 125590 642500 125680 642520
rect 125590 642450 125610 642500
rect 125660 642450 125680 642500
rect 125590 642400 125680 642450
rect 125590 642360 125610 642400
rect 125660 642360 125680 642400
rect 125590 642350 125680 642360
rect 125770 642500 125860 642520
rect 125770 642450 125790 642500
rect 125840 642450 125860 642500
rect 125770 642400 125860 642450
rect 125770 642360 125790 642400
rect 125840 642360 125860 642400
rect 125770 642350 125860 642360
rect 125950 642500 126040 642520
rect 125950 642450 125970 642500
rect 126020 642450 126040 642500
rect 125950 642400 126040 642450
rect 125950 642360 125970 642400
rect 126020 642360 126040 642400
rect 125950 642350 126040 642360
rect 126130 642500 126220 642520
rect 126130 642450 126150 642500
rect 126200 642450 126220 642500
rect 126130 642400 126220 642450
rect 126130 642360 126150 642400
rect 126200 642360 126220 642400
rect 126130 642350 126220 642360
rect 126310 642500 126400 642520
rect 126310 642450 126330 642500
rect 126380 642450 126400 642500
rect 126310 642400 126400 642450
rect 126310 642360 126330 642400
rect 126380 642360 126400 642400
rect 126310 642350 126400 642360
rect 126490 642500 126580 642520
rect 126490 642450 126510 642500
rect 126560 642450 126580 642500
rect 126490 642400 126580 642450
rect 126490 642360 126510 642400
rect 126560 642360 126580 642400
rect 126490 642350 126580 642360
rect 126670 642500 126760 642520
rect 126670 642450 126690 642500
rect 126740 642450 126760 642500
rect 126670 642400 126760 642450
rect 126670 642360 126690 642400
rect 126740 642360 126760 642400
rect 126670 642350 126760 642360
rect 126850 642500 126940 642520
rect 126850 642450 126870 642500
rect 126920 642450 126940 642500
rect 126850 642400 126940 642450
rect 126850 642360 126870 642400
rect 126920 642360 126940 642400
rect 126850 642350 126940 642360
rect 127030 642500 127120 642520
rect 127030 642450 127050 642500
rect 127100 642450 127120 642500
rect 127030 642400 127120 642450
rect 127030 642360 127050 642400
rect 127100 642360 127120 642400
rect 127030 642350 127120 642360
rect 127210 642500 127300 642520
rect 127210 642450 127230 642500
rect 127280 642450 127300 642500
rect 127210 642400 127300 642450
rect 127210 642360 127230 642400
rect 127280 642360 127300 642400
rect 127210 642350 127300 642360
rect 127390 642500 127480 642520
rect 127390 642450 127410 642500
rect 127460 642450 127480 642500
rect 127390 642400 127480 642450
rect 127390 642360 127410 642400
rect 127460 642360 127480 642400
rect 127390 642350 127480 642360
rect 127570 642500 127660 642520
rect 127570 642450 127590 642500
rect 127640 642450 127660 642500
rect 127570 642400 127660 642450
rect 127570 642360 127590 642400
rect 127640 642360 127660 642400
rect 127570 642350 127660 642360
rect 127750 642500 127840 642520
rect 127750 642450 127770 642500
rect 127820 642450 127840 642500
rect 127750 642400 127840 642450
rect 127750 642360 127770 642400
rect 127820 642360 127840 642400
rect 127750 642350 127840 642360
rect 127930 642500 128020 642520
rect 127930 642450 127950 642500
rect 128000 642450 128020 642500
rect 127930 642400 128020 642450
rect 127930 642360 127950 642400
rect 128000 642360 128020 642400
rect 127930 642350 128020 642360
rect 128110 642500 128200 642520
rect 128110 642450 128130 642500
rect 128180 642450 128200 642500
rect 128110 642400 128200 642450
rect 128110 642360 128130 642400
rect 128180 642360 128200 642400
rect 128110 642350 128200 642360
rect 128290 642500 128380 642520
rect 128290 642450 128310 642500
rect 128360 642450 128380 642500
rect 128290 642400 128380 642450
rect 128290 642360 128310 642400
rect 128360 642360 128380 642400
rect 128290 642350 128380 642360
rect 128470 642500 128560 642520
rect 128470 642450 128490 642500
rect 128540 642450 128560 642500
rect 128470 642400 128560 642450
rect 128470 642360 128490 642400
rect 128540 642360 128560 642400
rect 128470 642350 128560 642360
rect 128650 642500 128740 642520
rect 128650 642450 128670 642500
rect 128720 642450 128740 642500
rect 128650 642400 128740 642450
rect 128650 642360 128670 642400
rect 128720 642360 128740 642400
rect 128650 642350 128740 642360
rect 128830 642500 128920 642520
rect 128830 642450 128850 642500
rect 128900 642450 128920 642500
rect 128830 642400 128920 642450
rect 128830 642360 128850 642400
rect 128900 642360 128920 642400
rect 128830 642350 128920 642360
rect 129010 642500 129100 642520
rect 129010 642450 129030 642500
rect 129080 642450 129100 642500
rect 129010 642400 129100 642450
rect 129010 642360 129030 642400
rect 129080 642360 129100 642400
rect 129010 642350 129100 642360
rect 129190 642500 129280 642520
rect 129190 642450 129210 642500
rect 129260 642450 129280 642500
rect 129190 642400 129280 642450
rect 129190 642360 129210 642400
rect 129260 642360 129280 642400
rect 129190 642350 129280 642360
rect 129370 642500 129460 642520
rect 129370 642450 129390 642500
rect 129440 642450 129460 642500
rect 129370 642400 129460 642450
rect 129370 642360 129390 642400
rect 129440 642360 129460 642400
rect 129370 642350 129460 642360
rect 129550 642500 129640 642520
rect 129550 642450 129570 642500
rect 129620 642450 129640 642500
rect 129550 642400 129640 642450
rect 129550 642360 129570 642400
rect 129620 642360 129640 642400
rect 129550 642350 129640 642360
rect 129730 642500 129820 642520
rect 129730 642450 129750 642500
rect 129800 642450 129820 642500
rect 129730 642400 129820 642450
rect 129730 642360 129750 642400
rect 129800 642360 129820 642400
rect 129730 642350 129820 642360
rect 129910 642500 130000 642520
rect 129910 642450 129930 642500
rect 129980 642450 130000 642500
rect 129910 642400 130000 642450
rect 129910 642360 129930 642400
rect 129980 642360 130000 642400
rect 129910 642350 130000 642360
rect 130090 642500 130180 642520
rect 130090 642450 130110 642500
rect 130160 642450 130180 642500
rect 130090 642400 130180 642450
rect 130090 642360 130110 642400
rect 130160 642360 130180 642400
rect 130090 642350 130180 642360
rect 130270 642500 130360 642520
rect 130270 642450 130290 642500
rect 130340 642450 130360 642500
rect 130270 642400 130360 642450
rect 130270 642360 130290 642400
rect 130340 642360 130360 642400
rect 130270 642350 130360 642360
rect 130450 642500 130540 642520
rect 130450 642450 130470 642500
rect 130520 642450 130540 642500
rect 130450 642400 130540 642450
rect 130450 642360 130470 642400
rect 130520 642360 130540 642400
rect 130450 642350 130540 642360
rect 130630 642500 130720 642520
rect 130630 642450 130650 642500
rect 130700 642450 130720 642500
rect 130630 642400 130720 642450
rect 130630 642360 130650 642400
rect 130700 642360 130720 642400
rect 130630 642350 130720 642360
rect 130810 642500 130900 642520
rect 130810 642450 130830 642500
rect 130880 642450 130900 642500
rect 130810 642400 130900 642450
rect 130810 642360 130830 642400
rect 130880 642360 130900 642400
rect 130810 642350 130900 642360
rect 130990 642500 131080 642520
rect 130990 642450 131010 642500
rect 131060 642450 131080 642500
rect 130990 642400 131080 642450
rect 130990 642360 131010 642400
rect 131060 642360 131080 642400
rect 130990 642350 131080 642360
rect 131170 642500 131260 642520
rect 131170 642450 131190 642500
rect 131240 642450 131260 642500
rect 131170 642400 131260 642450
rect 131170 642360 131190 642400
rect 131240 642360 131260 642400
rect 131170 642350 131260 642360
rect 124150 642290 124240 642300
rect 124150 642250 124170 642290
rect 124220 642250 124240 642290
rect 124150 642200 124240 642250
rect 124150 642150 124170 642200
rect 124220 642150 124240 642200
rect 124150 642130 124240 642150
rect 124330 642290 124420 642300
rect 124330 642250 124350 642290
rect 124400 642250 124420 642290
rect 124330 642200 124420 642250
rect 124330 642150 124350 642200
rect 124400 642150 124420 642200
rect 124330 642130 124420 642150
rect 124510 642290 124600 642300
rect 124510 642250 124530 642290
rect 124580 642250 124600 642290
rect 124510 642200 124600 642250
rect 124510 642150 124530 642200
rect 124580 642150 124600 642200
rect 124510 642130 124600 642150
rect 124690 642290 124780 642300
rect 124690 642250 124710 642290
rect 124760 642250 124780 642290
rect 124690 642200 124780 642250
rect 124690 642150 124710 642200
rect 124760 642150 124780 642200
rect 124690 642130 124780 642150
rect 124870 642290 124960 642300
rect 124870 642250 124890 642290
rect 124940 642250 124960 642290
rect 124870 642200 124960 642250
rect 124870 642150 124890 642200
rect 124940 642150 124960 642200
rect 124870 642130 124960 642150
rect 125050 642290 125140 642300
rect 125050 642250 125070 642290
rect 125120 642250 125140 642290
rect 125050 642200 125140 642250
rect 125050 642150 125070 642200
rect 125120 642150 125140 642200
rect 125050 642130 125140 642150
rect 125230 642290 125320 642300
rect 125230 642250 125250 642290
rect 125300 642250 125320 642290
rect 125230 642200 125320 642250
rect 125230 642150 125250 642200
rect 125300 642150 125320 642200
rect 125230 642130 125320 642150
rect 125410 642290 125500 642300
rect 125410 642250 125430 642290
rect 125480 642250 125500 642290
rect 125410 642200 125500 642250
rect 125410 642150 125430 642200
rect 125480 642150 125500 642200
rect 125410 642130 125500 642150
rect 125590 642290 125680 642300
rect 125590 642250 125610 642290
rect 125660 642250 125680 642290
rect 125590 642200 125680 642250
rect 125590 642150 125610 642200
rect 125660 642150 125680 642200
rect 125590 642130 125680 642150
rect 125770 642290 125860 642300
rect 125770 642250 125790 642290
rect 125840 642250 125860 642290
rect 125770 642200 125860 642250
rect 125770 642150 125790 642200
rect 125840 642150 125860 642200
rect 125770 642130 125860 642150
rect 125950 642290 126040 642300
rect 125950 642250 125970 642290
rect 126020 642250 126040 642290
rect 125950 642200 126040 642250
rect 125950 642150 125970 642200
rect 126020 642150 126040 642200
rect 125950 642130 126040 642150
rect 126130 642290 126220 642300
rect 126130 642250 126150 642290
rect 126200 642250 126220 642290
rect 126130 642200 126220 642250
rect 126130 642150 126150 642200
rect 126200 642150 126220 642200
rect 126130 642130 126220 642150
rect 126310 642290 126400 642300
rect 126310 642250 126330 642290
rect 126380 642250 126400 642290
rect 126310 642200 126400 642250
rect 126310 642150 126330 642200
rect 126380 642150 126400 642200
rect 126310 642130 126400 642150
rect 126490 642290 126580 642300
rect 126490 642250 126510 642290
rect 126560 642250 126580 642290
rect 126490 642200 126580 642250
rect 126490 642150 126510 642200
rect 126560 642150 126580 642200
rect 126490 642130 126580 642150
rect 126670 642290 126760 642300
rect 126670 642250 126690 642290
rect 126740 642250 126760 642290
rect 126670 642200 126760 642250
rect 126670 642150 126690 642200
rect 126740 642150 126760 642200
rect 126670 642130 126760 642150
rect 126850 642290 126940 642300
rect 126850 642250 126870 642290
rect 126920 642250 126940 642290
rect 126850 642200 126940 642250
rect 126850 642150 126870 642200
rect 126920 642150 126940 642200
rect 126850 642130 126940 642150
rect 127030 642290 127120 642300
rect 127030 642250 127050 642290
rect 127100 642250 127120 642290
rect 127030 642200 127120 642250
rect 127030 642150 127050 642200
rect 127100 642150 127120 642200
rect 127030 642130 127120 642150
rect 127210 642290 127300 642300
rect 127210 642250 127230 642290
rect 127280 642250 127300 642290
rect 127210 642200 127300 642250
rect 127210 642150 127230 642200
rect 127280 642150 127300 642200
rect 127210 642130 127300 642150
rect 127390 642290 127480 642300
rect 127390 642250 127410 642290
rect 127460 642250 127480 642290
rect 127390 642200 127480 642250
rect 127390 642150 127410 642200
rect 127460 642150 127480 642200
rect 127390 642130 127480 642150
rect 127570 642290 127660 642300
rect 127570 642250 127590 642290
rect 127640 642250 127660 642290
rect 127570 642200 127660 642250
rect 127570 642150 127590 642200
rect 127640 642150 127660 642200
rect 127570 642130 127660 642150
rect 127750 642290 127840 642300
rect 127750 642250 127770 642290
rect 127820 642250 127840 642290
rect 127750 642200 127840 642250
rect 127750 642150 127770 642200
rect 127820 642150 127840 642200
rect 127750 642130 127840 642150
rect 127930 642290 128020 642300
rect 127930 642250 127950 642290
rect 128000 642250 128020 642290
rect 127930 642200 128020 642250
rect 127930 642150 127950 642200
rect 128000 642150 128020 642200
rect 127930 642130 128020 642150
rect 128110 642290 128200 642300
rect 128110 642250 128130 642290
rect 128180 642250 128200 642290
rect 128110 642200 128200 642250
rect 128110 642150 128130 642200
rect 128180 642150 128200 642200
rect 128110 642130 128200 642150
rect 128290 642290 128380 642300
rect 128290 642250 128310 642290
rect 128360 642250 128380 642290
rect 128290 642200 128380 642250
rect 128290 642150 128310 642200
rect 128360 642150 128380 642200
rect 128290 642130 128380 642150
rect 128470 642290 128560 642300
rect 128470 642250 128490 642290
rect 128540 642250 128560 642290
rect 128470 642200 128560 642250
rect 128470 642150 128490 642200
rect 128540 642150 128560 642200
rect 128470 642130 128560 642150
rect 128650 642290 128740 642300
rect 128650 642250 128670 642290
rect 128720 642250 128740 642290
rect 128650 642200 128740 642250
rect 128650 642150 128670 642200
rect 128720 642150 128740 642200
rect 128650 642130 128740 642150
rect 128830 642290 128920 642300
rect 128830 642250 128850 642290
rect 128900 642250 128920 642290
rect 128830 642200 128920 642250
rect 128830 642150 128850 642200
rect 128900 642150 128920 642200
rect 128830 642130 128920 642150
rect 129010 642290 129100 642300
rect 129010 642250 129030 642290
rect 129080 642250 129100 642290
rect 129010 642200 129100 642250
rect 129010 642150 129030 642200
rect 129080 642150 129100 642200
rect 129010 642130 129100 642150
rect 129190 642290 129280 642300
rect 129190 642250 129210 642290
rect 129260 642250 129280 642290
rect 129190 642200 129280 642250
rect 129190 642150 129210 642200
rect 129260 642150 129280 642200
rect 129190 642130 129280 642150
rect 129370 642290 129460 642300
rect 129370 642250 129390 642290
rect 129440 642250 129460 642290
rect 129370 642200 129460 642250
rect 129370 642150 129390 642200
rect 129440 642150 129460 642200
rect 129370 642130 129460 642150
rect 129550 642290 129640 642300
rect 129550 642250 129570 642290
rect 129620 642250 129640 642290
rect 129550 642200 129640 642250
rect 129550 642150 129570 642200
rect 129620 642150 129640 642200
rect 129550 642130 129640 642150
rect 129730 642290 129820 642300
rect 129730 642250 129750 642290
rect 129800 642250 129820 642290
rect 129730 642200 129820 642250
rect 129730 642150 129750 642200
rect 129800 642150 129820 642200
rect 129730 642130 129820 642150
rect 129910 642290 130000 642300
rect 129910 642250 129930 642290
rect 129980 642250 130000 642290
rect 129910 642200 130000 642250
rect 129910 642150 129930 642200
rect 129980 642150 130000 642200
rect 129910 642130 130000 642150
rect 130090 642290 130180 642300
rect 130090 642250 130110 642290
rect 130160 642250 130180 642290
rect 130090 642200 130180 642250
rect 130090 642150 130110 642200
rect 130160 642150 130180 642200
rect 130090 642130 130180 642150
rect 130270 642290 130360 642300
rect 130270 642250 130290 642290
rect 130340 642250 130360 642290
rect 130270 642200 130360 642250
rect 130270 642150 130290 642200
rect 130340 642150 130360 642200
rect 130270 642130 130360 642150
rect 130450 642290 130540 642300
rect 130450 642250 130470 642290
rect 130520 642250 130540 642290
rect 130450 642200 130540 642250
rect 130450 642150 130470 642200
rect 130520 642150 130540 642200
rect 130450 642130 130540 642150
rect 130630 642290 130720 642300
rect 130630 642250 130650 642290
rect 130700 642250 130720 642290
rect 130630 642200 130720 642250
rect 130630 642150 130650 642200
rect 130700 642150 130720 642200
rect 130630 642130 130720 642150
rect 130810 642290 130900 642300
rect 130810 642250 130830 642290
rect 130880 642250 130900 642290
rect 130810 642200 130900 642250
rect 130810 642150 130830 642200
rect 130880 642150 130900 642200
rect 130810 642130 130900 642150
rect 130990 642290 131080 642300
rect 130990 642250 131010 642290
rect 131060 642250 131080 642290
rect 130990 642200 131080 642250
rect 130990 642150 131010 642200
rect 131060 642150 131080 642200
rect 130990 642130 131080 642150
rect 131170 642290 131260 642300
rect 131170 642250 131190 642290
rect 131240 642250 131260 642290
rect 131170 642200 131260 642250
rect 131170 642150 131190 642200
rect 131240 642150 131260 642200
rect 131170 642130 131260 642150
rect 123830 641930 123960 642040
rect 123830 641760 123960 641810
rect 131500 641760 131630 642060
rect 123830 641640 123980 641760
rect 124110 641640 124280 641760
rect 124410 641640 124580 641760
rect 124710 641640 124880 641760
rect 125010 641640 125180 641760
rect 125310 641640 125480 641760
rect 125610 641640 125780 641760
rect 125910 641640 126080 641760
rect 126210 641640 126380 641760
rect 126510 641640 126680 641760
rect 126810 641640 126980 641760
rect 127110 641640 127280 641760
rect 127410 641640 127580 641760
rect 127710 641640 127880 641760
rect 128010 641640 128180 641760
rect 128310 641640 128480 641760
rect 128610 641640 128780 641760
rect 128910 641640 129080 641760
rect 129210 641640 129380 641760
rect 129510 641640 129680 641760
rect 129810 641640 129980 641760
rect 130110 641640 130280 641760
rect 130410 641640 130580 641760
rect 130710 641640 130880 641760
rect 131010 641640 131180 641760
rect 131310 641640 131470 641760
rect 131600 641640 131630 641760
rect 123830 641620 131630 641640
rect 123880 636810 129230 636820
rect 123880 636690 124020 636810
rect 124150 636690 124320 636810
rect 124450 636690 124620 636810
rect 124750 636690 124920 636810
rect 125050 636690 125220 636810
rect 125350 636690 125520 636810
rect 125650 636690 125820 636810
rect 125950 636690 126120 636810
rect 126250 636690 126420 636810
rect 126550 636690 126720 636810
rect 126850 636690 127020 636810
rect 127150 636690 127320 636810
rect 127450 636690 127620 636810
rect 127750 636690 127920 636810
rect 128050 636690 128220 636810
rect 128350 636690 128520 636810
rect 128650 636690 128820 636810
rect 128950 636700 129230 636810
rect 128950 636690 129100 636700
rect 123880 636680 129100 636690
rect 123880 636610 124010 636680
rect 123880 636360 124010 636490
rect 129100 636470 129230 636580
rect 123880 636100 124010 636240
rect 124180 636330 124360 636350
rect 124180 636280 124200 636330
rect 124340 636280 124360 636330
rect 124180 636230 124360 636280
rect 124180 636190 124200 636230
rect 124340 636190 124360 636230
rect 124050 636170 124130 636190
rect 124180 636180 124360 636190
rect 124420 636330 124600 636350
rect 124420 636280 124440 636330
rect 124580 636280 124600 636330
rect 124420 636230 124600 636280
rect 124420 636190 124440 636230
rect 124580 636190 124600 636230
rect 124420 636180 124600 636190
rect 124660 636330 124840 636350
rect 124660 636280 124680 636330
rect 124820 636280 124840 636330
rect 124660 636230 124840 636280
rect 124660 636190 124680 636230
rect 124820 636190 124840 636230
rect 124660 636180 124840 636190
rect 124900 636330 125080 636350
rect 124900 636280 124920 636330
rect 125060 636280 125080 636330
rect 124900 636230 125080 636280
rect 124900 636190 124920 636230
rect 125060 636190 125080 636230
rect 124900 636180 125080 636190
rect 125140 636330 125320 636350
rect 125140 636280 125160 636330
rect 125300 636280 125320 636330
rect 125140 636230 125320 636280
rect 125140 636190 125160 636230
rect 125300 636190 125320 636230
rect 125140 636180 125320 636190
rect 125380 636330 125560 636350
rect 125380 636280 125400 636330
rect 125540 636280 125560 636330
rect 125380 636230 125560 636280
rect 125380 636190 125400 636230
rect 125540 636190 125560 636230
rect 125380 636180 125560 636190
rect 125620 636330 125800 636350
rect 125620 636280 125640 636330
rect 125780 636280 125800 636330
rect 125620 636230 125800 636280
rect 125620 636190 125640 636230
rect 125780 636190 125800 636230
rect 125620 636180 125800 636190
rect 125860 636330 126040 636350
rect 125860 636280 125880 636330
rect 126020 636280 126040 636330
rect 125860 636230 126040 636280
rect 125860 636190 125880 636230
rect 126020 636190 126040 636230
rect 125860 636180 126040 636190
rect 126100 636330 126280 636350
rect 126100 636280 126120 636330
rect 126260 636280 126280 636330
rect 126100 636230 126280 636280
rect 126100 636190 126120 636230
rect 126260 636190 126280 636230
rect 126100 636180 126280 636190
rect 126340 636330 126520 636350
rect 126340 636280 126360 636330
rect 126500 636280 126520 636330
rect 126340 636230 126520 636280
rect 126340 636190 126360 636230
rect 126500 636190 126520 636230
rect 126340 636180 126520 636190
rect 126580 636330 126760 636350
rect 126580 636280 126600 636330
rect 126740 636280 126760 636330
rect 126580 636230 126760 636280
rect 126580 636190 126600 636230
rect 126740 636190 126760 636230
rect 126580 636180 126760 636190
rect 126820 636330 127000 636350
rect 126820 636280 126840 636330
rect 126980 636280 127000 636330
rect 126820 636230 127000 636280
rect 126820 636190 126840 636230
rect 126980 636190 127000 636230
rect 126820 636180 127000 636190
rect 127060 636330 127240 636350
rect 127060 636280 127080 636330
rect 127220 636280 127240 636330
rect 127060 636230 127240 636280
rect 127060 636190 127080 636230
rect 127220 636190 127240 636230
rect 127060 636180 127240 636190
rect 127300 636330 127480 636350
rect 127300 636280 127320 636330
rect 127460 636280 127480 636330
rect 127300 636230 127480 636280
rect 127300 636190 127320 636230
rect 127460 636190 127480 636230
rect 127300 636180 127480 636190
rect 127540 636330 127720 636350
rect 127540 636280 127560 636330
rect 127700 636280 127720 636330
rect 127540 636230 127720 636280
rect 127540 636190 127560 636230
rect 127700 636190 127720 636230
rect 127540 636180 127720 636190
rect 127780 636330 127960 636350
rect 127780 636280 127800 636330
rect 127940 636280 127960 636330
rect 127780 636230 127960 636280
rect 127780 636190 127800 636230
rect 127940 636190 127960 636230
rect 127780 636180 127960 636190
rect 128020 636330 128200 636350
rect 128020 636280 128040 636330
rect 128180 636280 128200 636330
rect 128020 636230 128200 636280
rect 128020 636190 128040 636230
rect 128180 636190 128200 636230
rect 128020 636180 128200 636190
rect 128260 636330 128440 636350
rect 128260 636280 128280 636330
rect 128420 636280 128440 636330
rect 128260 636230 128440 636280
rect 128260 636190 128280 636230
rect 128420 636190 128440 636230
rect 128260 636180 128440 636190
rect 128500 636330 128680 636350
rect 128500 636280 128520 636330
rect 128660 636280 128680 636330
rect 128500 636230 128680 636280
rect 128500 636190 128520 636230
rect 128660 636190 128680 636230
rect 128500 636180 128680 636190
rect 128740 636330 128920 636350
rect 128740 636280 128760 636330
rect 128900 636280 128920 636330
rect 128740 636230 128920 636280
rect 128740 636190 128760 636230
rect 128900 636190 128920 636230
rect 128740 636180 128920 636190
rect 124050 636130 124070 636170
rect 124110 636130 124130 636170
rect 124050 636110 124130 636130
rect 124180 636120 124360 636130
rect 123880 635820 124010 635980
rect 124180 636080 124200 636120
rect 124340 636080 124360 636120
rect 124180 636030 124360 636080
rect 124180 635980 124200 636030
rect 124340 635980 124360 636030
rect 124180 635960 124360 635980
rect 124420 636120 124600 636130
rect 124420 636080 124440 636120
rect 124580 636080 124600 636120
rect 124420 636030 124600 636080
rect 124420 635980 124440 636030
rect 124580 635980 124600 636030
rect 124420 635960 124600 635980
rect 124660 636120 124840 636130
rect 124660 636080 124680 636120
rect 124820 636080 124840 636120
rect 124660 636030 124840 636080
rect 124660 635980 124680 636030
rect 124820 635980 124840 636030
rect 124660 635960 124840 635980
rect 124900 636120 125080 636130
rect 124900 636080 124920 636120
rect 125060 636080 125080 636120
rect 124900 636030 125080 636080
rect 124900 635980 124920 636030
rect 125060 635980 125080 636030
rect 124900 635960 125080 635980
rect 125140 636120 125320 636130
rect 125140 636080 125160 636120
rect 125300 636080 125320 636120
rect 125140 636030 125320 636080
rect 125140 635980 125160 636030
rect 125300 635980 125320 636030
rect 125140 635960 125320 635980
rect 125380 636120 125560 636130
rect 125380 636080 125400 636120
rect 125540 636080 125560 636120
rect 125380 636030 125560 636080
rect 125380 635980 125400 636030
rect 125540 635980 125560 636030
rect 125380 635960 125560 635980
rect 125620 636120 125800 636130
rect 125620 636080 125640 636120
rect 125780 636080 125800 636120
rect 125620 636030 125800 636080
rect 125620 635980 125640 636030
rect 125780 635980 125800 636030
rect 125620 635960 125800 635980
rect 125860 636120 126040 636130
rect 125860 636080 125880 636120
rect 126020 636080 126040 636120
rect 125860 636030 126040 636080
rect 125860 635980 125880 636030
rect 126020 635980 126040 636030
rect 125860 635960 126040 635980
rect 126100 636120 126280 636130
rect 126100 636080 126120 636120
rect 126260 636080 126280 636120
rect 126100 636030 126280 636080
rect 126100 635980 126120 636030
rect 126260 635980 126280 636030
rect 126100 635960 126280 635980
rect 126340 636120 126520 636130
rect 126340 636080 126360 636120
rect 126500 636080 126520 636120
rect 126340 636030 126520 636080
rect 126340 635980 126360 636030
rect 126500 635980 126520 636030
rect 126340 635960 126520 635980
rect 126580 636120 126760 636130
rect 126580 636080 126600 636120
rect 126740 636080 126760 636120
rect 126580 636030 126760 636080
rect 126580 635980 126600 636030
rect 126740 635980 126760 636030
rect 126580 635960 126760 635980
rect 126820 636120 127000 636130
rect 126820 636080 126840 636120
rect 126980 636080 127000 636120
rect 126820 636030 127000 636080
rect 126820 635980 126840 636030
rect 126980 635980 127000 636030
rect 126820 635960 127000 635980
rect 127060 636120 127240 636130
rect 127060 636080 127080 636120
rect 127220 636080 127240 636120
rect 127060 636030 127240 636080
rect 127060 635980 127080 636030
rect 127220 635980 127240 636030
rect 127060 635960 127240 635980
rect 127300 636120 127480 636130
rect 127300 636080 127320 636120
rect 127460 636080 127480 636120
rect 127300 636030 127480 636080
rect 127300 635980 127320 636030
rect 127460 635980 127480 636030
rect 127300 635960 127480 635980
rect 127540 636120 127720 636130
rect 127540 636080 127560 636120
rect 127700 636080 127720 636120
rect 127540 636030 127720 636080
rect 127540 635980 127560 636030
rect 127700 635980 127720 636030
rect 127540 635960 127720 635980
rect 127780 636120 127960 636130
rect 127780 636080 127800 636120
rect 127940 636080 127960 636120
rect 127780 636030 127960 636080
rect 127780 635980 127800 636030
rect 127940 635980 127960 636030
rect 127780 635960 127960 635980
rect 128020 636120 128200 636130
rect 128020 636080 128040 636120
rect 128180 636080 128200 636120
rect 128020 636030 128200 636080
rect 128020 635980 128040 636030
rect 128180 635980 128200 636030
rect 128020 635960 128200 635980
rect 128260 636120 128440 636130
rect 128260 636080 128280 636120
rect 128420 636080 128440 636120
rect 128260 636030 128440 636080
rect 128260 635980 128280 636030
rect 128420 635980 128440 636030
rect 128260 635960 128440 635980
rect 128500 636120 128680 636130
rect 128500 636080 128520 636120
rect 128660 636080 128680 636120
rect 128500 636030 128680 636080
rect 128500 635980 128520 636030
rect 128660 635980 128680 636030
rect 128500 635960 128680 635980
rect 128740 636120 128920 636130
rect 128740 636080 128760 636120
rect 128900 636080 128920 636120
rect 128740 636030 128920 636080
rect 128740 635980 128760 636030
rect 128900 635980 128920 636030
rect 128740 635960 128920 635980
rect 123880 635660 124010 635700
rect 129100 635820 129230 635900
rect 129100 635660 129230 635700
rect 123880 635540 124020 635660
rect 124150 635540 124320 635660
rect 124450 635540 124620 635660
rect 124750 635540 124920 635660
rect 125050 635540 125220 635660
rect 125350 635540 125520 635660
rect 125650 635540 125820 635660
rect 125950 635540 126120 635660
rect 126250 635540 126420 635660
rect 126550 635540 126720 635660
rect 126850 635540 127020 635660
rect 127150 635540 127320 635660
rect 127450 635540 127620 635660
rect 127750 635540 127920 635660
rect 128050 635540 128220 635660
rect 128350 635540 128520 635660
rect 128650 635540 128820 635660
rect 128950 635540 129230 635660
rect 124240 632740 124640 632760
rect 124240 632690 124260 632740
rect 124620 632690 124640 632740
rect 124240 632640 124640 632690
rect 124240 632600 124260 632640
rect 124620 632600 124640 632640
rect 124240 632590 124640 632600
rect 124240 632530 124640 632540
rect 124240 632490 124260 632530
rect 124620 632490 124640 632530
rect 124240 632440 124640 632490
rect 124240 632390 124260 632440
rect 124620 632390 124640 632440
rect 124240 632370 124640 632390
rect 124160 630720 129300 630740
rect 124160 630600 124390 630720
rect 124520 630600 124690 630720
rect 124820 630600 124990 630720
rect 125120 630600 125290 630720
rect 125420 630600 125590 630720
rect 125720 630600 125890 630720
rect 126020 630600 126190 630720
rect 126320 630600 126490 630720
rect 126620 630600 126790 630720
rect 126920 630600 127090 630720
rect 127220 630600 127390 630720
rect 127520 630600 127690 630720
rect 127820 630600 127990 630720
rect 128120 630600 128290 630720
rect 128420 630600 128590 630720
rect 128720 630600 128890 630720
rect 129020 630620 129300 630720
rect 129020 630600 129170 630620
rect 124160 630590 129170 630600
rect 124160 630240 124290 630470
rect 129170 630410 129300 630500
rect 124450 630300 124850 630320
rect 124450 630250 124470 630300
rect 124830 630250 124850 630300
rect 124450 630200 124850 630250
rect 124450 630160 124470 630200
rect 124830 630160 124850 630200
rect 124160 629860 124290 630120
rect 124330 630140 124410 630160
rect 124450 630150 124850 630160
rect 124910 630300 125310 630320
rect 124910 630250 124930 630300
rect 125290 630250 125310 630300
rect 124910 630200 125310 630250
rect 124910 630160 124930 630200
rect 125290 630160 125310 630200
rect 124910 630150 125310 630160
rect 125370 630300 125770 630320
rect 125370 630250 125390 630300
rect 125750 630250 125770 630300
rect 125370 630200 125770 630250
rect 125370 630160 125390 630200
rect 125750 630160 125770 630200
rect 125370 630150 125770 630160
rect 125830 630300 126230 630320
rect 125830 630250 125850 630300
rect 126210 630250 126230 630300
rect 125830 630200 126230 630250
rect 125830 630160 125850 630200
rect 126210 630160 126230 630200
rect 125830 630150 126230 630160
rect 126290 630300 126690 630320
rect 126290 630250 126310 630300
rect 126670 630250 126690 630300
rect 126290 630200 126690 630250
rect 126290 630160 126310 630200
rect 126670 630160 126690 630200
rect 126290 630150 126690 630160
rect 126750 630300 127150 630320
rect 126750 630250 126770 630300
rect 127130 630250 127150 630300
rect 126750 630200 127150 630250
rect 126750 630160 126770 630200
rect 127130 630160 127150 630200
rect 126750 630150 127150 630160
rect 127210 630300 127610 630320
rect 127210 630250 127230 630300
rect 127590 630250 127610 630300
rect 127210 630200 127610 630250
rect 127210 630160 127230 630200
rect 127590 630160 127610 630200
rect 127210 630150 127610 630160
rect 127670 630300 128070 630320
rect 127670 630250 127690 630300
rect 128050 630250 128070 630300
rect 127670 630200 128070 630250
rect 127670 630160 127690 630200
rect 128050 630160 128070 630200
rect 127670 630150 128070 630160
rect 128130 630300 128530 630320
rect 128130 630250 128150 630300
rect 128510 630250 128530 630300
rect 128130 630200 128530 630250
rect 128130 630160 128150 630200
rect 128510 630160 128530 630200
rect 128130 630150 128530 630160
rect 128590 630300 128990 630320
rect 128590 630250 128610 630300
rect 128970 630250 128990 630300
rect 128590 630200 128990 630250
rect 128590 630160 128610 630200
rect 128970 630160 128990 630200
rect 128590 630150 128990 630160
rect 124330 630100 124350 630140
rect 124390 630100 124410 630140
rect 124330 630080 124410 630100
rect 124450 630090 124850 630100
rect 124450 630050 124470 630090
rect 124830 630050 124850 630090
rect 124450 630000 124850 630050
rect 124450 629950 124470 630000
rect 124830 629950 124850 630000
rect 124450 629930 124850 629950
rect 124910 630090 125310 630100
rect 124910 630050 124930 630090
rect 125290 630050 125310 630090
rect 124910 630000 125310 630050
rect 124910 629950 124930 630000
rect 125290 629950 125310 630000
rect 124910 629930 125310 629950
rect 125370 630090 125770 630100
rect 125370 630050 125390 630090
rect 125750 630050 125770 630090
rect 125370 630000 125770 630050
rect 125370 629950 125390 630000
rect 125750 629950 125770 630000
rect 125370 629930 125770 629950
rect 125830 630090 126230 630100
rect 125830 630050 125850 630090
rect 126210 630050 126230 630090
rect 125830 630000 126230 630050
rect 125830 629950 125850 630000
rect 126210 629950 126230 630000
rect 125830 629930 126230 629950
rect 126290 630090 126690 630100
rect 126290 630050 126310 630090
rect 126670 630050 126690 630090
rect 126290 630000 126690 630050
rect 126290 629950 126310 630000
rect 126670 629950 126690 630000
rect 126290 629930 126690 629950
rect 126750 630090 127150 630100
rect 126750 630050 126770 630090
rect 127130 630050 127150 630090
rect 126750 630000 127150 630050
rect 126750 629950 126770 630000
rect 127130 629950 127150 630000
rect 126750 629930 127150 629950
rect 127210 630090 127610 630100
rect 127210 630050 127230 630090
rect 127590 630050 127610 630090
rect 127210 630000 127610 630050
rect 127210 629950 127230 630000
rect 127590 629950 127610 630000
rect 127210 629930 127610 629950
rect 127670 630090 128070 630100
rect 127670 630050 127690 630090
rect 128050 630050 128070 630090
rect 127670 630000 128070 630050
rect 127670 629950 127690 630000
rect 128050 629950 128070 630000
rect 127670 629930 128070 629950
rect 128130 630090 128530 630100
rect 128130 630050 128150 630090
rect 128510 630050 128530 630090
rect 128130 630000 128530 630050
rect 128130 629950 128150 630000
rect 128510 629950 128530 630000
rect 128130 629930 128530 629950
rect 128590 630090 128990 630100
rect 128590 630050 128610 630090
rect 128970 630050 128990 630090
rect 128590 630000 128990 630050
rect 128590 629950 128610 630000
rect 128970 629950 128990 630000
rect 128590 629930 128990 629950
rect 124160 629690 124290 629740
rect 129170 629690 129300 629840
rect 124160 629680 129300 629690
rect 124160 629560 124390 629680
rect 124520 629560 124690 629680
rect 124820 629560 124990 629680
rect 125120 629560 125290 629680
rect 125420 629560 125590 629680
rect 125720 629560 125890 629680
rect 126020 629560 126190 629680
rect 126320 629560 126490 629680
rect 126620 629560 126790 629680
rect 126920 629560 127090 629680
rect 127220 629560 127390 629680
rect 127520 629560 127690 629680
rect 127820 629560 127990 629680
rect 128120 629560 128290 629680
rect 128420 629560 128590 629680
rect 128720 629560 128890 629680
rect 129020 629560 129300 629680
rect 124160 629540 129300 629560
rect 124220 625070 124820 625090
rect 124220 625020 124240 625070
rect 124800 625020 124820 625070
rect 124220 624970 124820 625020
rect 124220 624930 124240 624970
rect 124800 624930 124820 624970
rect 124220 624920 124820 624930
rect 124220 624860 124820 624870
rect 124220 624820 124240 624860
rect 124800 624820 124820 624860
rect 124220 624770 124820 624820
rect 124220 624720 124240 624770
rect 124800 624720 124820 624770
rect 124220 624700 124820 624720
rect 124410 624210 128950 624220
rect 124410 624140 124630 624210
rect 124540 624090 124630 624140
rect 124760 624090 124930 624210
rect 125060 624090 125230 624210
rect 125360 624090 125530 624210
rect 125660 624090 125830 624210
rect 125960 624090 126130 624210
rect 126260 624090 126430 624210
rect 126560 624090 126730 624210
rect 126860 624090 127030 624210
rect 127160 624090 127330 624210
rect 127460 624090 127630 624210
rect 127760 624090 127930 624210
rect 128060 624090 128230 624210
rect 128360 624090 128530 624210
rect 128660 624150 128950 624210
rect 128660 624090 128820 624150
rect 124540 624070 128820 624090
rect 124410 623840 124540 624020
rect 124580 624010 124660 624030
rect 124580 623970 124600 624010
rect 124640 623970 124660 624010
rect 124580 623950 124660 623970
rect 128820 623890 128950 624030
rect 124410 623540 124540 623720
rect 124780 623780 125380 623800
rect 124780 623730 124800 623780
rect 125360 623730 125380 623780
rect 124780 623680 125380 623730
rect 124780 623640 124800 623680
rect 125360 623640 125380 623680
rect 124780 623630 125380 623640
rect 125440 623780 126040 623800
rect 125440 623730 125460 623780
rect 126020 623730 126040 623780
rect 125440 623680 126040 623730
rect 125440 623640 125460 623680
rect 126020 623640 126040 623680
rect 125440 623630 126040 623640
rect 126100 623780 126700 623800
rect 126100 623730 126120 623780
rect 126680 623730 126700 623780
rect 126100 623680 126700 623730
rect 126100 623640 126120 623680
rect 126680 623640 126700 623680
rect 126100 623630 126700 623640
rect 126760 623780 127360 623800
rect 126760 623730 126780 623780
rect 127340 623730 127360 623780
rect 126760 623680 127360 623730
rect 126760 623640 126780 623680
rect 127340 623640 127360 623680
rect 126760 623630 127360 623640
rect 127420 623780 128020 623800
rect 127420 623730 127440 623780
rect 128000 623730 128020 623780
rect 127420 623680 128020 623730
rect 127420 623640 127440 623680
rect 128000 623640 128020 623680
rect 127420 623630 128020 623640
rect 128080 623780 128680 623800
rect 128080 623730 128100 623780
rect 128660 623730 128680 623780
rect 128080 623680 128680 623730
rect 128080 623640 128100 623680
rect 128660 623640 128680 623680
rect 128080 623630 128680 623640
rect 124410 623240 124540 623420
rect 124780 623570 125380 623580
rect 124780 623530 124800 623570
rect 125360 623530 125380 623570
rect 124780 623480 125380 623530
rect 124780 623430 124800 623480
rect 125360 623430 125380 623480
rect 124780 623410 125380 623430
rect 125440 623570 126040 623580
rect 125440 623530 125460 623570
rect 126020 623530 126040 623570
rect 125440 623480 126040 623530
rect 125440 623430 125460 623480
rect 126020 623430 126040 623480
rect 125440 623410 126040 623430
rect 126100 623570 126700 623580
rect 126100 623530 126120 623570
rect 126680 623530 126700 623570
rect 126100 623480 126700 623530
rect 126100 623430 126120 623480
rect 126680 623430 126700 623480
rect 126100 623410 126700 623430
rect 126760 623570 127360 623580
rect 126760 623530 126780 623570
rect 127340 623530 127360 623570
rect 126760 623480 127360 623530
rect 126760 623430 126780 623480
rect 127340 623430 127360 623480
rect 126760 623410 127360 623430
rect 127420 623570 128020 623580
rect 127420 623530 127440 623570
rect 128000 623530 128020 623570
rect 127420 623480 128020 623530
rect 127420 623430 127440 623480
rect 128000 623430 128020 623480
rect 127420 623410 128020 623430
rect 128080 623570 128680 623580
rect 128080 623530 128100 623570
rect 128660 623530 128680 623570
rect 128080 623480 128680 623530
rect 128080 623430 128100 623480
rect 128660 623430 128680 623480
rect 128080 623410 128680 623430
rect 128820 623170 128950 623320
rect 124540 623160 128950 623170
rect 124540 623120 124670 623160
rect 124410 623040 124670 623120
rect 124800 623040 124970 623160
rect 125100 623040 125270 623160
rect 125400 623040 125570 623160
rect 125700 623040 125870 623160
rect 126000 623040 126170 623160
rect 126300 623040 126470 623160
rect 126600 623040 126770 623160
rect 126900 623040 127070 623160
rect 127200 623040 127370 623160
rect 127500 623040 127670 623160
rect 127800 623040 127970 623160
rect 128100 623040 128270 623160
rect 128400 623040 128570 623160
rect 128700 623040 128950 623160
rect 124410 623020 128950 623040
rect 125510 619550 125570 619570
rect 125510 619510 125520 619550
rect 125560 619510 125570 619550
rect 125510 619490 125570 619510
rect 125350 619350 125410 619370
rect 125350 619310 125360 619350
rect 125400 619310 125410 619350
rect 125350 619290 125410 619310
rect 125450 619350 125530 619370
rect 125450 619310 125470 619350
rect 125510 619310 125530 619350
rect 125450 619300 125530 619310
rect 125570 619350 125630 619370
rect 125570 619310 125580 619350
rect 125620 619310 125630 619350
rect 125570 619290 125630 619310
rect 125040 618860 125230 618990
rect 125370 618860 125730 618990
rect 125870 618860 126230 618990
rect 126370 618860 126730 618990
rect 126870 618860 127230 618990
rect 127370 618860 127730 618990
rect 127870 618860 128230 618990
rect 128370 618860 128730 618990
rect 128870 618860 129230 618990
rect 129370 618860 129730 618990
rect 129870 618860 130230 618990
rect 130370 618860 130730 618990
rect 130870 618860 131230 618990
rect 131370 618860 131730 618990
rect 131870 618860 132080 618990
rect 125040 618770 125180 618860
rect 131940 618810 132080 618860
rect 132070 618790 132080 618810
rect 125580 618770 125640 618790
rect 125580 618730 125590 618770
rect 125630 618730 125640 618770
rect 125580 618710 125640 618730
rect 125920 618770 125980 618790
rect 125920 618730 125930 618770
rect 125970 618730 125980 618770
rect 125920 618710 125980 618730
rect 126260 618770 126320 618790
rect 126260 618730 126270 618770
rect 126310 618730 126320 618770
rect 126260 618710 126320 618730
rect 126600 618770 126660 618790
rect 126600 618730 126610 618770
rect 126650 618730 126660 618770
rect 126600 618710 126660 618730
rect 126940 618770 127000 618790
rect 126940 618730 126950 618770
rect 126990 618730 127000 618770
rect 126940 618710 127000 618730
rect 127280 618770 127340 618790
rect 127280 618730 127290 618770
rect 127330 618730 127340 618770
rect 127280 618710 127340 618730
rect 127620 618770 127680 618790
rect 127620 618730 127630 618770
rect 127670 618730 127680 618770
rect 127620 618710 127680 618730
rect 127960 618770 128020 618790
rect 127960 618730 127970 618770
rect 128010 618730 128020 618770
rect 127960 618710 128020 618730
rect 128300 618770 128360 618790
rect 128300 618730 128310 618770
rect 128350 618730 128360 618770
rect 128300 618710 128360 618730
rect 128640 618770 128700 618790
rect 128640 618730 128650 618770
rect 128690 618730 128700 618770
rect 128640 618710 128700 618730
rect 128980 618770 129040 618790
rect 128980 618730 128990 618770
rect 129030 618730 129040 618770
rect 128980 618710 129040 618730
rect 129320 618770 129380 618790
rect 129320 618730 129330 618770
rect 129370 618730 129380 618770
rect 129320 618710 129380 618730
rect 129660 618770 129720 618790
rect 129660 618730 129670 618770
rect 129710 618730 129720 618770
rect 129660 618710 129720 618730
rect 130000 618770 130060 618790
rect 130000 618730 130010 618770
rect 130050 618730 130060 618770
rect 130000 618710 130060 618730
rect 130340 618770 130400 618790
rect 130340 618730 130350 618770
rect 130390 618730 130400 618770
rect 130340 618710 130400 618730
rect 130680 618770 130740 618790
rect 130680 618730 130690 618770
rect 130730 618730 130740 618770
rect 130680 618710 130740 618730
rect 131020 618770 131080 618790
rect 131020 618730 131030 618770
rect 131070 618730 131080 618770
rect 131020 618710 131080 618730
rect 131360 618770 131420 618790
rect 131360 618730 131370 618770
rect 131410 618730 131420 618770
rect 131360 618710 131420 618730
rect 131700 618770 131760 618790
rect 131700 618730 131710 618770
rect 131750 618730 131760 618770
rect 131700 618710 131760 618730
rect 125040 618410 125180 618640
rect 125420 618570 125480 618590
rect 125420 618530 125430 618570
rect 125470 618530 125480 618570
rect 125420 618510 125480 618530
rect 125520 618570 125600 618590
rect 125520 618530 125540 618570
rect 125580 618530 125600 618570
rect 125520 618520 125600 618530
rect 125640 618570 125700 618590
rect 125640 618530 125650 618570
rect 125690 618530 125700 618570
rect 125640 618510 125700 618530
rect 125760 618570 125820 618590
rect 125760 618530 125770 618570
rect 125810 618530 125820 618570
rect 125760 618510 125820 618530
rect 125860 618570 125940 618590
rect 125860 618530 125880 618570
rect 125920 618530 125940 618570
rect 125860 618520 125940 618530
rect 125980 618570 126040 618590
rect 125980 618530 125990 618570
rect 126030 618530 126040 618570
rect 125980 618510 126040 618530
rect 126100 618570 126160 618590
rect 126100 618530 126110 618570
rect 126150 618530 126160 618570
rect 126100 618510 126160 618530
rect 126200 618570 126280 618590
rect 126200 618530 126220 618570
rect 126260 618530 126280 618570
rect 126200 618520 126280 618530
rect 126320 618570 126380 618590
rect 126320 618530 126330 618570
rect 126370 618530 126380 618570
rect 126320 618510 126380 618530
rect 126440 618570 126500 618590
rect 126440 618530 126450 618570
rect 126490 618530 126500 618570
rect 126440 618510 126500 618530
rect 126540 618570 126620 618590
rect 126540 618530 126560 618570
rect 126600 618530 126620 618570
rect 126540 618520 126620 618530
rect 126660 618570 126720 618590
rect 126660 618530 126670 618570
rect 126710 618530 126720 618570
rect 126660 618510 126720 618530
rect 126780 618570 126840 618590
rect 126780 618530 126790 618570
rect 126830 618530 126840 618570
rect 126780 618510 126840 618530
rect 126880 618570 126960 618590
rect 126880 618530 126900 618570
rect 126940 618530 126960 618570
rect 126880 618520 126960 618530
rect 127000 618570 127060 618590
rect 127000 618530 127010 618570
rect 127050 618530 127060 618570
rect 127000 618510 127060 618530
rect 127120 618570 127180 618590
rect 127120 618530 127130 618570
rect 127170 618530 127180 618570
rect 127120 618510 127180 618530
rect 127220 618570 127300 618590
rect 127220 618530 127240 618570
rect 127280 618530 127300 618570
rect 127220 618520 127300 618530
rect 127340 618570 127400 618590
rect 127340 618530 127350 618570
rect 127390 618530 127400 618570
rect 127340 618510 127400 618530
rect 127460 618570 127520 618590
rect 127460 618530 127470 618570
rect 127510 618530 127520 618570
rect 127460 618510 127520 618530
rect 127560 618570 127640 618590
rect 127560 618530 127580 618570
rect 127620 618530 127640 618570
rect 127560 618520 127640 618530
rect 127680 618570 127740 618590
rect 127680 618530 127690 618570
rect 127730 618530 127740 618570
rect 127680 618510 127740 618530
rect 127800 618570 127860 618590
rect 127800 618530 127810 618570
rect 127850 618530 127860 618570
rect 127800 618510 127860 618530
rect 127900 618570 127980 618590
rect 127900 618530 127920 618570
rect 127960 618530 127980 618570
rect 127900 618520 127980 618530
rect 128020 618570 128080 618590
rect 128020 618530 128030 618570
rect 128070 618530 128080 618570
rect 128020 618510 128080 618530
rect 128140 618570 128200 618590
rect 128140 618530 128150 618570
rect 128190 618530 128200 618570
rect 128140 618510 128200 618530
rect 128240 618570 128320 618590
rect 128240 618530 128260 618570
rect 128300 618530 128320 618570
rect 128240 618520 128320 618530
rect 128360 618570 128420 618590
rect 128360 618530 128370 618570
rect 128410 618530 128420 618570
rect 128360 618510 128420 618530
rect 128480 618570 128540 618590
rect 128480 618530 128490 618570
rect 128530 618530 128540 618570
rect 128480 618510 128540 618530
rect 128580 618570 128660 618590
rect 128580 618530 128600 618570
rect 128640 618530 128660 618570
rect 128580 618520 128660 618530
rect 128700 618570 128760 618590
rect 128700 618530 128710 618570
rect 128750 618530 128760 618570
rect 128700 618510 128760 618530
rect 128820 618570 128880 618590
rect 128820 618530 128830 618570
rect 128870 618530 128880 618570
rect 128820 618510 128880 618530
rect 128920 618570 129000 618590
rect 128920 618530 128940 618570
rect 128980 618530 129000 618570
rect 128920 618520 129000 618530
rect 129040 618570 129100 618590
rect 129040 618530 129050 618570
rect 129090 618530 129100 618570
rect 129040 618510 129100 618530
rect 129160 618570 129220 618590
rect 129160 618530 129170 618570
rect 129210 618530 129220 618570
rect 129160 618510 129220 618530
rect 129260 618570 129340 618590
rect 129260 618530 129280 618570
rect 129320 618530 129340 618570
rect 129260 618520 129340 618530
rect 129380 618570 129440 618590
rect 129380 618530 129390 618570
rect 129430 618530 129440 618570
rect 129380 618510 129440 618530
rect 129500 618570 129560 618590
rect 129500 618530 129510 618570
rect 129550 618530 129560 618570
rect 129500 618510 129560 618530
rect 129600 618570 129680 618590
rect 129600 618530 129620 618570
rect 129660 618530 129680 618570
rect 129600 618520 129680 618530
rect 129720 618570 129780 618590
rect 129720 618530 129730 618570
rect 129770 618530 129780 618570
rect 129720 618510 129780 618530
rect 129840 618570 129900 618590
rect 129840 618530 129850 618570
rect 129890 618530 129900 618570
rect 129840 618510 129900 618530
rect 129940 618570 130020 618590
rect 129940 618530 129960 618570
rect 130000 618530 130020 618570
rect 129940 618520 130020 618530
rect 130060 618570 130120 618590
rect 130060 618530 130070 618570
rect 130110 618530 130120 618570
rect 130060 618510 130120 618530
rect 130180 618570 130240 618590
rect 130180 618530 130190 618570
rect 130230 618530 130240 618570
rect 130180 618510 130240 618530
rect 130280 618570 130360 618590
rect 130280 618530 130300 618570
rect 130340 618530 130360 618570
rect 130280 618520 130360 618530
rect 130400 618570 130460 618590
rect 130400 618530 130410 618570
rect 130450 618530 130460 618570
rect 130400 618510 130460 618530
rect 130520 618570 130580 618590
rect 130520 618530 130530 618570
rect 130570 618530 130580 618570
rect 130520 618510 130580 618530
rect 130620 618570 130700 618590
rect 130620 618530 130640 618570
rect 130680 618530 130700 618570
rect 130620 618520 130700 618530
rect 130740 618570 130800 618590
rect 130740 618530 130750 618570
rect 130790 618530 130800 618570
rect 130740 618510 130800 618530
rect 130860 618570 130920 618590
rect 130860 618530 130870 618570
rect 130910 618530 130920 618570
rect 130860 618510 130920 618530
rect 130960 618570 131040 618590
rect 130960 618530 130980 618570
rect 131020 618530 131040 618570
rect 130960 618520 131040 618530
rect 131080 618570 131140 618590
rect 131080 618530 131090 618570
rect 131130 618530 131140 618570
rect 131080 618510 131140 618530
rect 131200 618570 131260 618590
rect 131200 618530 131210 618570
rect 131250 618530 131260 618570
rect 131200 618510 131260 618530
rect 131300 618570 131380 618590
rect 131300 618530 131320 618570
rect 131360 618530 131380 618570
rect 131300 618520 131380 618530
rect 131420 618570 131480 618590
rect 131420 618530 131430 618570
rect 131470 618530 131480 618570
rect 131420 618510 131480 618530
rect 131540 618570 131600 618590
rect 131540 618530 131550 618570
rect 131590 618530 131600 618570
rect 131540 618510 131600 618530
rect 131640 618570 131720 618590
rect 131640 618530 131660 618570
rect 131700 618530 131720 618570
rect 131640 618520 131720 618530
rect 131760 618570 131820 618590
rect 131760 618530 131770 618570
rect 131810 618530 131820 618570
rect 131760 618510 131820 618530
rect 125040 618190 125180 618280
rect 132070 618420 132080 618660
rect 132070 618240 132080 618290
rect 131940 618190 132080 618240
rect 125040 618060 125230 618190
rect 125370 618060 125730 618190
rect 125870 618060 126230 618190
rect 126370 618060 126730 618190
rect 126870 618060 127230 618190
rect 127370 618060 127730 618190
rect 127870 618060 128230 618190
rect 128370 618060 128730 618190
rect 128870 618060 129230 618190
rect 129370 618060 129730 618190
rect 129870 618060 130230 618190
rect 130370 618060 130730 618190
rect 130870 618060 131230 618190
rect 131370 618060 131730 618190
rect 131870 618060 132080 618190
rect 125160 612100 125220 612120
rect 125160 612060 125170 612100
rect 125210 612060 125220 612100
rect 125160 612040 125220 612060
rect 125000 611900 125060 611920
rect 125000 611860 125010 611900
rect 125050 611860 125060 611900
rect 125000 611840 125060 611860
rect 125100 611900 125180 611920
rect 125100 611860 125120 611900
rect 125160 611860 125180 611900
rect 125100 611850 125180 611860
rect 125220 611900 125280 611920
rect 125220 611860 125230 611900
rect 125270 611860 125280 611900
rect 125220 611840 125280 611860
rect 124690 611410 124880 611540
rect 125020 611410 125380 611540
rect 125520 611410 125880 611540
rect 126020 611410 126380 611540
rect 126520 611410 126880 611540
rect 127020 611410 127380 611540
rect 127520 611410 127880 611540
rect 128020 611410 128380 611540
rect 128520 611410 128880 611540
rect 129020 611410 129380 611540
rect 129520 611410 129880 611540
rect 130020 611410 130380 611540
rect 130520 611410 130880 611540
rect 131020 611410 131380 611540
rect 131520 611410 131730 611540
rect 124690 611320 124830 611410
rect 131590 611360 131730 611410
rect 131720 611340 131730 611360
rect 125230 611320 125290 611340
rect 125230 611280 125240 611320
rect 125280 611280 125290 611320
rect 125230 611260 125290 611280
rect 125570 611320 125630 611340
rect 125570 611280 125580 611320
rect 125620 611280 125630 611320
rect 125570 611260 125630 611280
rect 125910 611320 125970 611340
rect 125910 611280 125920 611320
rect 125960 611280 125970 611320
rect 125910 611260 125970 611280
rect 126250 611320 126310 611340
rect 126250 611280 126260 611320
rect 126300 611280 126310 611320
rect 126250 611260 126310 611280
rect 126590 611320 126650 611340
rect 126590 611280 126600 611320
rect 126640 611280 126650 611320
rect 126590 611260 126650 611280
rect 126930 611320 126990 611340
rect 126930 611280 126940 611320
rect 126980 611280 126990 611320
rect 126930 611260 126990 611280
rect 127270 611320 127330 611340
rect 127270 611280 127280 611320
rect 127320 611280 127330 611320
rect 127270 611260 127330 611280
rect 127610 611320 127670 611340
rect 127610 611280 127620 611320
rect 127660 611280 127670 611320
rect 127610 611260 127670 611280
rect 127950 611320 128010 611340
rect 127950 611280 127960 611320
rect 128000 611280 128010 611320
rect 127950 611260 128010 611280
rect 128290 611320 128350 611340
rect 128290 611280 128300 611320
rect 128340 611280 128350 611320
rect 128290 611260 128350 611280
rect 128630 611320 128690 611340
rect 128630 611280 128640 611320
rect 128680 611280 128690 611320
rect 128630 611260 128690 611280
rect 128970 611320 129030 611340
rect 128970 611280 128980 611320
rect 129020 611280 129030 611320
rect 128970 611260 129030 611280
rect 129310 611320 129370 611340
rect 129310 611280 129320 611320
rect 129360 611280 129370 611320
rect 129310 611260 129370 611280
rect 129650 611320 129710 611340
rect 129650 611280 129660 611320
rect 129700 611280 129710 611320
rect 129650 611260 129710 611280
rect 129990 611320 130050 611340
rect 129990 611280 130000 611320
rect 130040 611280 130050 611320
rect 129990 611260 130050 611280
rect 130330 611320 130390 611340
rect 130330 611280 130340 611320
rect 130380 611280 130390 611320
rect 130330 611260 130390 611280
rect 130670 611320 130730 611340
rect 130670 611280 130680 611320
rect 130720 611280 130730 611320
rect 130670 611260 130730 611280
rect 131010 611320 131070 611340
rect 131010 611280 131020 611320
rect 131060 611280 131070 611320
rect 131010 611260 131070 611280
rect 131350 611320 131410 611340
rect 131350 611280 131360 611320
rect 131400 611280 131410 611320
rect 131350 611260 131410 611280
rect 124690 610960 124830 611190
rect 125070 611120 125130 611140
rect 125070 610930 125080 611120
rect 125120 610930 125130 611120
rect 125070 610910 125130 610930
rect 125170 611120 125250 611140
rect 125170 610930 125190 611120
rect 125230 610930 125250 611120
rect 125170 610920 125250 610930
rect 125290 611120 125350 611140
rect 125290 610930 125300 611120
rect 125340 610930 125350 611120
rect 125290 610910 125350 610930
rect 125410 611120 125470 611140
rect 125410 610930 125420 611120
rect 125460 610930 125470 611120
rect 125410 610910 125470 610930
rect 125510 611120 125590 611140
rect 125510 610930 125530 611120
rect 125570 610930 125590 611120
rect 125510 610920 125590 610930
rect 125630 611120 125690 611140
rect 125630 610930 125640 611120
rect 125680 610930 125690 611120
rect 125630 610910 125690 610930
rect 125750 611120 125810 611140
rect 125750 610930 125760 611120
rect 125800 610930 125810 611120
rect 125750 610910 125810 610930
rect 125850 611120 125930 611140
rect 125850 610930 125870 611120
rect 125910 610930 125930 611120
rect 125850 610920 125930 610930
rect 125970 611120 126030 611140
rect 125970 610930 125980 611120
rect 126020 610930 126030 611120
rect 125970 610910 126030 610930
rect 126090 611120 126150 611140
rect 126090 610930 126100 611120
rect 126140 610930 126150 611120
rect 126090 610910 126150 610930
rect 126190 611120 126270 611140
rect 126190 610930 126210 611120
rect 126250 610930 126270 611120
rect 126190 610920 126270 610930
rect 126310 611120 126370 611140
rect 126310 610930 126320 611120
rect 126360 610930 126370 611120
rect 126310 610910 126370 610930
rect 126430 611120 126490 611140
rect 126430 610930 126440 611120
rect 126480 610930 126490 611120
rect 126430 610910 126490 610930
rect 126530 611120 126610 611140
rect 126530 610930 126550 611120
rect 126590 610930 126610 611120
rect 126530 610920 126610 610930
rect 126650 611120 126710 611140
rect 126650 610930 126660 611120
rect 126700 610930 126710 611120
rect 126650 610910 126710 610930
rect 126770 611120 126830 611140
rect 126770 610930 126780 611120
rect 126820 610930 126830 611120
rect 126770 610910 126830 610930
rect 126870 611120 126950 611140
rect 126870 610930 126890 611120
rect 126930 610930 126950 611120
rect 126870 610920 126950 610930
rect 126990 611120 127050 611140
rect 126990 610930 127000 611120
rect 127040 610930 127050 611120
rect 126990 610910 127050 610930
rect 127110 611120 127170 611140
rect 127110 610930 127120 611120
rect 127160 610930 127170 611120
rect 127110 610910 127170 610930
rect 127210 611120 127290 611140
rect 127210 610930 127230 611120
rect 127270 610930 127290 611120
rect 127210 610920 127290 610930
rect 127330 611120 127390 611140
rect 127330 610930 127340 611120
rect 127380 610930 127390 611120
rect 127330 610910 127390 610930
rect 127450 611120 127510 611140
rect 127450 610930 127460 611120
rect 127500 610930 127510 611120
rect 127450 610910 127510 610930
rect 127550 611120 127630 611140
rect 127550 610930 127570 611120
rect 127610 610930 127630 611120
rect 127550 610920 127630 610930
rect 127670 611120 127730 611140
rect 127670 610930 127680 611120
rect 127720 610930 127730 611120
rect 127670 610910 127730 610930
rect 127790 611120 127850 611140
rect 127790 610930 127800 611120
rect 127840 610930 127850 611120
rect 127790 610910 127850 610930
rect 127890 611120 127970 611140
rect 127890 610930 127910 611120
rect 127950 610930 127970 611120
rect 127890 610920 127970 610930
rect 128010 611120 128070 611140
rect 128010 610930 128020 611120
rect 128060 610930 128070 611120
rect 128010 610910 128070 610930
rect 128130 611120 128190 611140
rect 128130 610930 128140 611120
rect 128180 610930 128190 611120
rect 128130 610910 128190 610930
rect 128230 611120 128310 611140
rect 128230 610930 128250 611120
rect 128290 610930 128310 611120
rect 128230 610920 128310 610930
rect 128350 611120 128410 611140
rect 128350 610930 128360 611120
rect 128400 610930 128410 611120
rect 128350 610910 128410 610930
rect 128470 611120 128530 611140
rect 128470 610930 128480 611120
rect 128520 610930 128530 611120
rect 128470 610910 128530 610930
rect 128570 611120 128650 611140
rect 128570 610930 128590 611120
rect 128630 610930 128650 611120
rect 128570 610920 128650 610930
rect 128690 611120 128750 611140
rect 128690 610930 128700 611120
rect 128740 610930 128750 611120
rect 128690 610910 128750 610930
rect 128810 611120 128870 611140
rect 128810 610930 128820 611120
rect 128860 610930 128870 611120
rect 128810 610910 128870 610930
rect 128910 611120 128990 611140
rect 128910 610930 128930 611120
rect 128970 610930 128990 611120
rect 128910 610920 128990 610930
rect 129030 611120 129090 611140
rect 129030 610930 129040 611120
rect 129080 610930 129090 611120
rect 129030 610910 129090 610930
rect 129150 611120 129210 611140
rect 129150 610930 129160 611120
rect 129200 610930 129210 611120
rect 129150 610910 129210 610930
rect 129250 611120 129330 611140
rect 129250 610930 129270 611120
rect 129310 610930 129330 611120
rect 129250 610920 129330 610930
rect 129370 611120 129430 611140
rect 129370 610930 129380 611120
rect 129420 610930 129430 611120
rect 129370 610910 129430 610930
rect 129490 611120 129550 611140
rect 129490 610930 129500 611120
rect 129540 610930 129550 611120
rect 129490 610910 129550 610930
rect 129590 611120 129670 611140
rect 129590 610930 129610 611120
rect 129650 610930 129670 611120
rect 129590 610920 129670 610930
rect 129710 611120 129770 611140
rect 129710 610930 129720 611120
rect 129760 610930 129770 611120
rect 129710 610910 129770 610930
rect 129830 611120 129890 611140
rect 129830 610930 129840 611120
rect 129880 610930 129890 611120
rect 129830 610910 129890 610930
rect 129930 611120 130010 611140
rect 129930 610930 129950 611120
rect 129990 610930 130010 611120
rect 129930 610920 130010 610930
rect 130050 611120 130110 611140
rect 130050 610930 130060 611120
rect 130100 610930 130110 611120
rect 130050 610910 130110 610930
rect 130170 611120 130230 611140
rect 130170 610930 130180 611120
rect 130220 610930 130230 611120
rect 130170 610910 130230 610930
rect 130270 611120 130350 611140
rect 130270 610930 130290 611120
rect 130330 610930 130350 611120
rect 130270 610920 130350 610930
rect 130390 611120 130450 611140
rect 130390 610930 130400 611120
rect 130440 610930 130450 611120
rect 130390 610910 130450 610930
rect 130510 611120 130570 611140
rect 130510 610930 130520 611120
rect 130560 610930 130570 611120
rect 130510 610910 130570 610930
rect 130610 611120 130690 611140
rect 130610 610930 130630 611120
rect 130670 610930 130690 611120
rect 130610 610920 130690 610930
rect 130730 611120 130790 611140
rect 130730 610930 130740 611120
rect 130780 610930 130790 611120
rect 130730 610910 130790 610930
rect 130850 611120 130910 611140
rect 130850 610930 130860 611120
rect 130900 610930 130910 611120
rect 130850 610910 130910 610930
rect 130950 611120 131030 611140
rect 130950 610930 130970 611120
rect 131010 610930 131030 611120
rect 130950 610920 131030 610930
rect 131070 611120 131130 611140
rect 131070 610930 131080 611120
rect 131120 610930 131130 611120
rect 131070 610910 131130 610930
rect 131190 611120 131250 611140
rect 131190 610930 131200 611120
rect 131240 610930 131250 611120
rect 131190 610910 131250 610930
rect 131290 611120 131370 611140
rect 131290 610930 131310 611120
rect 131350 610930 131370 611120
rect 131290 610920 131370 610930
rect 131410 611120 131470 611140
rect 131410 610930 131420 611120
rect 131460 610930 131470 611120
rect 131410 610910 131470 610930
rect 131720 610970 131730 611210
rect 124690 610740 124830 610830
rect 131720 610790 131730 610840
rect 131590 610740 131730 610790
rect 124690 610610 124880 610740
rect 125020 610610 125380 610740
rect 125520 610610 125880 610740
rect 126020 610610 126380 610740
rect 126520 610610 126880 610740
rect 127020 610610 127380 610740
rect 127520 610610 127880 610740
rect 128020 610610 128380 610740
rect 128520 610610 128880 610740
rect 129020 610610 129380 610740
rect 129520 610610 129880 610740
rect 130020 610610 130380 610740
rect 130520 610610 130880 610740
rect 131020 610610 131380 610740
rect 131520 610610 131730 610740
rect 125290 606050 125350 606070
rect 125290 606010 125300 606050
rect 125340 606010 125350 606050
rect 125290 605990 125350 606010
rect 125130 605850 125190 605870
rect 125130 605810 125140 605850
rect 125180 605810 125190 605850
rect 125130 605790 125190 605810
rect 125230 605850 125310 605870
rect 125230 605810 125250 605850
rect 125290 605810 125310 605850
rect 125230 605800 125310 605810
rect 125350 605850 125410 605870
rect 125350 605810 125360 605850
rect 125400 605810 125410 605850
rect 125350 605790 125410 605810
rect 124820 605360 125010 605490
rect 125150 605360 125510 605490
rect 125650 605360 126010 605490
rect 126150 605360 126510 605490
rect 126650 605360 127010 605490
rect 127150 605360 127510 605490
rect 127650 605360 128010 605490
rect 128150 605360 128510 605490
rect 128650 605360 129010 605490
rect 129150 605360 129510 605490
rect 129650 605360 130010 605490
rect 130150 605360 130510 605490
rect 130650 605360 131010 605490
rect 131150 605360 131510 605490
rect 131650 605360 131860 605490
rect 124820 605270 124960 605360
rect 131720 605310 131860 605360
rect 131850 605290 131860 605310
rect 125360 605270 125420 605290
rect 125360 605230 125370 605270
rect 125410 605230 125420 605270
rect 125360 605210 125420 605230
rect 125700 605270 125760 605290
rect 125700 605230 125710 605270
rect 125750 605230 125760 605270
rect 125700 605210 125760 605230
rect 126040 605270 126100 605290
rect 126040 605230 126050 605270
rect 126090 605230 126100 605270
rect 126040 605210 126100 605230
rect 126380 605270 126440 605290
rect 126380 605230 126390 605270
rect 126430 605230 126440 605270
rect 126380 605210 126440 605230
rect 126720 605270 126780 605290
rect 126720 605230 126730 605270
rect 126770 605230 126780 605270
rect 126720 605210 126780 605230
rect 127060 605270 127120 605290
rect 127060 605230 127070 605270
rect 127110 605230 127120 605270
rect 127060 605210 127120 605230
rect 127400 605270 127460 605290
rect 127400 605230 127410 605270
rect 127450 605230 127460 605270
rect 127400 605210 127460 605230
rect 127740 605270 127800 605290
rect 127740 605230 127750 605270
rect 127790 605230 127800 605270
rect 127740 605210 127800 605230
rect 128080 605270 128140 605290
rect 128080 605230 128090 605270
rect 128130 605230 128140 605270
rect 128080 605210 128140 605230
rect 128420 605270 128480 605290
rect 128420 605230 128430 605270
rect 128470 605230 128480 605270
rect 128420 605210 128480 605230
rect 128760 605270 128820 605290
rect 128760 605230 128770 605270
rect 128810 605230 128820 605270
rect 128760 605210 128820 605230
rect 129100 605270 129160 605290
rect 129100 605230 129110 605270
rect 129150 605230 129160 605270
rect 129100 605210 129160 605230
rect 129440 605270 129500 605290
rect 129440 605230 129450 605270
rect 129490 605230 129500 605270
rect 129440 605210 129500 605230
rect 129780 605270 129840 605290
rect 129780 605230 129790 605270
rect 129830 605230 129840 605270
rect 129780 605210 129840 605230
rect 130120 605270 130180 605290
rect 130120 605230 130130 605270
rect 130170 605230 130180 605270
rect 130120 605210 130180 605230
rect 130460 605270 130520 605290
rect 130460 605230 130470 605270
rect 130510 605230 130520 605270
rect 130460 605210 130520 605230
rect 130800 605270 130860 605290
rect 130800 605230 130810 605270
rect 130850 605230 130860 605270
rect 130800 605210 130860 605230
rect 131140 605270 131200 605290
rect 131140 605230 131150 605270
rect 131190 605230 131200 605270
rect 131140 605210 131200 605230
rect 131480 605270 131540 605290
rect 131480 605230 131490 605270
rect 131530 605230 131540 605270
rect 131480 605210 131540 605230
rect 124820 604810 124960 605140
rect 125200 605070 125260 605090
rect 125200 604780 125210 605070
rect 125250 604780 125260 605070
rect 125200 604760 125260 604780
rect 125300 605070 125380 605090
rect 125300 604780 125320 605070
rect 125360 604780 125380 605070
rect 125300 604770 125380 604780
rect 125420 605070 125480 605090
rect 125420 604780 125430 605070
rect 125470 604780 125480 605070
rect 125420 604760 125480 604780
rect 125540 605070 125600 605090
rect 125540 604780 125550 605070
rect 125590 604780 125600 605070
rect 125540 604760 125600 604780
rect 125640 605070 125720 605090
rect 125640 604780 125660 605070
rect 125700 604780 125720 605070
rect 125640 604770 125720 604780
rect 125760 605070 125820 605090
rect 125760 604780 125770 605070
rect 125810 604780 125820 605070
rect 125760 604760 125820 604780
rect 125880 605070 125940 605090
rect 125880 604780 125890 605070
rect 125930 604780 125940 605070
rect 125880 604760 125940 604780
rect 125980 605070 126060 605090
rect 125980 604780 126000 605070
rect 126040 604780 126060 605070
rect 125980 604770 126060 604780
rect 126100 605070 126160 605090
rect 126100 604780 126110 605070
rect 126150 604780 126160 605070
rect 126100 604760 126160 604780
rect 126220 605070 126280 605090
rect 126220 604780 126230 605070
rect 126270 604780 126280 605070
rect 126220 604760 126280 604780
rect 126320 605070 126400 605090
rect 126320 604780 126340 605070
rect 126380 604780 126400 605070
rect 126320 604770 126400 604780
rect 126440 605070 126500 605090
rect 126440 604780 126450 605070
rect 126490 604780 126500 605070
rect 126440 604760 126500 604780
rect 126560 605070 126620 605090
rect 126560 604780 126570 605070
rect 126610 604780 126620 605070
rect 126560 604760 126620 604780
rect 126660 605070 126740 605090
rect 126660 604780 126680 605070
rect 126720 604780 126740 605070
rect 126660 604770 126740 604780
rect 126780 605070 126840 605090
rect 126780 604780 126790 605070
rect 126830 604780 126840 605070
rect 126780 604760 126840 604780
rect 126900 605070 126960 605090
rect 126900 604780 126910 605070
rect 126950 604780 126960 605070
rect 126900 604760 126960 604780
rect 127000 605070 127080 605090
rect 127000 604780 127020 605070
rect 127060 604780 127080 605070
rect 127000 604770 127080 604780
rect 127120 605070 127180 605090
rect 127120 604780 127130 605070
rect 127170 604780 127180 605070
rect 127120 604760 127180 604780
rect 127240 605070 127300 605090
rect 127240 604780 127250 605070
rect 127290 604780 127300 605070
rect 127240 604760 127300 604780
rect 127340 605070 127420 605090
rect 127340 604780 127360 605070
rect 127400 604780 127420 605070
rect 127340 604770 127420 604780
rect 127460 605070 127520 605090
rect 127460 604780 127470 605070
rect 127510 604780 127520 605070
rect 127460 604760 127520 604780
rect 127580 605070 127640 605090
rect 127580 604780 127590 605070
rect 127630 604780 127640 605070
rect 127580 604760 127640 604780
rect 127680 605070 127760 605090
rect 127680 604780 127700 605070
rect 127740 604780 127760 605070
rect 127680 604770 127760 604780
rect 127800 605070 127860 605090
rect 127800 604780 127810 605070
rect 127850 604780 127860 605070
rect 127800 604760 127860 604780
rect 127920 605070 127980 605090
rect 127920 604780 127930 605070
rect 127970 604780 127980 605070
rect 127920 604760 127980 604780
rect 128020 605070 128100 605090
rect 128020 604780 128040 605070
rect 128080 604780 128100 605070
rect 128020 604770 128100 604780
rect 128140 605070 128200 605090
rect 128140 604780 128150 605070
rect 128190 604780 128200 605070
rect 128140 604760 128200 604780
rect 128260 605070 128320 605090
rect 128260 604780 128270 605070
rect 128310 604780 128320 605070
rect 128260 604760 128320 604780
rect 128360 605070 128440 605090
rect 128360 604780 128380 605070
rect 128420 604780 128440 605070
rect 128360 604770 128440 604780
rect 128480 605070 128540 605090
rect 128480 604780 128490 605070
rect 128530 604780 128540 605070
rect 128480 604760 128540 604780
rect 128600 605070 128660 605090
rect 128600 604780 128610 605070
rect 128650 604780 128660 605070
rect 128600 604760 128660 604780
rect 128700 605070 128780 605090
rect 128700 604780 128720 605070
rect 128760 604780 128780 605070
rect 128700 604770 128780 604780
rect 128820 605070 128880 605090
rect 128820 604780 128830 605070
rect 128870 604780 128880 605070
rect 128820 604760 128880 604780
rect 128940 605070 129000 605090
rect 128940 604780 128950 605070
rect 128990 604780 129000 605070
rect 128940 604760 129000 604780
rect 129040 605070 129120 605090
rect 129040 604780 129060 605070
rect 129100 604780 129120 605070
rect 129040 604770 129120 604780
rect 129160 605070 129220 605090
rect 129160 604780 129170 605070
rect 129210 604780 129220 605070
rect 129160 604760 129220 604780
rect 129280 605070 129340 605090
rect 129280 604780 129290 605070
rect 129330 604780 129340 605070
rect 129280 604760 129340 604780
rect 129380 605070 129460 605090
rect 129380 604780 129400 605070
rect 129440 604780 129460 605070
rect 129380 604770 129460 604780
rect 129500 605070 129560 605090
rect 129500 604780 129510 605070
rect 129550 604780 129560 605070
rect 129500 604760 129560 604780
rect 129620 605070 129680 605090
rect 129620 604780 129630 605070
rect 129670 604780 129680 605070
rect 129620 604760 129680 604780
rect 129720 605070 129800 605090
rect 129720 604780 129740 605070
rect 129780 604780 129800 605070
rect 129720 604770 129800 604780
rect 129840 605070 129900 605090
rect 129840 604780 129850 605070
rect 129890 604780 129900 605070
rect 129840 604760 129900 604780
rect 129960 605070 130020 605090
rect 129960 604780 129970 605070
rect 130010 604780 130020 605070
rect 129960 604760 130020 604780
rect 130060 605070 130140 605090
rect 130060 604780 130080 605070
rect 130120 604780 130140 605070
rect 130060 604770 130140 604780
rect 130180 605070 130240 605090
rect 130180 604780 130190 605070
rect 130230 604780 130240 605070
rect 130180 604760 130240 604780
rect 130300 605070 130360 605090
rect 130300 604780 130310 605070
rect 130350 604780 130360 605070
rect 130300 604760 130360 604780
rect 130400 605070 130480 605090
rect 130400 604780 130420 605070
rect 130460 604780 130480 605070
rect 130400 604770 130480 604780
rect 130520 605070 130580 605090
rect 130520 604780 130530 605070
rect 130570 604780 130580 605070
rect 130520 604760 130580 604780
rect 130640 605070 130700 605090
rect 130640 604780 130650 605070
rect 130690 604780 130700 605070
rect 130640 604760 130700 604780
rect 130740 605070 130820 605090
rect 130740 604780 130760 605070
rect 130800 604780 130820 605070
rect 130740 604770 130820 604780
rect 130860 605070 130920 605090
rect 130860 604780 130870 605070
rect 130910 604780 130920 605070
rect 130860 604760 130920 604780
rect 130980 605070 131040 605090
rect 130980 604780 130990 605070
rect 131030 604780 131040 605070
rect 130980 604760 131040 604780
rect 131080 605070 131160 605090
rect 131080 604780 131100 605070
rect 131140 604780 131160 605070
rect 131080 604770 131160 604780
rect 131200 605070 131260 605090
rect 131200 604780 131210 605070
rect 131250 604780 131260 605070
rect 131200 604760 131260 604780
rect 131320 605070 131380 605090
rect 131320 604780 131330 605070
rect 131370 604780 131380 605070
rect 131320 604760 131380 604780
rect 131420 605070 131500 605090
rect 131420 604780 131440 605070
rect 131480 604780 131500 605070
rect 131420 604770 131500 604780
rect 131540 605070 131600 605090
rect 131540 604780 131550 605070
rect 131590 604780 131600 605070
rect 131540 604760 131600 604780
rect 131850 604820 131860 605160
rect 124820 604590 124960 604680
rect 131850 604640 131860 604690
rect 131720 604590 131860 604640
rect 124820 604460 125010 604590
rect 125150 604460 125510 604590
rect 125650 604460 126010 604590
rect 126150 604460 126510 604590
rect 126650 604460 127010 604590
rect 127150 604460 127510 604590
rect 127650 604460 128010 604590
rect 128150 604460 128510 604590
rect 128650 604460 129010 604590
rect 129150 604460 129510 604590
rect 129650 604460 130010 604590
rect 130150 604460 130510 604590
rect 130650 604460 131010 604590
rect 131150 604460 131510 604590
rect 131650 604460 131860 604590
rect 125090 599790 125150 599810
rect 125090 599750 125100 599790
rect 125140 599750 125150 599790
rect 125090 599730 125150 599750
rect 124930 599590 124990 599610
rect 124930 599550 124940 599590
rect 124980 599550 124990 599590
rect 124930 599530 124990 599550
rect 125030 599590 125110 599610
rect 125030 599550 125050 599590
rect 125090 599550 125110 599590
rect 125030 599540 125110 599550
rect 125150 599590 125210 599610
rect 125150 599550 125160 599590
rect 125200 599550 125210 599590
rect 125150 599530 125210 599550
rect 124620 599100 124810 599230
rect 124950 599100 125310 599230
rect 125450 599100 125810 599230
rect 125950 599100 126310 599230
rect 126450 599100 126810 599230
rect 126950 599100 127310 599230
rect 127450 599100 127810 599230
rect 127950 599100 128310 599230
rect 128450 599100 128810 599230
rect 128950 599100 129310 599230
rect 129450 599100 129810 599230
rect 129950 599100 130310 599230
rect 130450 599100 130810 599230
rect 130950 599100 131310 599230
rect 131450 599100 131660 599230
rect 124620 599010 124760 599100
rect 131520 599050 131660 599100
rect 131650 599030 131660 599050
rect 125160 599010 125220 599030
rect 125160 598970 125170 599010
rect 125210 598970 125220 599010
rect 125160 598950 125220 598970
rect 125500 599010 125560 599030
rect 125500 598970 125510 599010
rect 125550 598970 125560 599010
rect 125500 598950 125560 598970
rect 125840 599010 125900 599030
rect 125840 598970 125850 599010
rect 125890 598970 125900 599010
rect 125840 598950 125900 598970
rect 126180 599010 126240 599030
rect 126180 598970 126190 599010
rect 126230 598970 126240 599010
rect 126180 598950 126240 598970
rect 126520 599010 126580 599030
rect 126520 598970 126530 599010
rect 126570 598970 126580 599010
rect 126520 598950 126580 598970
rect 126860 599010 126920 599030
rect 126860 598970 126870 599010
rect 126910 598970 126920 599010
rect 126860 598950 126920 598970
rect 127200 599010 127260 599030
rect 127200 598970 127210 599010
rect 127250 598970 127260 599010
rect 127200 598950 127260 598970
rect 127540 599010 127600 599030
rect 127540 598970 127550 599010
rect 127590 598970 127600 599010
rect 127540 598950 127600 598970
rect 127880 599010 127940 599030
rect 127880 598970 127890 599010
rect 127930 598970 127940 599010
rect 127880 598950 127940 598970
rect 128220 599010 128280 599030
rect 128220 598970 128230 599010
rect 128270 598970 128280 599010
rect 128220 598950 128280 598970
rect 128560 599010 128620 599030
rect 128560 598970 128570 599010
rect 128610 598970 128620 599010
rect 128560 598950 128620 598970
rect 128900 599010 128960 599030
rect 128900 598970 128910 599010
rect 128950 598970 128960 599010
rect 128900 598950 128960 598970
rect 129240 599010 129300 599030
rect 129240 598970 129250 599010
rect 129290 598970 129300 599010
rect 129240 598950 129300 598970
rect 129580 599010 129640 599030
rect 129580 598970 129590 599010
rect 129630 598970 129640 599010
rect 129580 598950 129640 598970
rect 129920 599010 129980 599030
rect 129920 598970 129930 599010
rect 129970 598970 129980 599010
rect 129920 598950 129980 598970
rect 130260 599010 130320 599030
rect 130260 598970 130270 599010
rect 130310 598970 130320 599010
rect 130260 598950 130320 598970
rect 130600 599010 130660 599030
rect 130600 598970 130610 599010
rect 130650 598970 130660 599010
rect 130600 598950 130660 598970
rect 130940 599010 131000 599030
rect 130940 598970 130950 599010
rect 130990 598970 131000 599010
rect 130940 598950 131000 598970
rect 131280 599010 131340 599030
rect 131280 598970 131290 599010
rect 131330 598970 131340 599010
rect 131280 598950 131340 598970
rect 124620 598450 124760 598880
rect 125000 598810 125060 598830
rect 125000 598420 125010 598810
rect 125050 598420 125060 598810
rect 125000 598400 125060 598420
rect 125100 598810 125180 598830
rect 125100 598420 125120 598810
rect 125160 598420 125180 598810
rect 125100 598410 125180 598420
rect 125220 598810 125280 598830
rect 125220 598420 125230 598810
rect 125270 598420 125280 598810
rect 125220 598400 125280 598420
rect 125340 598810 125400 598830
rect 125340 598420 125350 598810
rect 125390 598420 125400 598810
rect 125340 598400 125400 598420
rect 125440 598810 125520 598830
rect 125440 598420 125460 598810
rect 125500 598420 125520 598810
rect 125440 598410 125520 598420
rect 125560 598810 125620 598830
rect 125560 598420 125570 598810
rect 125610 598420 125620 598810
rect 125560 598400 125620 598420
rect 125680 598810 125740 598830
rect 125680 598420 125690 598810
rect 125730 598420 125740 598810
rect 125680 598400 125740 598420
rect 125780 598810 125860 598830
rect 125780 598420 125800 598810
rect 125840 598420 125860 598810
rect 125780 598410 125860 598420
rect 125900 598810 125960 598830
rect 125900 598420 125910 598810
rect 125950 598420 125960 598810
rect 125900 598400 125960 598420
rect 126020 598810 126080 598830
rect 126020 598420 126030 598810
rect 126070 598420 126080 598810
rect 126020 598400 126080 598420
rect 126120 598810 126200 598830
rect 126120 598420 126140 598810
rect 126180 598420 126200 598810
rect 126120 598410 126200 598420
rect 126240 598810 126300 598830
rect 126240 598420 126250 598810
rect 126290 598420 126300 598810
rect 126240 598400 126300 598420
rect 126360 598810 126420 598830
rect 126360 598420 126370 598810
rect 126410 598420 126420 598810
rect 126360 598400 126420 598420
rect 126460 598810 126540 598830
rect 126460 598420 126480 598810
rect 126520 598420 126540 598810
rect 126460 598410 126540 598420
rect 126580 598810 126640 598830
rect 126580 598420 126590 598810
rect 126630 598420 126640 598810
rect 126580 598400 126640 598420
rect 126700 598810 126760 598830
rect 126700 598420 126710 598810
rect 126750 598420 126760 598810
rect 126700 598400 126760 598420
rect 126800 598810 126880 598830
rect 126800 598420 126820 598810
rect 126860 598420 126880 598810
rect 126800 598410 126880 598420
rect 126920 598810 126980 598830
rect 126920 598420 126930 598810
rect 126970 598420 126980 598810
rect 126920 598400 126980 598420
rect 127040 598810 127100 598830
rect 127040 598420 127050 598810
rect 127090 598420 127100 598810
rect 127040 598400 127100 598420
rect 127140 598810 127220 598830
rect 127140 598420 127160 598810
rect 127200 598420 127220 598810
rect 127140 598410 127220 598420
rect 127260 598810 127320 598830
rect 127260 598420 127270 598810
rect 127310 598420 127320 598810
rect 127260 598400 127320 598420
rect 127380 598810 127440 598830
rect 127380 598420 127390 598810
rect 127430 598420 127440 598810
rect 127380 598400 127440 598420
rect 127480 598810 127560 598830
rect 127480 598420 127500 598810
rect 127540 598420 127560 598810
rect 127480 598410 127560 598420
rect 127600 598810 127660 598830
rect 127600 598420 127610 598810
rect 127650 598420 127660 598810
rect 127600 598400 127660 598420
rect 127720 598810 127780 598830
rect 127720 598420 127730 598810
rect 127770 598420 127780 598810
rect 127720 598400 127780 598420
rect 127820 598810 127900 598830
rect 127820 598420 127840 598810
rect 127880 598420 127900 598810
rect 127820 598410 127900 598420
rect 127940 598810 128000 598830
rect 127940 598420 127950 598810
rect 127990 598420 128000 598810
rect 127940 598400 128000 598420
rect 128060 598810 128120 598830
rect 128060 598420 128070 598810
rect 128110 598420 128120 598810
rect 128060 598400 128120 598420
rect 128160 598810 128240 598830
rect 128160 598420 128180 598810
rect 128220 598420 128240 598810
rect 128160 598410 128240 598420
rect 128280 598810 128340 598830
rect 128280 598420 128290 598810
rect 128330 598420 128340 598810
rect 128280 598400 128340 598420
rect 128400 598810 128460 598830
rect 128400 598420 128410 598810
rect 128450 598420 128460 598810
rect 128400 598400 128460 598420
rect 128500 598810 128580 598830
rect 128500 598420 128520 598810
rect 128560 598420 128580 598810
rect 128500 598410 128580 598420
rect 128620 598810 128680 598830
rect 128620 598420 128630 598810
rect 128670 598420 128680 598810
rect 128620 598400 128680 598420
rect 128740 598810 128800 598830
rect 128740 598420 128750 598810
rect 128790 598420 128800 598810
rect 128740 598400 128800 598420
rect 128840 598810 128920 598830
rect 128840 598420 128860 598810
rect 128900 598420 128920 598810
rect 128840 598410 128920 598420
rect 128960 598810 129020 598830
rect 128960 598420 128970 598810
rect 129010 598420 129020 598810
rect 128960 598400 129020 598420
rect 129080 598810 129140 598830
rect 129080 598420 129090 598810
rect 129130 598420 129140 598810
rect 129080 598400 129140 598420
rect 129180 598810 129260 598830
rect 129180 598420 129200 598810
rect 129240 598420 129260 598810
rect 129180 598410 129260 598420
rect 129300 598810 129360 598830
rect 129300 598420 129310 598810
rect 129350 598420 129360 598810
rect 129300 598400 129360 598420
rect 129420 598810 129480 598830
rect 129420 598420 129430 598810
rect 129470 598420 129480 598810
rect 129420 598400 129480 598420
rect 129520 598810 129600 598830
rect 129520 598420 129540 598810
rect 129580 598420 129600 598810
rect 129520 598410 129600 598420
rect 129640 598810 129700 598830
rect 129640 598420 129650 598810
rect 129690 598420 129700 598810
rect 129640 598400 129700 598420
rect 129760 598810 129820 598830
rect 129760 598420 129770 598810
rect 129810 598420 129820 598810
rect 129760 598400 129820 598420
rect 129860 598810 129940 598830
rect 129860 598420 129880 598810
rect 129920 598420 129940 598810
rect 129860 598410 129940 598420
rect 129980 598810 130040 598830
rect 129980 598420 129990 598810
rect 130030 598420 130040 598810
rect 129980 598400 130040 598420
rect 130100 598810 130160 598830
rect 130100 598420 130110 598810
rect 130150 598420 130160 598810
rect 130100 598400 130160 598420
rect 130200 598810 130280 598830
rect 130200 598420 130220 598810
rect 130260 598420 130280 598810
rect 130200 598410 130280 598420
rect 130320 598810 130380 598830
rect 130320 598420 130330 598810
rect 130370 598420 130380 598810
rect 130320 598400 130380 598420
rect 130440 598810 130500 598830
rect 130440 598420 130450 598810
rect 130490 598420 130500 598810
rect 130440 598400 130500 598420
rect 130540 598810 130620 598830
rect 130540 598420 130560 598810
rect 130600 598420 130620 598810
rect 130540 598410 130620 598420
rect 130660 598810 130720 598830
rect 130660 598420 130670 598810
rect 130710 598420 130720 598810
rect 130660 598400 130720 598420
rect 130780 598810 130840 598830
rect 130780 598420 130790 598810
rect 130830 598420 130840 598810
rect 130780 598400 130840 598420
rect 130880 598810 130960 598830
rect 130880 598420 130900 598810
rect 130940 598420 130960 598810
rect 130880 598410 130960 598420
rect 131000 598810 131060 598830
rect 131000 598420 131010 598810
rect 131050 598420 131060 598810
rect 131000 598400 131060 598420
rect 131120 598810 131180 598830
rect 131120 598420 131130 598810
rect 131170 598420 131180 598810
rect 131120 598400 131180 598420
rect 131220 598810 131300 598830
rect 131220 598420 131240 598810
rect 131280 598420 131300 598810
rect 131220 598410 131300 598420
rect 131340 598810 131400 598830
rect 131340 598420 131350 598810
rect 131390 598420 131400 598810
rect 131340 598400 131400 598420
rect 131650 598460 131660 598900
rect 124620 598230 124760 598320
rect 131650 598280 131660 598330
rect 131520 598230 131660 598280
rect 124620 598100 124810 598230
rect 124950 598100 125310 598230
rect 125450 598100 125810 598230
rect 125950 598100 126310 598230
rect 126450 598100 126810 598230
rect 126950 598100 127310 598230
rect 127450 598100 127810 598230
rect 127950 598100 128310 598230
rect 128450 598100 128810 598230
rect 128950 598100 129310 598230
rect 129450 598100 129810 598230
rect 129950 598100 130310 598230
rect 130450 598100 130810 598230
rect 130950 598100 131310 598230
rect 131450 598100 131660 598230
rect 119430 593550 119490 593560
rect 119420 593540 119500 593550
rect 119420 593480 119430 593540
rect 119490 593480 119500 593540
rect 119420 593470 119500 593480
rect 119100 593430 119180 593440
rect 119100 593370 119110 593430
rect 119170 593370 119180 593430
rect 119430 593380 119490 593470
rect 119100 593360 119180 593370
rect 119260 593330 120250 593380
rect 119260 593230 119320 593330
rect 119540 593260 119580 593330
rect 119260 593180 119270 593230
rect 119310 593180 119320 593230
rect 119260 593160 119320 593180
rect 119370 593230 119430 593250
rect 119370 593180 119380 593230
rect 119420 593180 119430 593230
rect 119370 593030 119430 593180
rect 119540 593080 119580 593100
rect 119620 593260 119680 593280
rect 119620 593100 119630 593260
rect 119670 593100 119680 593260
rect 119470 593030 119550 593040
rect 119370 593020 119550 593030
rect 119370 592980 119490 593020
rect 119530 592980 119550 593020
rect 119260 592950 119320 592970
rect 119260 592900 119270 592950
rect 119310 592900 119320 592950
rect 119260 592880 119320 592900
rect 119370 592950 119430 592980
rect 119470 592960 119550 592980
rect 119370 592900 119380 592950
rect 119420 592900 119430 592950
rect 119370 592880 119430 592900
rect 119620 592870 119680 593100
rect 119540 592750 119580 592770
rect 119260 592520 119340 592530
rect 119540 592520 119580 592590
rect 119620 592750 119680 592810
rect 119620 592590 119630 592750
rect 119670 592590 119680 592750
rect 119620 592570 119680 592590
rect 119730 593260 119790 593280
rect 119730 593100 119740 593260
rect 119780 593100 119790 593260
rect 119730 592870 119790 593100
rect 120000 593260 120060 593280
rect 120000 593100 120010 593260
rect 120050 593100 120060 593260
rect 119850 593040 119930 593050
rect 119850 592980 119860 593040
rect 119920 592980 119930 593040
rect 119850 592970 119930 592980
rect 119850 592870 119930 592880
rect 120000 592870 120060 593100
rect 119730 592810 119860 592870
rect 119920 592810 120060 592870
rect 119730 592750 119790 592810
rect 119850 592800 119930 592810
rect 119730 592590 119740 592750
rect 119780 592590 119790 592750
rect 119730 592570 119790 592590
rect 120000 592750 120060 592810
rect 120000 592590 120010 592750
rect 120050 592590 120060 592750
rect 120000 592570 120060 592590
rect 120110 593260 120170 593280
rect 120110 593100 120120 593260
rect 120160 593100 120170 593260
rect 120110 592750 120170 593100
rect 120210 593260 120250 593330
rect 120210 593080 120250 593100
rect 120220 593030 120300 593040
rect 120220 592970 120230 593030
rect 120290 592970 120300 593030
rect 120220 592960 120300 592970
rect 120110 592590 120120 592750
rect 120160 592590 120170 592750
rect 120110 592520 120170 592590
rect 120210 592750 120250 592770
rect 120210 592520 120250 592590
rect 119250 592460 119270 592520
rect 119330 592460 120250 592520
rect 119260 592450 119340 592460
rect 125050 592240 125110 592260
rect 125050 592200 125060 592240
rect 125100 592200 125110 592240
rect 125050 592180 125110 592200
rect 124890 592040 124950 592060
rect 124890 592000 124900 592040
rect 124940 592000 124950 592040
rect 124890 591980 124950 592000
rect 124990 592040 125070 592060
rect 124990 592000 125010 592040
rect 125050 592000 125070 592040
rect 124990 591990 125070 592000
rect 125110 592040 125170 592060
rect 125110 592000 125120 592040
rect 125160 592000 125170 592040
rect 125110 591980 125170 592000
rect 124580 591550 124770 591680
rect 124910 591550 125270 591680
rect 125410 591550 125770 591680
rect 125910 591550 126270 591680
rect 126410 591550 126770 591680
rect 126910 591550 127270 591680
rect 127410 591550 127770 591680
rect 127910 591550 128270 591680
rect 128410 591550 128770 591680
rect 128910 591550 129270 591680
rect 129410 591550 129770 591680
rect 129910 591550 130270 591680
rect 130410 591550 130770 591680
rect 130910 591550 131270 591680
rect 131410 591550 131620 591680
rect 124580 591460 124720 591550
rect 131480 591500 131620 591550
rect 131610 591480 131620 591500
rect 125120 591460 125180 591480
rect 125120 591420 125130 591460
rect 125170 591420 125180 591460
rect 125120 591400 125180 591420
rect 125460 591460 125520 591480
rect 125460 591420 125470 591460
rect 125510 591420 125520 591460
rect 125460 591400 125520 591420
rect 125800 591460 125860 591480
rect 125800 591420 125810 591460
rect 125850 591420 125860 591460
rect 125800 591400 125860 591420
rect 126140 591460 126200 591480
rect 126140 591420 126150 591460
rect 126190 591420 126200 591460
rect 126140 591400 126200 591420
rect 126480 591460 126540 591480
rect 126480 591420 126490 591460
rect 126530 591420 126540 591460
rect 126480 591400 126540 591420
rect 126820 591460 126880 591480
rect 126820 591420 126830 591460
rect 126870 591420 126880 591460
rect 126820 591400 126880 591420
rect 127160 591460 127220 591480
rect 127160 591420 127170 591460
rect 127210 591420 127220 591460
rect 127160 591400 127220 591420
rect 127500 591460 127560 591480
rect 127500 591420 127510 591460
rect 127550 591420 127560 591460
rect 127500 591400 127560 591420
rect 127840 591460 127900 591480
rect 127840 591420 127850 591460
rect 127890 591420 127900 591460
rect 127840 591400 127900 591420
rect 128180 591460 128240 591480
rect 128180 591420 128190 591460
rect 128230 591420 128240 591460
rect 128180 591400 128240 591420
rect 128520 591460 128580 591480
rect 128520 591420 128530 591460
rect 128570 591420 128580 591460
rect 128520 591400 128580 591420
rect 128860 591460 128920 591480
rect 128860 591420 128870 591460
rect 128910 591420 128920 591460
rect 128860 591400 128920 591420
rect 129200 591460 129260 591480
rect 129200 591420 129210 591460
rect 129250 591420 129260 591460
rect 129200 591400 129260 591420
rect 129540 591460 129600 591480
rect 129540 591420 129550 591460
rect 129590 591420 129600 591460
rect 129540 591400 129600 591420
rect 129880 591460 129940 591480
rect 129880 591420 129890 591460
rect 129930 591420 129940 591460
rect 129880 591400 129940 591420
rect 130220 591460 130280 591480
rect 130220 591420 130230 591460
rect 130270 591420 130280 591460
rect 130220 591400 130280 591420
rect 130560 591460 130620 591480
rect 130560 591420 130570 591460
rect 130610 591420 130620 591460
rect 130560 591400 130620 591420
rect 130900 591460 130960 591480
rect 130900 591420 130910 591460
rect 130950 591420 130960 591460
rect 130900 591400 130960 591420
rect 131240 591460 131300 591480
rect 131240 591420 131250 591460
rect 131290 591420 131300 591460
rect 131240 591400 131300 591420
rect 124580 590800 124720 591330
rect 124960 591260 125020 591280
rect 124960 590770 124970 591260
rect 125010 590770 125020 591260
rect 124960 590750 125020 590770
rect 125060 591260 125140 591280
rect 125060 590770 125080 591260
rect 125120 590770 125140 591260
rect 125060 590760 125140 590770
rect 125180 591260 125240 591280
rect 125180 590770 125190 591260
rect 125230 590770 125240 591260
rect 125180 590750 125240 590770
rect 125300 591260 125360 591280
rect 125300 590770 125310 591260
rect 125350 590770 125360 591260
rect 125300 590750 125360 590770
rect 125400 591260 125480 591280
rect 125400 590770 125420 591260
rect 125460 590770 125480 591260
rect 125400 590760 125480 590770
rect 125520 591260 125580 591280
rect 125520 590770 125530 591260
rect 125570 590770 125580 591260
rect 125520 590750 125580 590770
rect 125640 591260 125700 591280
rect 125640 590770 125650 591260
rect 125690 590770 125700 591260
rect 125640 590750 125700 590770
rect 125740 591260 125820 591280
rect 125740 590770 125760 591260
rect 125800 590770 125820 591260
rect 125740 590760 125820 590770
rect 125860 591260 125920 591280
rect 125860 590770 125870 591260
rect 125910 590770 125920 591260
rect 125860 590750 125920 590770
rect 125980 591260 126040 591280
rect 125980 590770 125990 591260
rect 126030 590770 126040 591260
rect 125980 590750 126040 590770
rect 126080 591260 126160 591280
rect 126080 590770 126100 591260
rect 126140 590770 126160 591260
rect 126080 590760 126160 590770
rect 126200 591260 126260 591280
rect 126200 590770 126210 591260
rect 126250 590770 126260 591260
rect 126200 590750 126260 590770
rect 126320 591260 126380 591280
rect 126320 590770 126330 591260
rect 126370 590770 126380 591260
rect 126320 590750 126380 590770
rect 126420 591260 126500 591280
rect 126420 590770 126440 591260
rect 126480 590770 126500 591260
rect 126420 590760 126500 590770
rect 126540 591260 126600 591280
rect 126540 590770 126550 591260
rect 126590 590770 126600 591260
rect 126540 590750 126600 590770
rect 126660 591260 126720 591280
rect 126660 590770 126670 591260
rect 126710 590770 126720 591260
rect 126660 590750 126720 590770
rect 126760 591260 126840 591280
rect 126760 590770 126780 591260
rect 126820 590770 126840 591260
rect 126760 590760 126840 590770
rect 126880 591260 126940 591280
rect 126880 590770 126890 591260
rect 126930 590770 126940 591260
rect 126880 590750 126940 590770
rect 127000 591260 127060 591280
rect 127000 590770 127010 591260
rect 127050 590770 127060 591260
rect 127000 590750 127060 590770
rect 127100 591260 127180 591280
rect 127100 590770 127120 591260
rect 127160 590770 127180 591260
rect 127100 590760 127180 590770
rect 127220 591260 127280 591280
rect 127220 590770 127230 591260
rect 127270 590770 127280 591260
rect 127220 590750 127280 590770
rect 127340 591260 127400 591280
rect 127340 590770 127350 591260
rect 127390 590770 127400 591260
rect 127340 590750 127400 590770
rect 127440 591260 127520 591280
rect 127440 590770 127460 591260
rect 127500 590770 127520 591260
rect 127440 590760 127520 590770
rect 127560 591260 127620 591280
rect 127560 590770 127570 591260
rect 127610 590770 127620 591260
rect 127560 590750 127620 590770
rect 127680 591260 127740 591280
rect 127680 590770 127690 591260
rect 127730 590770 127740 591260
rect 127680 590750 127740 590770
rect 127780 591260 127860 591280
rect 127780 590770 127800 591260
rect 127840 590770 127860 591260
rect 127780 590760 127860 590770
rect 127900 591260 127960 591280
rect 127900 590770 127910 591260
rect 127950 590770 127960 591260
rect 127900 590750 127960 590770
rect 128020 591260 128080 591280
rect 128020 590770 128030 591260
rect 128070 590770 128080 591260
rect 128020 590750 128080 590770
rect 128120 591260 128200 591280
rect 128120 590770 128140 591260
rect 128180 590770 128200 591260
rect 128120 590760 128200 590770
rect 128240 591260 128300 591280
rect 128240 590770 128250 591260
rect 128290 590770 128300 591260
rect 128240 590750 128300 590770
rect 128360 591260 128420 591280
rect 128360 590770 128370 591260
rect 128410 590770 128420 591260
rect 128360 590750 128420 590770
rect 128460 591260 128540 591280
rect 128460 590770 128480 591260
rect 128520 590770 128540 591260
rect 128460 590760 128540 590770
rect 128580 591260 128640 591280
rect 128580 590770 128590 591260
rect 128630 590770 128640 591260
rect 128580 590750 128640 590770
rect 128700 591260 128760 591280
rect 128700 590770 128710 591260
rect 128750 590770 128760 591260
rect 128700 590750 128760 590770
rect 128800 591260 128880 591280
rect 128800 590770 128820 591260
rect 128860 590770 128880 591260
rect 128800 590760 128880 590770
rect 128920 591260 128980 591280
rect 128920 590770 128930 591260
rect 128970 590770 128980 591260
rect 128920 590750 128980 590770
rect 129040 591260 129100 591280
rect 129040 590770 129050 591260
rect 129090 590770 129100 591260
rect 129040 590750 129100 590770
rect 129140 591260 129220 591280
rect 129140 590770 129160 591260
rect 129200 590770 129220 591260
rect 129140 590760 129220 590770
rect 129260 591260 129320 591280
rect 129260 590770 129270 591260
rect 129310 590770 129320 591260
rect 129260 590750 129320 590770
rect 129380 591260 129440 591280
rect 129380 590770 129390 591260
rect 129430 590770 129440 591260
rect 129380 590750 129440 590770
rect 129480 591260 129560 591280
rect 129480 590770 129500 591260
rect 129540 590770 129560 591260
rect 129480 590760 129560 590770
rect 129600 591260 129660 591280
rect 129600 590770 129610 591260
rect 129650 590770 129660 591260
rect 129600 590750 129660 590770
rect 129720 591260 129780 591280
rect 129720 590770 129730 591260
rect 129770 590770 129780 591260
rect 129720 590750 129780 590770
rect 129820 591260 129900 591280
rect 129820 590770 129840 591260
rect 129880 590770 129900 591260
rect 129820 590760 129900 590770
rect 129940 591260 130000 591280
rect 129940 590770 129950 591260
rect 129990 590770 130000 591260
rect 129940 590750 130000 590770
rect 130060 591260 130120 591280
rect 130060 590770 130070 591260
rect 130110 590770 130120 591260
rect 130060 590750 130120 590770
rect 130160 591260 130240 591280
rect 130160 590770 130180 591260
rect 130220 590770 130240 591260
rect 130160 590760 130240 590770
rect 130280 591260 130340 591280
rect 130280 590770 130290 591260
rect 130330 590770 130340 591260
rect 130280 590750 130340 590770
rect 130400 591260 130460 591280
rect 130400 590770 130410 591260
rect 130450 590770 130460 591260
rect 130400 590750 130460 590770
rect 130500 591260 130580 591280
rect 130500 590770 130520 591260
rect 130560 590770 130580 591260
rect 130500 590760 130580 590770
rect 130620 591260 130680 591280
rect 130620 590770 130630 591260
rect 130670 590770 130680 591260
rect 130620 590750 130680 590770
rect 130740 591260 130800 591280
rect 130740 590770 130750 591260
rect 130790 590770 130800 591260
rect 130740 590750 130800 590770
rect 130840 591260 130920 591280
rect 130840 590770 130860 591260
rect 130900 590770 130920 591260
rect 130840 590760 130920 590770
rect 130960 591260 131020 591280
rect 130960 590770 130970 591260
rect 131010 590770 131020 591260
rect 130960 590750 131020 590770
rect 131080 591260 131140 591280
rect 131080 590770 131090 591260
rect 131130 590770 131140 591260
rect 131080 590750 131140 590770
rect 131180 591260 131260 591280
rect 131180 590770 131200 591260
rect 131240 590770 131260 591260
rect 131180 590760 131260 590770
rect 131300 591260 131360 591280
rect 131300 590770 131310 591260
rect 131350 590770 131360 591260
rect 131300 590750 131360 590770
rect 131610 590810 131620 591350
rect 124580 590580 124720 590670
rect 131610 590630 131620 590680
rect 131480 590580 131620 590630
rect 124580 590450 124770 590580
rect 124910 590450 125270 590580
rect 125410 590450 125770 590580
rect 125910 590450 126270 590580
rect 126410 590450 126770 590580
rect 126910 590450 127270 590580
rect 127410 590450 127770 590580
rect 127910 590450 128270 590580
rect 128410 590450 128770 590580
rect 128910 590450 129270 590580
rect 129410 590450 129770 590580
rect 129910 590450 130270 590580
rect 130410 590450 130770 590580
rect 130910 590450 131270 590580
rect 131410 590450 131620 590580
rect 119470 584010 119530 584020
rect 119460 584000 119540 584010
rect 119460 583940 119470 584000
rect 119530 583940 119540 584000
rect 119460 583930 119540 583940
rect 119140 583890 119220 583900
rect 119140 583830 119150 583890
rect 119210 583830 119220 583890
rect 119470 583840 119530 583930
rect 119140 583820 119220 583830
rect 119300 583790 120290 583840
rect 119300 583690 119360 583790
rect 119580 583720 119620 583790
rect 119300 583640 119310 583690
rect 119350 583640 119360 583690
rect 119300 583620 119360 583640
rect 119410 583690 119470 583710
rect 119410 583640 119420 583690
rect 119460 583640 119470 583690
rect 119410 583490 119470 583640
rect 119580 583540 119620 583560
rect 119660 583720 119720 583740
rect 119660 583560 119670 583720
rect 119710 583560 119720 583720
rect 119510 583490 119590 583500
rect 119410 583480 119590 583490
rect 119410 583440 119530 583480
rect 119570 583440 119590 583480
rect 119300 583410 119360 583430
rect 119300 583360 119310 583410
rect 119350 583360 119360 583410
rect 119300 583340 119360 583360
rect 119410 583410 119470 583440
rect 119510 583420 119590 583440
rect 119410 583360 119420 583410
rect 119460 583360 119470 583410
rect 119410 583340 119470 583360
rect 119660 583330 119720 583560
rect 119580 583210 119620 583230
rect 119300 582980 119380 582990
rect 119580 582980 119620 583050
rect 119660 583210 119720 583270
rect 119660 583050 119670 583210
rect 119710 583050 119720 583210
rect 119660 583030 119720 583050
rect 119770 583720 119830 583740
rect 119770 583560 119780 583720
rect 119820 583560 119830 583720
rect 119770 583330 119830 583560
rect 120040 583720 120100 583740
rect 120040 583560 120050 583720
rect 120090 583560 120100 583720
rect 119890 583500 119970 583510
rect 119890 583440 119900 583500
rect 119960 583440 119970 583500
rect 119890 583430 119970 583440
rect 119890 583330 119970 583340
rect 120040 583330 120100 583560
rect 119770 583270 119900 583330
rect 119960 583270 120100 583330
rect 119770 583210 119830 583270
rect 119890 583260 119970 583270
rect 119770 583050 119780 583210
rect 119820 583050 119830 583210
rect 119770 583030 119830 583050
rect 120040 583210 120100 583270
rect 120040 583050 120050 583210
rect 120090 583050 120100 583210
rect 120040 583030 120100 583050
rect 120150 583720 120210 583740
rect 120150 583560 120160 583720
rect 120200 583560 120210 583720
rect 120150 583210 120210 583560
rect 120250 583720 120290 583790
rect 120250 583540 120290 583560
rect 120260 583490 120340 583500
rect 120260 583430 120270 583490
rect 120330 583430 120340 583490
rect 120260 583420 120340 583430
rect 125510 583260 125570 583280
rect 120150 583050 120160 583210
rect 120200 583050 120210 583210
rect 120150 582980 120210 583050
rect 120250 583210 120290 583230
rect 125510 583220 125520 583260
rect 125560 583220 125570 583260
rect 125510 583200 125570 583220
rect 120250 582980 120290 583050
rect 125350 583060 125410 583080
rect 125350 583020 125360 583060
rect 125400 583020 125410 583060
rect 125350 583000 125410 583020
rect 125450 583060 125530 583080
rect 125450 583020 125470 583060
rect 125510 583020 125530 583060
rect 125450 583010 125530 583020
rect 125570 583060 125630 583080
rect 125570 583020 125580 583060
rect 125620 583020 125630 583060
rect 125570 583000 125630 583020
rect 119290 582920 119310 582980
rect 119370 582920 120290 582980
rect 119300 582910 119380 582920
rect 125040 582570 125230 582700
rect 125370 582570 125780 582700
rect 125920 582570 126330 582700
rect 126520 582570 126930 582700
rect 127070 582570 127480 582700
rect 127670 582570 128080 582700
rect 128220 582570 128630 582700
rect 128820 582570 129230 582700
rect 129370 582570 129780 582700
rect 129970 582570 130380 582700
rect 130520 582570 130930 582700
rect 131120 582570 131530 582700
rect 131670 582570 132080 582700
rect 132270 582570 132680 582700
rect 132820 582570 133030 582700
rect 125040 582480 125180 582570
rect 132890 582520 133030 582570
rect 133020 582500 133030 582520
rect 125630 582480 125690 582500
rect 125630 582440 125640 582480
rect 125680 582440 125690 582480
rect 125630 582420 125690 582440
rect 126020 582480 126080 582500
rect 126020 582440 126030 582480
rect 126070 582440 126080 582480
rect 126020 582420 126080 582440
rect 126410 582480 126470 582500
rect 126410 582440 126420 582480
rect 126460 582440 126470 582480
rect 126410 582420 126470 582440
rect 126800 582480 126860 582500
rect 126800 582440 126810 582480
rect 126850 582440 126860 582480
rect 126800 582420 126860 582440
rect 127190 582480 127250 582500
rect 127190 582440 127200 582480
rect 127240 582440 127250 582480
rect 127190 582420 127250 582440
rect 127580 582480 127640 582500
rect 127580 582440 127590 582480
rect 127630 582440 127640 582480
rect 127580 582420 127640 582440
rect 127970 582480 128030 582500
rect 127970 582440 127980 582480
rect 128020 582440 128030 582480
rect 127970 582420 128030 582440
rect 128360 582480 128420 582500
rect 128360 582440 128370 582480
rect 128410 582440 128420 582480
rect 128360 582420 128420 582440
rect 128750 582480 128810 582500
rect 128750 582440 128760 582480
rect 128800 582440 128810 582480
rect 128750 582420 128810 582440
rect 129140 582480 129200 582500
rect 129140 582440 129150 582480
rect 129190 582440 129200 582480
rect 129140 582420 129200 582440
rect 129530 582480 129590 582500
rect 129530 582440 129540 582480
rect 129580 582440 129590 582480
rect 129530 582420 129590 582440
rect 129920 582480 129980 582500
rect 129920 582440 129930 582480
rect 129970 582440 129980 582480
rect 129920 582420 129980 582440
rect 130310 582480 130370 582500
rect 130310 582440 130320 582480
rect 130360 582440 130370 582480
rect 130310 582420 130370 582440
rect 130700 582480 130760 582500
rect 130700 582440 130710 582480
rect 130750 582440 130760 582480
rect 130700 582420 130760 582440
rect 131090 582480 131150 582500
rect 131090 582440 131100 582480
rect 131140 582440 131150 582480
rect 131090 582420 131150 582440
rect 131480 582480 131540 582500
rect 131480 582440 131490 582480
rect 131530 582440 131540 582480
rect 131480 582420 131540 582440
rect 131870 582480 131930 582500
rect 131870 582440 131880 582480
rect 131920 582440 131930 582480
rect 131870 582420 131930 582440
rect 132260 582480 132320 582500
rect 132260 582440 132270 582480
rect 132310 582440 132320 582480
rect 132260 582420 132320 582440
rect 132650 582480 132710 582500
rect 132650 582440 132660 582480
rect 132700 582440 132710 582480
rect 132650 582420 132710 582440
rect 125040 582120 125180 582350
rect 125420 582280 125480 582300
rect 125420 582240 125430 582280
rect 125470 582240 125480 582280
rect 125420 582220 125480 582240
rect 125520 582280 125650 582300
rect 125520 582240 125540 582280
rect 125630 582240 125650 582280
rect 125520 582230 125650 582240
rect 125690 582280 125750 582300
rect 125690 582240 125700 582280
rect 125740 582240 125750 582280
rect 125690 582220 125750 582240
rect 125810 582280 125870 582300
rect 125810 582240 125820 582280
rect 125860 582240 125870 582280
rect 125810 582220 125870 582240
rect 125910 582280 126040 582300
rect 125910 582240 125930 582280
rect 126020 582240 126040 582280
rect 125910 582230 126040 582240
rect 126080 582280 126140 582300
rect 126080 582240 126090 582280
rect 126130 582240 126140 582280
rect 126080 582220 126140 582240
rect 126200 582280 126260 582300
rect 126200 582240 126210 582280
rect 126250 582240 126260 582280
rect 126200 582220 126260 582240
rect 126300 582280 126430 582300
rect 126300 582240 126320 582280
rect 126410 582240 126430 582280
rect 126300 582230 126430 582240
rect 126470 582280 126530 582300
rect 126470 582240 126480 582280
rect 126520 582240 126530 582280
rect 126470 582220 126530 582240
rect 126590 582280 126650 582300
rect 126590 582240 126600 582280
rect 126640 582240 126650 582280
rect 126590 582220 126650 582240
rect 126690 582280 126820 582300
rect 126690 582240 126710 582280
rect 126800 582240 126820 582280
rect 126690 582230 126820 582240
rect 126860 582280 126920 582300
rect 126860 582240 126870 582280
rect 126910 582240 126920 582280
rect 126860 582220 126920 582240
rect 126980 582280 127040 582300
rect 126980 582240 126990 582280
rect 127030 582240 127040 582280
rect 126980 582220 127040 582240
rect 127080 582280 127210 582300
rect 127080 582240 127100 582280
rect 127190 582240 127210 582280
rect 127080 582230 127210 582240
rect 127250 582280 127310 582300
rect 127250 582240 127260 582280
rect 127300 582240 127310 582280
rect 127250 582220 127310 582240
rect 127370 582280 127430 582300
rect 127370 582240 127380 582280
rect 127420 582240 127430 582280
rect 127370 582220 127430 582240
rect 127470 582280 127600 582300
rect 127470 582240 127490 582280
rect 127580 582240 127600 582280
rect 127470 582230 127600 582240
rect 127640 582280 127700 582300
rect 127640 582240 127650 582280
rect 127690 582240 127700 582280
rect 127640 582220 127700 582240
rect 127760 582280 127820 582300
rect 127760 582240 127770 582280
rect 127810 582240 127820 582280
rect 127760 582220 127820 582240
rect 127860 582280 127990 582300
rect 127860 582240 127880 582280
rect 127970 582240 127990 582280
rect 127860 582230 127990 582240
rect 128030 582280 128090 582300
rect 128030 582240 128040 582280
rect 128080 582240 128090 582280
rect 128030 582220 128090 582240
rect 128150 582280 128210 582300
rect 128150 582240 128160 582280
rect 128200 582240 128210 582280
rect 128150 582220 128210 582240
rect 128250 582280 128380 582300
rect 128250 582240 128270 582280
rect 128360 582240 128380 582280
rect 128250 582230 128380 582240
rect 128420 582280 128480 582300
rect 128420 582240 128430 582280
rect 128470 582240 128480 582280
rect 128420 582220 128480 582240
rect 128540 582280 128600 582300
rect 128540 582240 128550 582280
rect 128590 582240 128600 582280
rect 128540 582220 128600 582240
rect 128640 582280 128770 582300
rect 128640 582240 128660 582280
rect 128750 582240 128770 582280
rect 128640 582230 128770 582240
rect 128810 582280 128870 582300
rect 128810 582240 128820 582280
rect 128860 582240 128870 582280
rect 128810 582220 128870 582240
rect 128930 582280 128990 582300
rect 128930 582240 128940 582280
rect 128980 582240 128990 582280
rect 128930 582220 128990 582240
rect 129030 582280 129160 582300
rect 129030 582240 129050 582280
rect 129140 582240 129160 582280
rect 129030 582230 129160 582240
rect 129200 582280 129260 582300
rect 129200 582240 129210 582280
rect 129250 582240 129260 582280
rect 129200 582220 129260 582240
rect 129320 582280 129380 582300
rect 129320 582240 129330 582280
rect 129370 582240 129380 582280
rect 129320 582220 129380 582240
rect 129420 582280 129550 582300
rect 129420 582240 129440 582280
rect 129530 582240 129550 582280
rect 129420 582230 129550 582240
rect 129590 582280 129650 582300
rect 129590 582240 129600 582280
rect 129640 582240 129650 582280
rect 129590 582220 129650 582240
rect 129710 582280 129770 582300
rect 129710 582240 129720 582280
rect 129760 582240 129770 582280
rect 129710 582220 129770 582240
rect 129810 582280 129940 582300
rect 129810 582240 129830 582280
rect 129920 582240 129940 582280
rect 129810 582230 129940 582240
rect 129980 582280 130040 582300
rect 129980 582240 129990 582280
rect 130030 582240 130040 582280
rect 129980 582220 130040 582240
rect 130100 582280 130160 582300
rect 130100 582240 130110 582280
rect 130150 582240 130160 582280
rect 130100 582220 130160 582240
rect 130200 582280 130330 582300
rect 130200 582240 130220 582280
rect 130310 582240 130330 582280
rect 130200 582230 130330 582240
rect 130370 582280 130430 582300
rect 130370 582240 130380 582280
rect 130420 582240 130430 582280
rect 130370 582220 130430 582240
rect 130490 582280 130550 582300
rect 130490 582240 130500 582280
rect 130540 582240 130550 582280
rect 130490 582220 130550 582240
rect 130590 582280 130720 582300
rect 130590 582240 130610 582280
rect 130700 582240 130720 582280
rect 130590 582230 130720 582240
rect 130760 582280 130820 582300
rect 130760 582240 130770 582280
rect 130810 582240 130820 582280
rect 130760 582220 130820 582240
rect 130880 582280 130940 582300
rect 130880 582240 130890 582280
rect 130930 582240 130940 582280
rect 130880 582220 130940 582240
rect 130980 582280 131110 582300
rect 130980 582240 131000 582280
rect 131090 582240 131110 582280
rect 130980 582230 131110 582240
rect 131150 582280 131210 582300
rect 131150 582240 131160 582280
rect 131200 582240 131210 582280
rect 131150 582220 131210 582240
rect 131270 582280 131330 582300
rect 131270 582240 131280 582280
rect 131320 582240 131330 582280
rect 131270 582220 131330 582240
rect 131370 582280 131500 582300
rect 131370 582240 131390 582280
rect 131480 582240 131500 582280
rect 131370 582230 131500 582240
rect 131540 582280 131600 582300
rect 131540 582240 131550 582280
rect 131590 582240 131600 582280
rect 131540 582220 131600 582240
rect 131660 582280 131720 582300
rect 131660 582240 131670 582280
rect 131710 582240 131720 582280
rect 131660 582220 131720 582240
rect 131760 582280 131890 582300
rect 131760 582240 131780 582280
rect 131870 582240 131890 582280
rect 131760 582230 131890 582240
rect 131930 582280 131990 582300
rect 131930 582240 131940 582280
rect 131980 582240 131990 582280
rect 131930 582220 131990 582240
rect 132050 582280 132110 582300
rect 132050 582240 132060 582280
rect 132100 582240 132110 582280
rect 132050 582220 132110 582240
rect 132150 582280 132280 582300
rect 132150 582240 132170 582280
rect 132260 582240 132280 582280
rect 132150 582230 132280 582240
rect 132320 582280 132380 582300
rect 132320 582240 132330 582280
rect 132370 582240 132380 582280
rect 132320 582220 132380 582240
rect 132440 582280 132500 582300
rect 132440 582240 132450 582280
rect 132490 582240 132500 582280
rect 132440 582220 132500 582240
rect 132540 582280 132670 582300
rect 132540 582240 132560 582280
rect 132650 582240 132670 582280
rect 132540 582230 132670 582240
rect 132710 582280 132770 582300
rect 132710 582240 132720 582280
rect 132760 582240 132770 582280
rect 132710 582220 132770 582240
rect 125040 581900 125180 581990
rect 133020 582130 133030 582370
rect 133020 581950 133030 582000
rect 132890 581900 133030 581950
rect 125040 581770 125230 581900
rect 125370 581770 125780 581900
rect 125920 581770 126330 581900
rect 126520 581770 126930 581900
rect 127070 581770 127480 581900
rect 127670 581770 128080 581900
rect 128220 581770 128630 581900
rect 128820 581770 129230 581900
rect 129370 581770 129780 581900
rect 129970 581770 130380 581900
rect 130520 581770 130930 581900
rect 131120 581770 131530 581900
rect 131670 581770 132080 581900
rect 132270 581770 132680 581900
rect 132820 581770 133030 581900
rect 119510 574990 119570 575000
rect 119500 574980 119580 574990
rect 119500 574920 119510 574980
rect 119570 574920 119580 574980
rect 119500 574910 119580 574920
rect 119180 574870 119260 574880
rect 119180 574810 119190 574870
rect 119250 574810 119260 574870
rect 119510 574820 119570 574910
rect 119180 574800 119260 574810
rect 119340 574770 120330 574820
rect 119340 574670 119400 574770
rect 119620 574700 119660 574770
rect 119340 574620 119350 574670
rect 119390 574620 119400 574670
rect 119340 574600 119400 574620
rect 119450 574670 119510 574690
rect 119450 574620 119460 574670
rect 119500 574620 119510 574670
rect 119450 574470 119510 574620
rect 119620 574520 119660 574540
rect 119700 574700 119760 574720
rect 119700 574540 119710 574700
rect 119750 574540 119760 574700
rect 119550 574470 119630 574480
rect 119450 574460 119630 574470
rect 119450 574420 119570 574460
rect 119610 574420 119630 574460
rect 119340 574390 119400 574410
rect 119340 574340 119350 574390
rect 119390 574340 119400 574390
rect 119340 574320 119400 574340
rect 119450 574390 119510 574420
rect 119550 574400 119630 574420
rect 119450 574340 119460 574390
rect 119500 574340 119510 574390
rect 119450 574320 119510 574340
rect 119700 574310 119760 574540
rect 119620 574190 119660 574210
rect 119340 573960 119420 573970
rect 119620 573960 119660 574030
rect 119700 574190 119760 574250
rect 119700 574030 119710 574190
rect 119750 574030 119760 574190
rect 119700 574010 119760 574030
rect 119810 574700 119870 574720
rect 119810 574540 119820 574700
rect 119860 574540 119870 574700
rect 119810 574310 119870 574540
rect 120080 574700 120140 574720
rect 120080 574540 120090 574700
rect 120130 574540 120140 574700
rect 119930 574480 120010 574490
rect 119930 574420 119940 574480
rect 120000 574420 120010 574480
rect 119930 574410 120010 574420
rect 119930 574310 120010 574320
rect 120080 574310 120140 574540
rect 119810 574250 119940 574310
rect 120000 574250 120140 574310
rect 119810 574190 119870 574250
rect 119930 574240 120010 574250
rect 119810 574030 119820 574190
rect 119860 574030 119870 574190
rect 119810 574010 119870 574030
rect 120080 574190 120140 574250
rect 120080 574030 120090 574190
rect 120130 574030 120140 574190
rect 120080 574010 120140 574030
rect 120190 574700 120250 574720
rect 120190 574540 120200 574700
rect 120240 574540 120250 574700
rect 120190 574190 120250 574540
rect 120290 574700 120330 574770
rect 120290 574520 120330 574540
rect 120300 574470 120380 574480
rect 120300 574410 120310 574470
rect 120370 574410 120380 574470
rect 120300 574400 120380 574410
rect 125550 574240 125610 574260
rect 120190 574030 120200 574190
rect 120240 574030 120250 574190
rect 120190 573960 120250 574030
rect 120290 574190 120330 574210
rect 125550 574200 125560 574240
rect 125600 574200 125610 574240
rect 125550 574180 125610 574200
rect 120290 573960 120330 574030
rect 125390 574040 125450 574060
rect 125390 574000 125400 574040
rect 125440 574000 125450 574040
rect 125390 573980 125450 574000
rect 125490 574040 125570 574060
rect 125490 574000 125510 574040
rect 125550 574000 125570 574040
rect 125490 573990 125570 574000
rect 125610 574040 125670 574060
rect 125610 574000 125620 574040
rect 125660 574000 125670 574040
rect 125610 573980 125670 574000
rect 119330 573900 119350 573960
rect 119410 573900 120330 573960
rect 119340 573890 119420 573900
rect 125080 573550 125270 573680
rect 125410 573550 125820 573680
rect 125960 573550 126370 573680
rect 126560 573550 126970 573680
rect 127110 573550 127520 573680
rect 127710 573550 128120 573680
rect 128260 573550 128670 573680
rect 128860 573550 129270 573680
rect 129410 573550 129820 573680
rect 130010 573550 130420 573680
rect 130560 573550 130970 573680
rect 131160 573550 131570 573680
rect 131710 573550 132120 573680
rect 132310 573550 132720 573680
rect 132860 573550 133070 573680
rect 125080 573460 125220 573550
rect 132930 573500 133070 573550
rect 133060 573480 133070 573500
rect 125670 573460 125730 573480
rect 125670 573420 125680 573460
rect 125720 573420 125730 573460
rect 125670 573400 125730 573420
rect 126060 573460 126120 573480
rect 126060 573420 126070 573460
rect 126110 573420 126120 573460
rect 126060 573400 126120 573420
rect 126450 573460 126510 573480
rect 126450 573420 126460 573460
rect 126500 573420 126510 573460
rect 126450 573400 126510 573420
rect 126840 573460 126900 573480
rect 126840 573420 126850 573460
rect 126890 573420 126900 573460
rect 126840 573400 126900 573420
rect 127230 573460 127290 573480
rect 127230 573420 127240 573460
rect 127280 573420 127290 573460
rect 127230 573400 127290 573420
rect 127620 573460 127680 573480
rect 127620 573420 127630 573460
rect 127670 573420 127680 573460
rect 127620 573400 127680 573420
rect 128010 573460 128070 573480
rect 128010 573420 128020 573460
rect 128060 573420 128070 573460
rect 128010 573400 128070 573420
rect 128400 573460 128460 573480
rect 128400 573420 128410 573460
rect 128450 573420 128460 573460
rect 128400 573400 128460 573420
rect 128790 573460 128850 573480
rect 128790 573420 128800 573460
rect 128840 573420 128850 573460
rect 128790 573400 128850 573420
rect 129180 573460 129240 573480
rect 129180 573420 129190 573460
rect 129230 573420 129240 573460
rect 129180 573400 129240 573420
rect 129570 573460 129630 573480
rect 129570 573420 129580 573460
rect 129620 573420 129630 573460
rect 129570 573400 129630 573420
rect 129960 573460 130020 573480
rect 129960 573420 129970 573460
rect 130010 573420 130020 573460
rect 129960 573400 130020 573420
rect 130350 573460 130410 573480
rect 130350 573420 130360 573460
rect 130400 573420 130410 573460
rect 130350 573400 130410 573420
rect 130740 573460 130800 573480
rect 130740 573420 130750 573460
rect 130790 573420 130800 573460
rect 130740 573400 130800 573420
rect 131130 573460 131190 573480
rect 131130 573420 131140 573460
rect 131180 573420 131190 573460
rect 131130 573400 131190 573420
rect 131520 573460 131580 573480
rect 131520 573420 131530 573460
rect 131570 573420 131580 573460
rect 131520 573400 131580 573420
rect 131910 573460 131970 573480
rect 131910 573420 131920 573460
rect 131960 573420 131970 573460
rect 131910 573400 131970 573420
rect 132300 573460 132360 573480
rect 132300 573420 132310 573460
rect 132350 573420 132360 573460
rect 132300 573400 132360 573420
rect 132690 573460 132750 573480
rect 132690 573420 132700 573460
rect 132740 573420 132750 573460
rect 132690 573400 132750 573420
rect 125080 573000 125220 573330
rect 125460 573260 125520 573280
rect 125460 573120 125470 573260
rect 125510 573120 125520 573260
rect 125460 573100 125520 573120
rect 125560 573260 125690 573280
rect 125560 573120 125580 573260
rect 125670 573120 125690 573260
rect 125560 573110 125690 573120
rect 125730 573260 125790 573280
rect 125730 573120 125740 573260
rect 125780 573120 125790 573260
rect 125730 573100 125790 573120
rect 125850 573260 125910 573280
rect 125850 573120 125860 573260
rect 125900 573120 125910 573260
rect 125850 573100 125910 573120
rect 125950 573260 126080 573280
rect 125950 573120 125970 573260
rect 126060 573120 126080 573260
rect 125950 573110 126080 573120
rect 126120 573260 126180 573280
rect 126120 573120 126130 573260
rect 126170 573120 126180 573260
rect 126120 573100 126180 573120
rect 126240 573260 126300 573280
rect 126240 573120 126250 573260
rect 126290 573120 126300 573260
rect 126240 573100 126300 573120
rect 126340 573260 126470 573280
rect 126340 573120 126360 573260
rect 126450 573120 126470 573260
rect 126340 573110 126470 573120
rect 126510 573260 126570 573280
rect 126510 573120 126520 573260
rect 126560 573120 126570 573260
rect 126510 573100 126570 573120
rect 126630 573260 126690 573280
rect 126630 573120 126640 573260
rect 126680 573120 126690 573260
rect 126630 573100 126690 573120
rect 126730 573260 126860 573280
rect 126730 573120 126750 573260
rect 126840 573120 126860 573260
rect 126730 573110 126860 573120
rect 126900 573260 126960 573280
rect 126900 573120 126910 573260
rect 126950 573120 126960 573260
rect 126900 573100 126960 573120
rect 127020 573260 127080 573280
rect 127020 573120 127030 573260
rect 127070 573120 127080 573260
rect 127020 573100 127080 573120
rect 127120 573260 127250 573280
rect 127120 573120 127140 573260
rect 127230 573120 127250 573260
rect 127120 573110 127250 573120
rect 127290 573260 127350 573280
rect 127290 573120 127300 573260
rect 127340 573120 127350 573260
rect 127290 573100 127350 573120
rect 127410 573260 127470 573280
rect 127410 573120 127420 573260
rect 127460 573120 127470 573260
rect 127410 573100 127470 573120
rect 127510 573260 127640 573280
rect 127510 573120 127530 573260
rect 127620 573120 127640 573260
rect 127510 573110 127640 573120
rect 127680 573260 127740 573280
rect 127680 573120 127690 573260
rect 127730 573120 127740 573260
rect 127680 573100 127740 573120
rect 127800 573260 127860 573280
rect 127800 573120 127810 573260
rect 127850 573120 127860 573260
rect 127800 573100 127860 573120
rect 127900 573260 128030 573280
rect 127900 573120 127920 573260
rect 128010 573120 128030 573260
rect 127900 573110 128030 573120
rect 128070 573260 128130 573280
rect 128070 573120 128080 573260
rect 128120 573120 128130 573260
rect 128070 573100 128130 573120
rect 128190 573260 128250 573280
rect 128190 573120 128200 573260
rect 128240 573120 128250 573260
rect 128190 573100 128250 573120
rect 128290 573260 128420 573280
rect 128290 573120 128310 573260
rect 128400 573120 128420 573260
rect 128290 573110 128420 573120
rect 128460 573260 128520 573280
rect 128460 573120 128470 573260
rect 128510 573120 128520 573260
rect 128460 573100 128520 573120
rect 128580 573260 128640 573280
rect 128580 573120 128590 573260
rect 128630 573120 128640 573260
rect 128580 573100 128640 573120
rect 128680 573260 128810 573280
rect 128680 573120 128700 573260
rect 128790 573120 128810 573260
rect 128680 573110 128810 573120
rect 128850 573260 128910 573280
rect 128850 573120 128860 573260
rect 128900 573120 128910 573260
rect 128850 573100 128910 573120
rect 128970 573260 129030 573280
rect 128970 573120 128980 573260
rect 129020 573120 129030 573260
rect 128970 573100 129030 573120
rect 129070 573260 129200 573280
rect 129070 573120 129090 573260
rect 129180 573120 129200 573260
rect 129070 573110 129200 573120
rect 129240 573260 129300 573280
rect 129240 573120 129250 573260
rect 129290 573120 129300 573260
rect 129240 573100 129300 573120
rect 129360 573260 129420 573280
rect 129360 573120 129370 573260
rect 129410 573120 129420 573260
rect 129360 573100 129420 573120
rect 129460 573260 129590 573280
rect 129460 573120 129480 573260
rect 129570 573120 129590 573260
rect 129460 573110 129590 573120
rect 129630 573260 129690 573280
rect 129630 573120 129640 573260
rect 129680 573120 129690 573260
rect 129630 573100 129690 573120
rect 129750 573260 129810 573280
rect 129750 573120 129760 573260
rect 129800 573120 129810 573260
rect 129750 573100 129810 573120
rect 129850 573260 129980 573280
rect 129850 573120 129870 573260
rect 129960 573120 129980 573260
rect 129850 573110 129980 573120
rect 130020 573260 130080 573280
rect 130020 573120 130030 573260
rect 130070 573120 130080 573260
rect 130020 573100 130080 573120
rect 130140 573260 130200 573280
rect 130140 573120 130150 573260
rect 130190 573120 130200 573260
rect 130140 573100 130200 573120
rect 130240 573260 130370 573280
rect 130240 573120 130260 573260
rect 130350 573120 130370 573260
rect 130240 573110 130370 573120
rect 130410 573260 130470 573280
rect 130410 573120 130420 573260
rect 130460 573120 130470 573260
rect 130410 573100 130470 573120
rect 130530 573260 130590 573280
rect 130530 573120 130540 573260
rect 130580 573120 130590 573260
rect 130530 573100 130590 573120
rect 130630 573260 130760 573280
rect 130630 573120 130650 573260
rect 130740 573120 130760 573260
rect 130630 573110 130760 573120
rect 130800 573260 130860 573280
rect 130800 573120 130810 573260
rect 130850 573120 130860 573260
rect 130800 573100 130860 573120
rect 130920 573260 130980 573280
rect 130920 573120 130930 573260
rect 130970 573120 130980 573260
rect 130920 573100 130980 573120
rect 131020 573260 131150 573280
rect 131020 573120 131040 573260
rect 131130 573120 131150 573260
rect 131020 573110 131150 573120
rect 131190 573260 131250 573280
rect 131190 573120 131200 573260
rect 131240 573120 131250 573260
rect 131190 573100 131250 573120
rect 131310 573260 131370 573280
rect 131310 573120 131320 573260
rect 131360 573120 131370 573260
rect 131310 573100 131370 573120
rect 131410 573260 131540 573280
rect 131410 573120 131430 573260
rect 131520 573120 131540 573260
rect 131410 573110 131540 573120
rect 131580 573260 131640 573280
rect 131580 573120 131590 573260
rect 131630 573120 131640 573260
rect 131580 573100 131640 573120
rect 131700 573260 131760 573280
rect 131700 573120 131710 573260
rect 131750 573120 131760 573260
rect 131700 573100 131760 573120
rect 131800 573260 131930 573280
rect 131800 573120 131820 573260
rect 131910 573120 131930 573260
rect 131800 573110 131930 573120
rect 131970 573260 132030 573280
rect 131970 573120 131980 573260
rect 132020 573120 132030 573260
rect 131970 573100 132030 573120
rect 132090 573260 132150 573280
rect 132090 573120 132100 573260
rect 132140 573120 132150 573260
rect 132090 573100 132150 573120
rect 132190 573260 132320 573280
rect 132190 573120 132210 573260
rect 132300 573120 132320 573260
rect 132190 573110 132320 573120
rect 132360 573260 132420 573280
rect 132360 573120 132370 573260
rect 132410 573120 132420 573260
rect 132360 573100 132420 573120
rect 132480 573260 132540 573280
rect 132480 573120 132490 573260
rect 132530 573120 132540 573260
rect 132480 573100 132540 573120
rect 132580 573260 132710 573280
rect 132580 573120 132600 573260
rect 132690 573120 132710 573260
rect 132580 573110 132710 573120
rect 132750 573260 132810 573280
rect 132750 573120 132760 573260
rect 132800 573120 132810 573260
rect 132750 573100 132810 573120
rect 125080 572780 125220 572870
rect 133060 573010 133070 573350
rect 133060 572830 133070 572880
rect 132930 572780 133070 572830
rect 125080 572650 125270 572780
rect 125410 572650 125820 572780
rect 125960 572650 126370 572780
rect 126560 572650 126970 572780
rect 127110 572650 127520 572780
rect 127710 572650 128120 572780
rect 128260 572650 128670 572780
rect 128860 572650 129270 572780
rect 129410 572650 129820 572780
rect 130010 572650 130420 572780
rect 130560 572650 130970 572780
rect 131160 572650 131570 572780
rect 131710 572650 132120 572780
rect 132310 572650 132720 572780
rect 132860 572650 133070 572780
rect 119460 567320 119520 567330
rect 119450 567310 119530 567320
rect 119450 567250 119460 567310
rect 119520 567250 119530 567310
rect 119450 567240 119530 567250
rect 119130 567200 119210 567210
rect 119130 567140 119140 567200
rect 119200 567140 119210 567200
rect 119460 567150 119520 567240
rect 119130 567130 119210 567140
rect 119290 567100 120280 567150
rect 119290 567000 119350 567100
rect 119570 567030 119610 567100
rect 119290 566950 119300 567000
rect 119340 566950 119350 567000
rect 119290 566930 119350 566950
rect 119400 567000 119460 567020
rect 119400 566950 119410 567000
rect 119450 566950 119460 567000
rect 119400 566800 119460 566950
rect 119570 566850 119610 566870
rect 119650 567030 119710 567050
rect 119650 566870 119660 567030
rect 119700 566870 119710 567030
rect 119500 566800 119580 566810
rect 119400 566790 119580 566800
rect 119400 566750 119520 566790
rect 119560 566750 119580 566790
rect 119290 566720 119350 566740
rect 119290 566670 119300 566720
rect 119340 566670 119350 566720
rect 119290 566650 119350 566670
rect 119400 566720 119460 566750
rect 119500 566730 119580 566750
rect 119400 566670 119410 566720
rect 119450 566670 119460 566720
rect 119400 566650 119460 566670
rect 119650 566640 119710 566870
rect 119570 566520 119610 566540
rect 119290 566290 119370 566300
rect 119570 566290 119610 566360
rect 119650 566520 119710 566580
rect 119650 566360 119660 566520
rect 119700 566360 119710 566520
rect 119650 566340 119710 566360
rect 119760 567030 119820 567050
rect 119760 566870 119770 567030
rect 119810 566870 119820 567030
rect 119760 566640 119820 566870
rect 120030 567030 120090 567050
rect 120030 566870 120040 567030
rect 120080 566870 120090 567030
rect 119880 566810 119960 566820
rect 119880 566750 119890 566810
rect 119950 566750 119960 566810
rect 119880 566740 119960 566750
rect 119880 566640 119960 566650
rect 120030 566640 120090 566870
rect 119760 566580 119890 566640
rect 119950 566580 120090 566640
rect 119760 566520 119820 566580
rect 119880 566570 119960 566580
rect 119760 566360 119770 566520
rect 119810 566360 119820 566520
rect 119760 566340 119820 566360
rect 120030 566520 120090 566580
rect 120030 566360 120040 566520
rect 120080 566360 120090 566520
rect 120030 566340 120090 566360
rect 120140 567030 120200 567050
rect 120140 566870 120150 567030
rect 120190 566870 120200 567030
rect 120140 566520 120200 566870
rect 120240 567030 120280 567100
rect 120240 566850 120280 566870
rect 120250 566800 120330 566810
rect 120250 566740 120260 566800
rect 120320 566740 120330 566800
rect 120250 566730 120330 566740
rect 125500 566570 125560 566590
rect 120140 566360 120150 566520
rect 120190 566360 120200 566520
rect 120140 566290 120200 566360
rect 120240 566520 120280 566540
rect 125500 566530 125510 566570
rect 125550 566530 125560 566570
rect 125500 566510 125560 566530
rect 120240 566290 120280 566360
rect 125340 566370 125400 566390
rect 125340 566330 125350 566370
rect 125390 566330 125400 566370
rect 125340 566310 125400 566330
rect 125440 566370 125520 566390
rect 125440 566330 125460 566370
rect 125500 566330 125520 566370
rect 125440 566320 125520 566330
rect 125560 566370 125620 566390
rect 125560 566330 125570 566370
rect 125610 566330 125620 566370
rect 125560 566310 125620 566330
rect 119280 566230 119300 566290
rect 119360 566230 120280 566290
rect 119290 566220 119370 566230
rect 125030 565880 125220 566010
rect 125360 565880 125770 566010
rect 125910 565880 126320 566010
rect 126510 565880 126920 566010
rect 127060 565880 127470 566010
rect 127660 565880 128070 566010
rect 128210 565880 128620 566010
rect 128810 565880 129220 566010
rect 129360 565880 129770 566010
rect 129960 565880 130370 566010
rect 130510 565880 130920 566010
rect 131110 565880 131520 566010
rect 131660 565880 132070 566010
rect 132260 565880 132670 566010
rect 132810 565880 133020 566010
rect 125030 565790 125170 565880
rect 132880 565830 133020 565880
rect 133010 565810 133020 565830
rect 125620 565790 125680 565810
rect 125620 565750 125630 565790
rect 125670 565750 125680 565790
rect 125620 565730 125680 565750
rect 126010 565790 126070 565810
rect 126010 565750 126020 565790
rect 126060 565750 126070 565790
rect 126010 565730 126070 565750
rect 126400 565790 126460 565810
rect 126400 565750 126410 565790
rect 126450 565750 126460 565790
rect 126400 565730 126460 565750
rect 126790 565790 126850 565810
rect 126790 565750 126800 565790
rect 126840 565750 126850 565790
rect 126790 565730 126850 565750
rect 127180 565790 127240 565810
rect 127180 565750 127190 565790
rect 127230 565750 127240 565790
rect 127180 565730 127240 565750
rect 127570 565790 127630 565810
rect 127570 565750 127580 565790
rect 127620 565750 127630 565790
rect 127570 565730 127630 565750
rect 127960 565790 128020 565810
rect 127960 565750 127970 565790
rect 128010 565750 128020 565790
rect 127960 565730 128020 565750
rect 128350 565790 128410 565810
rect 128350 565750 128360 565790
rect 128400 565750 128410 565790
rect 128350 565730 128410 565750
rect 128740 565790 128800 565810
rect 128740 565750 128750 565790
rect 128790 565750 128800 565790
rect 128740 565730 128800 565750
rect 129130 565790 129190 565810
rect 129130 565750 129140 565790
rect 129180 565750 129190 565790
rect 129130 565730 129190 565750
rect 129520 565790 129580 565810
rect 129520 565750 129530 565790
rect 129570 565750 129580 565790
rect 129520 565730 129580 565750
rect 129910 565790 129970 565810
rect 129910 565750 129920 565790
rect 129960 565750 129970 565790
rect 129910 565730 129970 565750
rect 130300 565790 130360 565810
rect 130300 565750 130310 565790
rect 130350 565750 130360 565790
rect 130300 565730 130360 565750
rect 130690 565790 130750 565810
rect 130690 565750 130700 565790
rect 130740 565750 130750 565790
rect 130690 565730 130750 565750
rect 131080 565790 131140 565810
rect 131080 565750 131090 565790
rect 131130 565750 131140 565790
rect 131080 565730 131140 565750
rect 131470 565790 131530 565810
rect 131470 565750 131480 565790
rect 131520 565750 131530 565790
rect 131470 565730 131530 565750
rect 131860 565790 131920 565810
rect 131860 565750 131870 565790
rect 131910 565750 131920 565790
rect 131860 565730 131920 565750
rect 132250 565790 132310 565810
rect 132250 565750 132260 565790
rect 132300 565750 132310 565790
rect 132250 565730 132310 565750
rect 132640 565790 132700 565810
rect 132640 565750 132650 565790
rect 132690 565750 132700 565790
rect 132640 565730 132700 565750
rect 125030 565230 125170 565660
rect 125410 565590 125470 565610
rect 125410 565350 125420 565590
rect 125460 565350 125470 565590
rect 125410 565330 125470 565350
rect 125510 565590 125640 565610
rect 125510 565350 125530 565590
rect 125620 565350 125640 565590
rect 125510 565340 125640 565350
rect 125680 565590 125740 565610
rect 125680 565350 125690 565590
rect 125730 565350 125740 565590
rect 125680 565330 125740 565350
rect 125800 565590 125860 565610
rect 125800 565350 125810 565590
rect 125850 565350 125860 565590
rect 125800 565330 125860 565350
rect 125900 565590 126030 565610
rect 125900 565350 125920 565590
rect 126010 565350 126030 565590
rect 125900 565340 126030 565350
rect 126070 565590 126130 565610
rect 126070 565350 126080 565590
rect 126120 565350 126130 565590
rect 126070 565330 126130 565350
rect 126190 565590 126250 565610
rect 126190 565350 126200 565590
rect 126240 565350 126250 565590
rect 126190 565330 126250 565350
rect 126290 565590 126420 565610
rect 126290 565350 126310 565590
rect 126400 565350 126420 565590
rect 126290 565340 126420 565350
rect 126460 565590 126520 565610
rect 126460 565350 126470 565590
rect 126510 565350 126520 565590
rect 126460 565330 126520 565350
rect 126580 565590 126640 565610
rect 126580 565350 126590 565590
rect 126630 565350 126640 565590
rect 126580 565330 126640 565350
rect 126680 565590 126810 565610
rect 126680 565350 126700 565590
rect 126790 565350 126810 565590
rect 126680 565340 126810 565350
rect 126850 565590 126910 565610
rect 126850 565350 126860 565590
rect 126900 565350 126910 565590
rect 126850 565330 126910 565350
rect 126970 565590 127030 565610
rect 126970 565350 126980 565590
rect 127020 565350 127030 565590
rect 126970 565330 127030 565350
rect 127070 565590 127200 565610
rect 127070 565350 127090 565590
rect 127180 565350 127200 565590
rect 127070 565340 127200 565350
rect 127240 565590 127300 565610
rect 127240 565350 127250 565590
rect 127290 565350 127300 565590
rect 127240 565330 127300 565350
rect 127360 565590 127420 565610
rect 127360 565350 127370 565590
rect 127410 565350 127420 565590
rect 127360 565330 127420 565350
rect 127460 565590 127590 565610
rect 127460 565350 127480 565590
rect 127570 565350 127590 565590
rect 127460 565340 127590 565350
rect 127630 565590 127690 565610
rect 127630 565350 127640 565590
rect 127680 565350 127690 565590
rect 127630 565330 127690 565350
rect 127750 565590 127810 565610
rect 127750 565350 127760 565590
rect 127800 565350 127810 565590
rect 127750 565330 127810 565350
rect 127850 565590 127980 565610
rect 127850 565350 127870 565590
rect 127960 565350 127980 565590
rect 127850 565340 127980 565350
rect 128020 565590 128080 565610
rect 128020 565350 128030 565590
rect 128070 565350 128080 565590
rect 128020 565330 128080 565350
rect 128140 565590 128200 565610
rect 128140 565350 128150 565590
rect 128190 565350 128200 565590
rect 128140 565330 128200 565350
rect 128240 565590 128370 565610
rect 128240 565350 128260 565590
rect 128350 565350 128370 565590
rect 128240 565340 128370 565350
rect 128410 565590 128470 565610
rect 128410 565350 128420 565590
rect 128460 565350 128470 565590
rect 128410 565330 128470 565350
rect 128530 565590 128590 565610
rect 128530 565350 128540 565590
rect 128580 565350 128590 565590
rect 128530 565330 128590 565350
rect 128630 565590 128760 565610
rect 128630 565350 128650 565590
rect 128740 565350 128760 565590
rect 128630 565340 128760 565350
rect 128800 565590 128860 565610
rect 128800 565350 128810 565590
rect 128850 565350 128860 565590
rect 128800 565330 128860 565350
rect 128920 565590 128980 565610
rect 128920 565350 128930 565590
rect 128970 565350 128980 565590
rect 128920 565330 128980 565350
rect 129020 565590 129150 565610
rect 129020 565350 129040 565590
rect 129130 565350 129150 565590
rect 129020 565340 129150 565350
rect 129190 565590 129250 565610
rect 129190 565350 129200 565590
rect 129240 565350 129250 565590
rect 129190 565330 129250 565350
rect 129310 565590 129370 565610
rect 129310 565350 129320 565590
rect 129360 565350 129370 565590
rect 129310 565330 129370 565350
rect 129410 565590 129540 565610
rect 129410 565350 129430 565590
rect 129520 565350 129540 565590
rect 129410 565340 129540 565350
rect 129580 565590 129640 565610
rect 129580 565350 129590 565590
rect 129630 565350 129640 565590
rect 129580 565330 129640 565350
rect 129700 565590 129760 565610
rect 129700 565350 129710 565590
rect 129750 565350 129760 565590
rect 129700 565330 129760 565350
rect 129800 565590 129930 565610
rect 129800 565350 129820 565590
rect 129910 565350 129930 565590
rect 129800 565340 129930 565350
rect 129970 565590 130030 565610
rect 129970 565350 129980 565590
rect 130020 565350 130030 565590
rect 129970 565330 130030 565350
rect 130090 565590 130150 565610
rect 130090 565350 130100 565590
rect 130140 565350 130150 565590
rect 130090 565330 130150 565350
rect 130190 565590 130320 565610
rect 130190 565350 130210 565590
rect 130300 565350 130320 565590
rect 130190 565340 130320 565350
rect 130360 565590 130420 565610
rect 130360 565350 130370 565590
rect 130410 565350 130420 565590
rect 130360 565330 130420 565350
rect 130480 565590 130540 565610
rect 130480 565350 130490 565590
rect 130530 565350 130540 565590
rect 130480 565330 130540 565350
rect 130580 565590 130710 565610
rect 130580 565350 130600 565590
rect 130690 565350 130710 565590
rect 130580 565340 130710 565350
rect 130750 565590 130810 565610
rect 130750 565350 130760 565590
rect 130800 565350 130810 565590
rect 130750 565330 130810 565350
rect 130870 565590 130930 565610
rect 130870 565350 130880 565590
rect 130920 565350 130930 565590
rect 130870 565330 130930 565350
rect 130970 565590 131100 565610
rect 130970 565350 130990 565590
rect 131080 565350 131100 565590
rect 130970 565340 131100 565350
rect 131140 565590 131200 565610
rect 131140 565350 131150 565590
rect 131190 565350 131200 565590
rect 131140 565330 131200 565350
rect 131260 565590 131320 565610
rect 131260 565350 131270 565590
rect 131310 565350 131320 565590
rect 131260 565330 131320 565350
rect 131360 565590 131490 565610
rect 131360 565350 131380 565590
rect 131470 565350 131490 565590
rect 131360 565340 131490 565350
rect 131530 565590 131590 565610
rect 131530 565350 131540 565590
rect 131580 565350 131590 565590
rect 131530 565330 131590 565350
rect 131650 565590 131710 565610
rect 131650 565350 131660 565590
rect 131700 565350 131710 565590
rect 131650 565330 131710 565350
rect 131750 565590 131880 565610
rect 131750 565350 131770 565590
rect 131860 565350 131880 565590
rect 131750 565340 131880 565350
rect 131920 565590 131980 565610
rect 131920 565350 131930 565590
rect 131970 565350 131980 565590
rect 131920 565330 131980 565350
rect 132040 565590 132100 565610
rect 132040 565350 132050 565590
rect 132090 565350 132100 565590
rect 132040 565330 132100 565350
rect 132140 565590 132270 565610
rect 132140 565350 132160 565590
rect 132250 565350 132270 565590
rect 132140 565340 132270 565350
rect 132310 565590 132370 565610
rect 132310 565350 132320 565590
rect 132360 565350 132370 565590
rect 132310 565330 132370 565350
rect 132430 565590 132490 565610
rect 132430 565350 132440 565590
rect 132480 565350 132490 565590
rect 132430 565330 132490 565350
rect 132530 565590 132660 565610
rect 132530 565350 132550 565590
rect 132640 565350 132660 565590
rect 132530 565340 132660 565350
rect 132700 565590 132760 565610
rect 132700 565350 132710 565590
rect 132750 565350 132760 565590
rect 132700 565330 132760 565350
rect 125030 565010 125170 565100
rect 133010 565240 133020 565680
rect 133010 565060 133020 565110
rect 132880 565010 133020 565060
rect 125030 564880 125220 565010
rect 125360 564880 125770 565010
rect 125910 564880 126320 565010
rect 126510 564880 126920 565010
rect 127060 564880 127470 565010
rect 127660 564880 128070 565010
rect 128210 564880 128620 565010
rect 128810 564880 129220 565010
rect 129360 564880 129770 565010
rect 129960 564880 130370 565010
rect 130510 564880 130920 565010
rect 131110 564880 131520 565010
rect 131660 564880 132070 565010
rect 132260 564880 132670 565010
rect 132810 564880 133020 565010
rect 119460 560780 119520 560790
rect 119450 560770 119530 560780
rect 119450 560710 119460 560770
rect 119520 560710 119530 560770
rect 119450 560700 119530 560710
rect 119130 560660 119210 560670
rect 119130 560600 119140 560660
rect 119200 560600 119210 560660
rect 119460 560610 119520 560700
rect 119130 560590 119210 560600
rect 119290 560560 120280 560610
rect 119290 560460 119350 560560
rect 119570 560490 119610 560560
rect 119290 560410 119300 560460
rect 119340 560410 119350 560460
rect 119290 560390 119350 560410
rect 119400 560460 119460 560480
rect 119400 560410 119410 560460
rect 119450 560410 119460 560460
rect 119400 560260 119460 560410
rect 119570 560310 119610 560330
rect 119650 560490 119710 560510
rect 119650 560330 119660 560490
rect 119700 560330 119710 560490
rect 119500 560260 119580 560270
rect 119400 560250 119580 560260
rect 119400 560210 119520 560250
rect 119560 560210 119580 560250
rect 119290 560180 119350 560200
rect 119290 560130 119300 560180
rect 119340 560130 119350 560180
rect 119290 560110 119350 560130
rect 119400 560180 119460 560210
rect 119500 560190 119580 560210
rect 119400 560130 119410 560180
rect 119450 560130 119460 560180
rect 119400 560110 119460 560130
rect 119650 560100 119710 560330
rect 119570 559980 119610 560000
rect 119290 559750 119370 559760
rect 119570 559750 119610 559820
rect 119650 559980 119710 560040
rect 119650 559820 119660 559980
rect 119700 559820 119710 559980
rect 119650 559800 119710 559820
rect 119760 560490 119820 560510
rect 119760 560330 119770 560490
rect 119810 560330 119820 560490
rect 119760 560100 119820 560330
rect 120030 560490 120090 560510
rect 120030 560330 120040 560490
rect 120080 560330 120090 560490
rect 119880 560270 119960 560280
rect 119880 560210 119890 560270
rect 119950 560210 119960 560270
rect 119880 560200 119960 560210
rect 119880 560100 119960 560110
rect 120030 560100 120090 560330
rect 119760 560040 119890 560100
rect 119950 560040 120090 560100
rect 119760 559980 119820 560040
rect 119880 560030 119960 560040
rect 119760 559820 119770 559980
rect 119810 559820 119820 559980
rect 119760 559800 119820 559820
rect 120030 559980 120090 560040
rect 120030 559820 120040 559980
rect 120080 559820 120090 559980
rect 120030 559800 120090 559820
rect 120140 560490 120200 560510
rect 120140 560330 120150 560490
rect 120190 560330 120200 560490
rect 120140 559980 120200 560330
rect 120240 560490 120280 560560
rect 120240 560310 120280 560330
rect 120250 560260 120330 560270
rect 120250 560200 120260 560260
rect 120320 560200 120330 560260
rect 120250 560190 120330 560200
rect 125500 560030 125560 560050
rect 120140 559820 120150 559980
rect 120190 559820 120200 559980
rect 120140 559750 120200 559820
rect 120240 559980 120280 560000
rect 125500 559990 125510 560030
rect 125550 559990 125560 560030
rect 125500 559970 125560 559990
rect 120240 559750 120280 559820
rect 125340 559830 125400 559850
rect 125340 559790 125350 559830
rect 125390 559790 125400 559830
rect 125340 559770 125400 559790
rect 125440 559830 125520 559850
rect 125440 559790 125460 559830
rect 125500 559790 125520 559830
rect 125440 559780 125520 559790
rect 125560 559830 125620 559850
rect 125560 559790 125570 559830
rect 125610 559790 125620 559830
rect 125560 559770 125620 559790
rect 119280 559690 119300 559750
rect 119360 559690 120280 559750
rect 119290 559680 119370 559690
rect 125030 559340 125220 559470
rect 125360 559340 125770 559470
rect 125910 559340 126320 559470
rect 126510 559340 126920 559470
rect 127060 559340 127470 559470
rect 127660 559340 128070 559470
rect 128210 559340 128620 559470
rect 128810 559340 129220 559470
rect 129360 559340 129770 559470
rect 129960 559340 130370 559470
rect 130510 559340 130920 559470
rect 131110 559340 131520 559470
rect 131660 559340 132070 559470
rect 132260 559340 132670 559470
rect 132810 559340 133020 559470
rect 125030 559250 125170 559340
rect 132880 559290 133020 559340
rect 133010 559270 133020 559290
rect 125620 559250 125680 559270
rect 125620 559210 125630 559250
rect 125670 559210 125680 559250
rect 125620 559190 125680 559210
rect 126010 559250 126070 559270
rect 126010 559210 126020 559250
rect 126060 559210 126070 559250
rect 126010 559190 126070 559210
rect 126400 559250 126460 559270
rect 126400 559210 126410 559250
rect 126450 559210 126460 559250
rect 126400 559190 126460 559210
rect 126790 559250 126850 559270
rect 126790 559210 126800 559250
rect 126840 559210 126850 559250
rect 126790 559190 126850 559210
rect 127180 559250 127240 559270
rect 127180 559210 127190 559250
rect 127230 559210 127240 559250
rect 127180 559190 127240 559210
rect 127570 559250 127630 559270
rect 127570 559210 127580 559250
rect 127620 559210 127630 559250
rect 127570 559190 127630 559210
rect 127960 559250 128020 559270
rect 127960 559210 127970 559250
rect 128010 559210 128020 559250
rect 127960 559190 128020 559210
rect 128350 559250 128410 559270
rect 128350 559210 128360 559250
rect 128400 559210 128410 559250
rect 128350 559190 128410 559210
rect 128740 559250 128800 559270
rect 128740 559210 128750 559250
rect 128790 559210 128800 559250
rect 128740 559190 128800 559210
rect 129130 559250 129190 559270
rect 129130 559210 129140 559250
rect 129180 559210 129190 559250
rect 129130 559190 129190 559210
rect 129520 559250 129580 559270
rect 129520 559210 129530 559250
rect 129570 559210 129580 559250
rect 129520 559190 129580 559210
rect 129910 559250 129970 559270
rect 129910 559210 129920 559250
rect 129960 559210 129970 559250
rect 129910 559190 129970 559210
rect 130300 559250 130360 559270
rect 130300 559210 130310 559250
rect 130350 559210 130360 559250
rect 130300 559190 130360 559210
rect 130690 559250 130750 559270
rect 130690 559210 130700 559250
rect 130740 559210 130750 559250
rect 130690 559190 130750 559210
rect 131080 559250 131140 559270
rect 131080 559210 131090 559250
rect 131130 559210 131140 559250
rect 131080 559190 131140 559210
rect 131470 559250 131530 559270
rect 131470 559210 131480 559250
rect 131520 559210 131530 559250
rect 131470 559190 131530 559210
rect 131860 559250 131920 559270
rect 131860 559210 131870 559250
rect 131910 559210 131920 559250
rect 131860 559190 131920 559210
rect 132250 559250 132310 559270
rect 132250 559210 132260 559250
rect 132300 559210 132310 559250
rect 132250 559190 132310 559210
rect 132640 559250 132700 559270
rect 132640 559210 132650 559250
rect 132690 559210 132700 559250
rect 132640 559190 132700 559210
rect 125030 558590 125170 559120
rect 125410 559050 125470 559070
rect 125410 558710 125420 559050
rect 125460 558710 125470 559050
rect 125410 558690 125470 558710
rect 125510 559050 125640 559070
rect 125510 558710 125530 559050
rect 125620 558710 125640 559050
rect 125510 558700 125640 558710
rect 125680 559050 125740 559070
rect 125680 558710 125690 559050
rect 125730 558710 125740 559050
rect 125680 558690 125740 558710
rect 125800 559050 125860 559070
rect 125800 558710 125810 559050
rect 125850 558710 125860 559050
rect 125800 558690 125860 558710
rect 125900 559050 126030 559070
rect 125900 558710 125920 559050
rect 126010 558710 126030 559050
rect 125900 558700 126030 558710
rect 126070 559050 126130 559070
rect 126070 558710 126080 559050
rect 126120 558710 126130 559050
rect 126070 558690 126130 558710
rect 126190 559050 126250 559070
rect 126190 558710 126200 559050
rect 126240 558710 126250 559050
rect 126190 558690 126250 558710
rect 126290 559050 126420 559070
rect 126290 558710 126310 559050
rect 126400 558710 126420 559050
rect 126290 558700 126420 558710
rect 126460 559050 126520 559070
rect 126460 558710 126470 559050
rect 126510 558710 126520 559050
rect 126460 558690 126520 558710
rect 126580 559050 126640 559070
rect 126580 558710 126590 559050
rect 126630 558710 126640 559050
rect 126580 558690 126640 558710
rect 126680 559050 126810 559070
rect 126680 558710 126700 559050
rect 126790 558710 126810 559050
rect 126680 558700 126810 558710
rect 126850 559050 126910 559070
rect 126850 558710 126860 559050
rect 126900 558710 126910 559050
rect 126850 558690 126910 558710
rect 126970 559050 127030 559070
rect 126970 558710 126980 559050
rect 127020 558710 127030 559050
rect 126970 558690 127030 558710
rect 127070 559050 127200 559070
rect 127070 558710 127090 559050
rect 127180 558710 127200 559050
rect 127070 558700 127200 558710
rect 127240 559050 127300 559070
rect 127240 558710 127250 559050
rect 127290 558710 127300 559050
rect 127240 558690 127300 558710
rect 127360 559050 127420 559070
rect 127360 558710 127370 559050
rect 127410 558710 127420 559050
rect 127360 558690 127420 558710
rect 127460 559050 127590 559070
rect 127460 558710 127480 559050
rect 127570 558710 127590 559050
rect 127460 558700 127590 558710
rect 127630 559050 127690 559070
rect 127630 558710 127640 559050
rect 127680 558710 127690 559050
rect 127630 558690 127690 558710
rect 127750 559050 127810 559070
rect 127750 558710 127760 559050
rect 127800 558710 127810 559050
rect 127750 558690 127810 558710
rect 127850 559050 127980 559070
rect 127850 558710 127870 559050
rect 127960 558710 127980 559050
rect 127850 558700 127980 558710
rect 128020 559050 128080 559070
rect 128020 558710 128030 559050
rect 128070 558710 128080 559050
rect 128020 558690 128080 558710
rect 128140 559050 128200 559070
rect 128140 558710 128150 559050
rect 128190 558710 128200 559050
rect 128140 558690 128200 558710
rect 128240 559050 128370 559070
rect 128240 558710 128260 559050
rect 128350 558710 128370 559050
rect 128240 558700 128370 558710
rect 128410 559050 128470 559070
rect 128410 558710 128420 559050
rect 128460 558710 128470 559050
rect 128410 558690 128470 558710
rect 128530 559050 128590 559070
rect 128530 558710 128540 559050
rect 128580 558710 128590 559050
rect 128530 558690 128590 558710
rect 128630 559050 128760 559070
rect 128630 558710 128650 559050
rect 128740 558710 128760 559050
rect 128630 558700 128760 558710
rect 128800 559050 128860 559070
rect 128800 558710 128810 559050
rect 128850 558710 128860 559050
rect 128800 558690 128860 558710
rect 128920 559050 128980 559070
rect 128920 558710 128930 559050
rect 128970 558710 128980 559050
rect 128920 558690 128980 558710
rect 129020 559050 129150 559070
rect 129020 558710 129040 559050
rect 129130 558710 129150 559050
rect 129020 558700 129150 558710
rect 129190 559050 129250 559070
rect 129190 558710 129200 559050
rect 129240 558710 129250 559050
rect 129190 558690 129250 558710
rect 129310 559050 129370 559070
rect 129310 558710 129320 559050
rect 129360 558710 129370 559050
rect 129310 558690 129370 558710
rect 129410 559050 129540 559070
rect 129410 558710 129430 559050
rect 129520 558710 129540 559050
rect 129410 558700 129540 558710
rect 129580 559050 129640 559070
rect 129580 558710 129590 559050
rect 129630 558710 129640 559050
rect 129580 558690 129640 558710
rect 129700 559050 129760 559070
rect 129700 558710 129710 559050
rect 129750 558710 129760 559050
rect 129700 558690 129760 558710
rect 129800 559050 129930 559070
rect 129800 558710 129820 559050
rect 129910 558710 129930 559050
rect 129800 558700 129930 558710
rect 129970 559050 130030 559070
rect 129970 558710 129980 559050
rect 130020 558710 130030 559050
rect 129970 558690 130030 558710
rect 130090 559050 130150 559070
rect 130090 558710 130100 559050
rect 130140 558710 130150 559050
rect 130090 558690 130150 558710
rect 130190 559050 130320 559070
rect 130190 558710 130210 559050
rect 130300 558710 130320 559050
rect 130190 558700 130320 558710
rect 130360 559050 130420 559070
rect 130360 558710 130370 559050
rect 130410 558710 130420 559050
rect 130360 558690 130420 558710
rect 130480 559050 130540 559070
rect 130480 558710 130490 559050
rect 130530 558710 130540 559050
rect 130480 558690 130540 558710
rect 130580 559050 130710 559070
rect 130580 558710 130600 559050
rect 130690 558710 130710 559050
rect 130580 558700 130710 558710
rect 130750 559050 130810 559070
rect 130750 558710 130760 559050
rect 130800 558710 130810 559050
rect 130750 558690 130810 558710
rect 130870 559050 130930 559070
rect 130870 558710 130880 559050
rect 130920 558710 130930 559050
rect 130870 558690 130930 558710
rect 130970 559050 131100 559070
rect 130970 558710 130990 559050
rect 131080 558710 131100 559050
rect 130970 558700 131100 558710
rect 131140 559050 131200 559070
rect 131140 558710 131150 559050
rect 131190 558710 131200 559050
rect 131140 558690 131200 558710
rect 131260 559050 131320 559070
rect 131260 558710 131270 559050
rect 131310 558710 131320 559050
rect 131260 558690 131320 558710
rect 131360 559050 131490 559070
rect 131360 558710 131380 559050
rect 131470 558710 131490 559050
rect 131360 558700 131490 558710
rect 131530 559050 131590 559070
rect 131530 558710 131540 559050
rect 131580 558710 131590 559050
rect 131530 558690 131590 558710
rect 131650 559050 131710 559070
rect 131650 558710 131660 559050
rect 131700 558710 131710 559050
rect 131650 558690 131710 558710
rect 131750 559050 131880 559070
rect 131750 558710 131770 559050
rect 131860 558710 131880 559050
rect 131750 558700 131880 558710
rect 131920 559050 131980 559070
rect 131920 558710 131930 559050
rect 131970 558710 131980 559050
rect 131920 558690 131980 558710
rect 132040 559050 132100 559070
rect 132040 558710 132050 559050
rect 132090 558710 132100 559050
rect 132040 558690 132100 558710
rect 132140 559050 132270 559070
rect 132140 558710 132160 559050
rect 132250 558710 132270 559050
rect 132140 558700 132270 558710
rect 132310 559050 132370 559070
rect 132310 558710 132320 559050
rect 132360 558710 132370 559050
rect 132310 558690 132370 558710
rect 132430 559050 132490 559070
rect 132430 558710 132440 559050
rect 132480 558710 132490 559050
rect 132430 558690 132490 558710
rect 132530 559050 132660 559070
rect 132530 558710 132550 559050
rect 132640 558710 132660 559050
rect 132530 558700 132660 558710
rect 132700 559050 132760 559070
rect 132700 558710 132710 559050
rect 132750 558710 132760 559050
rect 132700 558690 132760 558710
rect 125030 558370 125170 558460
rect 133010 558600 133020 559140
rect 133010 558420 133020 558470
rect 132880 558370 133020 558420
rect 125030 558240 125220 558370
rect 125360 558240 125770 558370
rect 125910 558240 126320 558370
rect 126510 558240 126920 558370
rect 127060 558240 127470 558370
rect 127660 558240 128070 558370
rect 128210 558240 128620 558370
rect 128810 558240 129220 558370
rect 129360 558240 129770 558370
rect 129960 558240 130370 558370
rect 130510 558240 130920 558370
rect 131110 558240 131520 558370
rect 131660 558240 132070 558370
rect 132260 558240 132670 558370
rect 132810 558240 133020 558370
rect 125150 554170 125210 554190
rect 125150 554130 125160 554170
rect 125200 554130 125210 554170
rect 125150 554110 125210 554130
rect 124990 553970 125050 553990
rect 119530 553950 119590 553960
rect 119520 553940 119600 553950
rect 119520 553880 119530 553940
rect 119590 553880 119600 553940
rect 124990 553930 125000 553970
rect 125040 553930 125050 553970
rect 124990 553910 125050 553930
rect 125090 553970 125170 553990
rect 125090 553930 125110 553970
rect 125150 553930 125170 553970
rect 125090 553920 125170 553930
rect 125210 553970 125270 553990
rect 125210 553930 125220 553970
rect 125260 553930 125270 553970
rect 125210 553910 125270 553930
rect 119520 553870 119600 553880
rect 119200 553830 119280 553840
rect 119200 553770 119210 553830
rect 119270 553770 119280 553830
rect 119530 553780 119590 553870
rect 119200 553760 119280 553770
rect 119360 553730 120350 553780
rect 119360 553630 119420 553730
rect 119640 553660 119680 553730
rect 119360 553580 119370 553630
rect 119410 553580 119420 553630
rect 119360 553560 119420 553580
rect 119470 553630 119530 553650
rect 119470 553580 119480 553630
rect 119520 553580 119530 553630
rect 119470 553430 119530 553580
rect 119640 553480 119680 553500
rect 119720 553660 119780 553680
rect 119720 553500 119730 553660
rect 119770 553500 119780 553660
rect 119570 553430 119650 553440
rect 119470 553420 119650 553430
rect 119470 553380 119590 553420
rect 119630 553380 119650 553420
rect 119360 553350 119420 553370
rect 119360 553300 119370 553350
rect 119410 553300 119420 553350
rect 119360 553280 119420 553300
rect 119470 553350 119530 553380
rect 119570 553360 119650 553380
rect 119470 553300 119480 553350
rect 119520 553300 119530 553350
rect 119470 553280 119530 553300
rect 119720 553270 119780 553500
rect 119640 553150 119680 553170
rect 119360 552920 119440 552930
rect 119640 552920 119680 552990
rect 119720 553150 119780 553210
rect 119720 552990 119730 553150
rect 119770 552990 119780 553150
rect 119720 552970 119780 552990
rect 119830 553660 119890 553680
rect 119830 553500 119840 553660
rect 119880 553500 119890 553660
rect 119830 553270 119890 553500
rect 120100 553660 120160 553680
rect 120100 553500 120110 553660
rect 120150 553500 120160 553660
rect 119950 553440 120030 553450
rect 119950 553380 119960 553440
rect 120020 553380 120030 553440
rect 119950 553370 120030 553380
rect 119950 553270 120030 553280
rect 120100 553270 120160 553500
rect 119830 553210 119960 553270
rect 120020 553210 120160 553270
rect 119830 553150 119890 553210
rect 119950 553200 120030 553210
rect 119830 552990 119840 553150
rect 119880 552990 119890 553150
rect 119830 552970 119890 552990
rect 120100 553150 120160 553210
rect 120100 552990 120110 553150
rect 120150 552990 120160 553150
rect 120100 552970 120160 552990
rect 120210 553660 120270 553680
rect 120210 553500 120220 553660
rect 120260 553500 120270 553660
rect 120210 553150 120270 553500
rect 120310 553660 120350 553730
rect 120310 553480 120350 553500
rect 120320 553430 120400 553440
rect 120320 553370 120330 553430
rect 120390 553370 120400 553430
rect 120320 553360 120400 553370
rect 120210 552990 120220 553150
rect 120260 552990 120270 553150
rect 120210 552920 120270 552990
rect 120310 553150 120350 553170
rect 120310 552920 120350 552990
rect 119350 552860 119370 552920
rect 119430 552860 120350 552920
rect 119360 552850 119440 552860
rect 125100 552510 125290 552640
rect 125430 552510 125890 552640
rect 126030 552510 126490 552640
rect 126730 552510 127190 552640
rect 127330 552510 127790 552640
rect 128030 552510 128490 552640
rect 128630 552510 129090 552640
rect 129330 552510 129790 552640
rect 129930 552510 130390 552640
rect 130630 552510 131090 552640
rect 131230 552510 131690 552640
rect 131930 552510 132390 552640
rect 132530 552510 132990 552640
rect 133230 552510 133690 552640
rect 133830 552510 134040 552640
rect 125100 552420 125240 552510
rect 133900 552460 134040 552510
rect 134030 552440 134040 552460
rect 125740 552420 125800 552440
rect 125740 552380 125750 552420
rect 125790 552380 125800 552420
rect 125740 552360 125800 552380
rect 126180 552420 126240 552440
rect 126180 552380 126190 552420
rect 126230 552380 126240 552420
rect 126180 552360 126240 552380
rect 126620 552420 126680 552440
rect 126620 552380 126630 552420
rect 126670 552380 126680 552420
rect 126620 552360 126680 552380
rect 127060 552420 127120 552440
rect 127060 552380 127070 552420
rect 127110 552380 127120 552420
rect 127060 552360 127120 552380
rect 127500 552420 127560 552440
rect 127500 552380 127510 552420
rect 127550 552380 127560 552420
rect 127500 552360 127560 552380
rect 127940 552420 128000 552440
rect 127940 552380 127950 552420
rect 127990 552380 128000 552420
rect 127940 552360 128000 552380
rect 128380 552420 128440 552440
rect 128380 552380 128390 552420
rect 128430 552380 128440 552420
rect 128380 552360 128440 552380
rect 128820 552420 128880 552440
rect 128820 552380 128830 552420
rect 128870 552380 128880 552420
rect 128820 552360 128880 552380
rect 129260 552420 129320 552440
rect 129260 552380 129270 552420
rect 129310 552380 129320 552420
rect 129260 552360 129320 552380
rect 129700 552420 129760 552440
rect 129700 552380 129710 552420
rect 129750 552380 129760 552420
rect 129700 552360 129760 552380
rect 130140 552420 130200 552440
rect 130140 552380 130150 552420
rect 130190 552380 130200 552420
rect 130140 552360 130200 552380
rect 130580 552420 130640 552440
rect 130580 552380 130590 552420
rect 130630 552380 130640 552420
rect 130580 552360 130640 552380
rect 131020 552420 131080 552440
rect 131020 552380 131030 552420
rect 131070 552380 131080 552420
rect 131020 552360 131080 552380
rect 131460 552420 131520 552440
rect 131460 552380 131470 552420
rect 131510 552380 131520 552420
rect 131460 552360 131520 552380
rect 131900 552420 131960 552440
rect 131900 552380 131910 552420
rect 131950 552380 131960 552420
rect 131900 552360 131960 552380
rect 132340 552420 132400 552440
rect 132340 552380 132350 552420
rect 132390 552380 132400 552420
rect 132340 552360 132400 552380
rect 132780 552420 132840 552440
rect 132780 552380 132790 552420
rect 132830 552380 132840 552420
rect 132780 552360 132840 552380
rect 133220 552420 133280 552440
rect 133220 552380 133230 552420
rect 133270 552380 133280 552420
rect 133220 552360 133280 552380
rect 133660 552420 133720 552440
rect 133660 552380 133670 552420
rect 133710 552380 133720 552420
rect 133660 552360 133720 552380
rect 125100 552060 125240 552290
rect 125480 552220 125540 552240
rect 125480 552180 125490 552220
rect 125530 552180 125540 552220
rect 125480 552160 125540 552180
rect 125580 552220 125760 552240
rect 125580 552180 125600 552220
rect 125740 552180 125760 552220
rect 125580 552170 125760 552180
rect 125800 552220 125860 552240
rect 125800 552180 125810 552220
rect 125850 552180 125860 552220
rect 125800 552160 125860 552180
rect 125920 552220 125980 552240
rect 125920 552180 125930 552220
rect 125970 552180 125980 552220
rect 125920 552160 125980 552180
rect 126020 552220 126200 552240
rect 126020 552180 126040 552220
rect 126180 552180 126200 552220
rect 126020 552170 126200 552180
rect 126240 552220 126300 552240
rect 126240 552180 126250 552220
rect 126290 552180 126300 552220
rect 126240 552160 126300 552180
rect 126360 552220 126420 552240
rect 126360 552180 126370 552220
rect 126410 552180 126420 552220
rect 126360 552160 126420 552180
rect 126460 552220 126640 552240
rect 126460 552180 126480 552220
rect 126620 552180 126640 552220
rect 126460 552170 126640 552180
rect 126680 552220 126740 552240
rect 126680 552180 126690 552220
rect 126730 552180 126740 552220
rect 126680 552160 126740 552180
rect 126800 552220 126860 552240
rect 126800 552180 126810 552220
rect 126850 552180 126860 552220
rect 126800 552160 126860 552180
rect 126900 552220 127080 552240
rect 126900 552180 126920 552220
rect 127060 552180 127080 552220
rect 126900 552170 127080 552180
rect 127120 552220 127180 552240
rect 127120 552180 127130 552220
rect 127170 552180 127180 552220
rect 127120 552160 127180 552180
rect 127240 552220 127300 552240
rect 127240 552180 127250 552220
rect 127290 552180 127300 552220
rect 127240 552160 127300 552180
rect 127340 552220 127520 552240
rect 127340 552180 127360 552220
rect 127500 552180 127520 552220
rect 127340 552170 127520 552180
rect 127560 552220 127620 552240
rect 127560 552180 127570 552220
rect 127610 552180 127620 552220
rect 127560 552160 127620 552180
rect 127680 552220 127740 552240
rect 127680 552180 127690 552220
rect 127730 552180 127740 552220
rect 127680 552160 127740 552180
rect 127780 552220 127960 552240
rect 127780 552180 127800 552220
rect 127940 552180 127960 552220
rect 127780 552170 127960 552180
rect 128000 552220 128060 552240
rect 128000 552180 128010 552220
rect 128050 552180 128060 552220
rect 128000 552160 128060 552180
rect 128120 552220 128180 552240
rect 128120 552180 128130 552220
rect 128170 552180 128180 552220
rect 128120 552160 128180 552180
rect 128220 552220 128400 552240
rect 128220 552180 128240 552220
rect 128380 552180 128400 552220
rect 128220 552170 128400 552180
rect 128440 552220 128500 552240
rect 128440 552180 128450 552220
rect 128490 552180 128500 552220
rect 128440 552160 128500 552180
rect 128560 552220 128620 552240
rect 128560 552180 128570 552220
rect 128610 552180 128620 552220
rect 128560 552160 128620 552180
rect 128660 552220 128840 552240
rect 128660 552180 128680 552220
rect 128820 552180 128840 552220
rect 128660 552170 128840 552180
rect 128880 552220 128940 552240
rect 128880 552180 128890 552220
rect 128930 552180 128940 552220
rect 128880 552160 128940 552180
rect 129000 552220 129060 552240
rect 129000 552180 129010 552220
rect 129050 552180 129060 552220
rect 129000 552160 129060 552180
rect 129100 552220 129280 552240
rect 129100 552180 129120 552220
rect 129260 552180 129280 552220
rect 129100 552170 129280 552180
rect 129320 552220 129380 552240
rect 129320 552180 129330 552220
rect 129370 552180 129380 552220
rect 129320 552160 129380 552180
rect 129440 552220 129500 552240
rect 129440 552180 129450 552220
rect 129490 552180 129500 552220
rect 129440 552160 129500 552180
rect 129540 552220 129720 552240
rect 129540 552180 129560 552220
rect 129700 552180 129720 552220
rect 129540 552170 129720 552180
rect 129760 552220 129820 552240
rect 129760 552180 129770 552220
rect 129810 552180 129820 552220
rect 129760 552160 129820 552180
rect 129880 552220 129940 552240
rect 129880 552180 129890 552220
rect 129930 552180 129940 552220
rect 129880 552160 129940 552180
rect 129980 552220 130160 552240
rect 129980 552180 130000 552220
rect 130140 552180 130160 552220
rect 129980 552170 130160 552180
rect 130200 552220 130260 552240
rect 130200 552180 130210 552220
rect 130250 552180 130260 552220
rect 130200 552160 130260 552180
rect 130320 552220 130380 552240
rect 130320 552180 130330 552220
rect 130370 552180 130380 552220
rect 130320 552160 130380 552180
rect 130420 552220 130600 552240
rect 130420 552180 130440 552220
rect 130580 552180 130600 552220
rect 130420 552170 130600 552180
rect 130640 552220 130700 552240
rect 130640 552180 130650 552220
rect 130690 552180 130700 552220
rect 130640 552160 130700 552180
rect 130760 552220 130820 552240
rect 130760 552180 130770 552220
rect 130810 552180 130820 552220
rect 130760 552160 130820 552180
rect 130860 552220 131040 552240
rect 130860 552180 130880 552220
rect 131020 552180 131040 552220
rect 130860 552170 131040 552180
rect 131080 552220 131140 552240
rect 131080 552180 131090 552220
rect 131130 552180 131140 552220
rect 131080 552160 131140 552180
rect 131200 552220 131260 552240
rect 131200 552180 131210 552220
rect 131250 552180 131260 552220
rect 131200 552160 131260 552180
rect 131300 552220 131480 552240
rect 131300 552180 131320 552220
rect 131460 552180 131480 552220
rect 131300 552170 131480 552180
rect 131520 552220 131580 552240
rect 131520 552180 131530 552220
rect 131570 552180 131580 552220
rect 131520 552160 131580 552180
rect 131640 552220 131700 552240
rect 131640 552180 131650 552220
rect 131690 552180 131700 552220
rect 131640 552160 131700 552180
rect 131740 552220 131920 552240
rect 131740 552180 131760 552220
rect 131900 552180 131920 552220
rect 131740 552170 131920 552180
rect 131960 552220 132020 552240
rect 131960 552180 131970 552220
rect 132010 552180 132020 552220
rect 131960 552160 132020 552180
rect 132080 552220 132140 552240
rect 132080 552180 132090 552220
rect 132130 552180 132140 552220
rect 132080 552160 132140 552180
rect 132180 552220 132360 552240
rect 132180 552180 132200 552220
rect 132340 552180 132360 552220
rect 132180 552170 132360 552180
rect 132400 552220 132460 552240
rect 132400 552180 132410 552220
rect 132450 552180 132460 552220
rect 132400 552160 132460 552180
rect 132520 552220 132580 552240
rect 132520 552180 132530 552220
rect 132570 552180 132580 552220
rect 132520 552160 132580 552180
rect 132620 552220 132800 552240
rect 132620 552180 132640 552220
rect 132780 552180 132800 552220
rect 132620 552170 132800 552180
rect 132840 552220 132900 552240
rect 132840 552180 132850 552220
rect 132890 552180 132900 552220
rect 132840 552160 132900 552180
rect 132960 552220 133020 552240
rect 132960 552180 132970 552220
rect 133010 552180 133020 552220
rect 132960 552160 133020 552180
rect 133060 552220 133240 552240
rect 133060 552180 133080 552220
rect 133220 552180 133240 552220
rect 133060 552170 133240 552180
rect 133280 552220 133340 552240
rect 133280 552180 133290 552220
rect 133330 552180 133340 552220
rect 133280 552160 133340 552180
rect 133400 552220 133460 552240
rect 133400 552180 133410 552220
rect 133450 552180 133460 552220
rect 133400 552160 133460 552180
rect 133500 552220 133680 552240
rect 133500 552180 133520 552220
rect 133660 552180 133680 552220
rect 133500 552170 133680 552180
rect 133720 552220 133780 552240
rect 133720 552180 133730 552220
rect 133770 552180 133780 552220
rect 133720 552160 133780 552180
rect 125100 551840 125240 551930
rect 134030 552070 134040 552310
rect 134030 551890 134040 551940
rect 133900 551840 134040 551890
rect 125100 551710 125290 551840
rect 125430 551710 125890 551840
rect 126030 551710 126490 551840
rect 126730 551710 127190 551840
rect 127330 551710 127790 551840
rect 128030 551710 128490 551840
rect 128630 551710 129090 551840
rect 129330 551710 129790 551840
rect 129930 551710 130390 551840
rect 130630 551710 131090 551840
rect 131230 551710 131690 551840
rect 131930 551710 132390 551840
rect 132530 551710 132990 551840
rect 133230 551710 133690 551840
rect 133830 551710 134040 551840
rect 125150 546600 125210 546620
rect 125150 546560 125160 546600
rect 125200 546560 125210 546600
rect 125150 546540 125210 546560
rect 124990 546400 125050 546420
rect 119530 546380 119590 546390
rect 119520 546370 119600 546380
rect 119520 546310 119530 546370
rect 119590 546310 119600 546370
rect 124990 546360 125000 546400
rect 125040 546360 125050 546400
rect 124990 546340 125050 546360
rect 125090 546400 125170 546420
rect 125090 546360 125110 546400
rect 125150 546360 125170 546400
rect 125090 546350 125170 546360
rect 125210 546400 125270 546420
rect 125210 546360 125220 546400
rect 125260 546360 125270 546400
rect 125210 546340 125270 546360
rect 119520 546300 119600 546310
rect 119200 546260 119280 546270
rect 119200 546200 119210 546260
rect 119270 546200 119280 546260
rect 119530 546210 119590 546300
rect 119200 546190 119280 546200
rect 119360 546160 120350 546210
rect 119360 546060 119420 546160
rect 119640 546090 119680 546160
rect 119360 546010 119370 546060
rect 119410 546010 119420 546060
rect 119360 545990 119420 546010
rect 119470 546060 119530 546080
rect 119470 546010 119480 546060
rect 119520 546010 119530 546060
rect 119470 545860 119530 546010
rect 119640 545910 119680 545930
rect 119720 546090 119780 546110
rect 119720 545930 119730 546090
rect 119770 545930 119780 546090
rect 119570 545860 119650 545870
rect 119470 545850 119650 545860
rect 119470 545810 119590 545850
rect 119630 545810 119650 545850
rect 119360 545780 119420 545800
rect 119360 545730 119370 545780
rect 119410 545730 119420 545780
rect 119360 545710 119420 545730
rect 119470 545780 119530 545810
rect 119570 545790 119650 545810
rect 119470 545730 119480 545780
rect 119520 545730 119530 545780
rect 119470 545710 119530 545730
rect 119720 545700 119780 545930
rect 119640 545580 119680 545600
rect 119360 545350 119440 545360
rect 119640 545350 119680 545420
rect 119720 545580 119780 545640
rect 119720 545420 119730 545580
rect 119770 545420 119780 545580
rect 119720 545400 119780 545420
rect 119830 546090 119890 546110
rect 119830 545930 119840 546090
rect 119880 545930 119890 546090
rect 119830 545700 119890 545930
rect 120100 546090 120160 546110
rect 120100 545930 120110 546090
rect 120150 545930 120160 546090
rect 119950 545870 120030 545880
rect 119950 545810 119960 545870
rect 120020 545810 120030 545870
rect 119950 545800 120030 545810
rect 119950 545700 120030 545710
rect 120100 545700 120160 545930
rect 119830 545640 119960 545700
rect 120020 545640 120160 545700
rect 119830 545580 119890 545640
rect 119950 545630 120030 545640
rect 119830 545420 119840 545580
rect 119880 545420 119890 545580
rect 119830 545400 119890 545420
rect 120100 545580 120160 545640
rect 120100 545420 120110 545580
rect 120150 545420 120160 545580
rect 120100 545400 120160 545420
rect 120210 546090 120270 546110
rect 120210 545930 120220 546090
rect 120260 545930 120270 546090
rect 120210 545580 120270 545930
rect 120310 546090 120350 546160
rect 120310 545910 120350 545930
rect 120320 545860 120400 545870
rect 120320 545800 120330 545860
rect 120390 545800 120400 545860
rect 120320 545790 120400 545800
rect 120210 545420 120220 545580
rect 120260 545420 120270 545580
rect 120210 545350 120270 545420
rect 120310 545580 120350 545600
rect 120310 545350 120350 545420
rect 119350 545290 119370 545350
rect 119430 545290 120350 545350
rect 119360 545280 119440 545290
rect 125100 544940 125290 545070
rect 125430 544940 125890 545070
rect 126030 544940 126490 545070
rect 126730 544940 127190 545070
rect 127330 544940 127790 545070
rect 128030 544940 128490 545070
rect 128630 544940 129090 545070
rect 129330 544940 129790 545070
rect 129930 544940 130390 545070
rect 130630 544940 131090 545070
rect 131230 544940 131690 545070
rect 131930 544940 132390 545070
rect 132530 544940 132990 545070
rect 133230 544940 133690 545070
rect 133830 544940 134040 545070
rect 125100 544850 125240 544940
rect 133900 544890 134040 544940
rect 134030 544870 134040 544890
rect 125740 544850 125800 544870
rect 125740 544810 125750 544850
rect 125790 544810 125800 544850
rect 125740 544790 125800 544810
rect 126180 544850 126240 544870
rect 126180 544810 126190 544850
rect 126230 544810 126240 544850
rect 126180 544790 126240 544810
rect 126620 544850 126680 544870
rect 126620 544810 126630 544850
rect 126670 544810 126680 544850
rect 126620 544790 126680 544810
rect 127060 544850 127120 544870
rect 127060 544810 127070 544850
rect 127110 544810 127120 544850
rect 127060 544790 127120 544810
rect 127500 544850 127560 544870
rect 127500 544810 127510 544850
rect 127550 544810 127560 544850
rect 127500 544790 127560 544810
rect 127940 544850 128000 544870
rect 127940 544810 127950 544850
rect 127990 544810 128000 544850
rect 127940 544790 128000 544810
rect 128380 544850 128440 544870
rect 128380 544810 128390 544850
rect 128430 544810 128440 544850
rect 128380 544790 128440 544810
rect 128820 544850 128880 544870
rect 128820 544810 128830 544850
rect 128870 544810 128880 544850
rect 128820 544790 128880 544810
rect 129260 544850 129320 544870
rect 129260 544810 129270 544850
rect 129310 544810 129320 544850
rect 129260 544790 129320 544810
rect 129700 544850 129760 544870
rect 129700 544810 129710 544850
rect 129750 544810 129760 544850
rect 129700 544790 129760 544810
rect 130140 544850 130200 544870
rect 130140 544810 130150 544850
rect 130190 544810 130200 544850
rect 130140 544790 130200 544810
rect 130580 544850 130640 544870
rect 130580 544810 130590 544850
rect 130630 544810 130640 544850
rect 130580 544790 130640 544810
rect 131020 544850 131080 544870
rect 131020 544810 131030 544850
rect 131070 544810 131080 544850
rect 131020 544790 131080 544810
rect 131460 544850 131520 544870
rect 131460 544810 131470 544850
rect 131510 544810 131520 544850
rect 131460 544790 131520 544810
rect 131900 544850 131960 544870
rect 131900 544810 131910 544850
rect 131950 544810 131960 544850
rect 131900 544790 131960 544810
rect 132340 544850 132400 544870
rect 132340 544810 132350 544850
rect 132390 544810 132400 544850
rect 132340 544790 132400 544810
rect 132780 544850 132840 544870
rect 132780 544810 132790 544850
rect 132830 544810 132840 544850
rect 132780 544790 132840 544810
rect 133220 544850 133280 544870
rect 133220 544810 133230 544850
rect 133270 544810 133280 544850
rect 133220 544790 133280 544810
rect 133660 544850 133720 544870
rect 133660 544810 133670 544850
rect 133710 544810 133720 544850
rect 133660 544790 133720 544810
rect 125100 544290 125240 544720
rect 125480 544650 125540 544670
rect 125480 544410 125490 544650
rect 125530 544410 125540 544650
rect 125480 544390 125540 544410
rect 125580 544650 125760 544670
rect 125580 544410 125600 544650
rect 125740 544410 125760 544650
rect 125580 544400 125760 544410
rect 125800 544650 125860 544670
rect 125800 544410 125810 544650
rect 125850 544410 125860 544650
rect 125800 544390 125860 544410
rect 125920 544650 125980 544670
rect 125920 544410 125930 544650
rect 125970 544410 125980 544650
rect 125920 544390 125980 544410
rect 126020 544650 126200 544670
rect 126020 544410 126040 544650
rect 126180 544410 126200 544650
rect 126020 544400 126200 544410
rect 126240 544650 126300 544670
rect 126240 544410 126250 544650
rect 126290 544410 126300 544650
rect 126240 544390 126300 544410
rect 126360 544650 126420 544670
rect 126360 544410 126370 544650
rect 126410 544410 126420 544650
rect 126360 544390 126420 544410
rect 126460 544650 126640 544670
rect 126460 544410 126480 544650
rect 126620 544410 126640 544650
rect 126460 544400 126640 544410
rect 126680 544650 126740 544670
rect 126680 544410 126690 544650
rect 126730 544410 126740 544650
rect 126680 544390 126740 544410
rect 126800 544650 126860 544670
rect 126800 544410 126810 544650
rect 126850 544410 126860 544650
rect 126800 544390 126860 544410
rect 126900 544650 127080 544670
rect 126900 544410 126920 544650
rect 127060 544410 127080 544650
rect 126900 544400 127080 544410
rect 127120 544650 127180 544670
rect 127120 544410 127130 544650
rect 127170 544410 127180 544650
rect 127120 544390 127180 544410
rect 127240 544650 127300 544670
rect 127240 544410 127250 544650
rect 127290 544410 127300 544650
rect 127240 544390 127300 544410
rect 127340 544650 127520 544670
rect 127340 544410 127360 544650
rect 127500 544410 127520 544650
rect 127340 544400 127520 544410
rect 127560 544650 127620 544670
rect 127560 544410 127570 544650
rect 127610 544410 127620 544650
rect 127560 544390 127620 544410
rect 127680 544650 127740 544670
rect 127680 544410 127690 544650
rect 127730 544410 127740 544650
rect 127680 544390 127740 544410
rect 127780 544650 127960 544670
rect 127780 544410 127800 544650
rect 127940 544410 127960 544650
rect 127780 544400 127960 544410
rect 128000 544650 128060 544670
rect 128000 544410 128010 544650
rect 128050 544410 128060 544650
rect 128000 544390 128060 544410
rect 128120 544650 128180 544670
rect 128120 544410 128130 544650
rect 128170 544410 128180 544650
rect 128120 544390 128180 544410
rect 128220 544650 128400 544670
rect 128220 544410 128240 544650
rect 128380 544410 128400 544650
rect 128220 544400 128400 544410
rect 128440 544650 128500 544670
rect 128440 544410 128450 544650
rect 128490 544410 128500 544650
rect 128440 544390 128500 544410
rect 128560 544650 128620 544670
rect 128560 544410 128570 544650
rect 128610 544410 128620 544650
rect 128560 544390 128620 544410
rect 128660 544650 128840 544670
rect 128660 544410 128680 544650
rect 128820 544410 128840 544650
rect 128660 544400 128840 544410
rect 128880 544650 128940 544670
rect 128880 544410 128890 544650
rect 128930 544410 128940 544650
rect 128880 544390 128940 544410
rect 129000 544650 129060 544670
rect 129000 544410 129010 544650
rect 129050 544410 129060 544650
rect 129000 544390 129060 544410
rect 129100 544650 129280 544670
rect 129100 544410 129120 544650
rect 129260 544410 129280 544650
rect 129100 544400 129280 544410
rect 129320 544650 129380 544670
rect 129320 544410 129330 544650
rect 129370 544410 129380 544650
rect 129320 544390 129380 544410
rect 129440 544650 129500 544670
rect 129440 544410 129450 544650
rect 129490 544410 129500 544650
rect 129440 544390 129500 544410
rect 129540 544650 129720 544670
rect 129540 544410 129560 544650
rect 129700 544410 129720 544650
rect 129540 544400 129720 544410
rect 129760 544650 129820 544670
rect 129760 544410 129770 544650
rect 129810 544410 129820 544650
rect 129760 544390 129820 544410
rect 129880 544650 129940 544670
rect 129880 544410 129890 544650
rect 129930 544410 129940 544650
rect 129880 544390 129940 544410
rect 129980 544650 130160 544670
rect 129980 544410 130000 544650
rect 130140 544410 130160 544650
rect 129980 544400 130160 544410
rect 130200 544650 130260 544670
rect 130200 544410 130210 544650
rect 130250 544410 130260 544650
rect 130200 544390 130260 544410
rect 130320 544650 130380 544670
rect 130320 544410 130330 544650
rect 130370 544410 130380 544650
rect 130320 544390 130380 544410
rect 130420 544650 130600 544670
rect 130420 544410 130440 544650
rect 130580 544410 130600 544650
rect 130420 544400 130600 544410
rect 130640 544650 130700 544670
rect 130640 544410 130650 544650
rect 130690 544410 130700 544650
rect 130640 544390 130700 544410
rect 130760 544650 130820 544670
rect 130760 544410 130770 544650
rect 130810 544410 130820 544650
rect 130760 544390 130820 544410
rect 130860 544650 131040 544670
rect 130860 544410 130880 544650
rect 131020 544410 131040 544650
rect 130860 544400 131040 544410
rect 131080 544650 131140 544670
rect 131080 544410 131090 544650
rect 131130 544410 131140 544650
rect 131080 544390 131140 544410
rect 131200 544650 131260 544670
rect 131200 544410 131210 544650
rect 131250 544410 131260 544650
rect 131200 544390 131260 544410
rect 131300 544650 131480 544670
rect 131300 544410 131320 544650
rect 131460 544410 131480 544650
rect 131300 544400 131480 544410
rect 131520 544650 131580 544670
rect 131520 544410 131530 544650
rect 131570 544410 131580 544650
rect 131520 544390 131580 544410
rect 131640 544650 131700 544670
rect 131640 544410 131650 544650
rect 131690 544410 131700 544650
rect 131640 544390 131700 544410
rect 131740 544650 131920 544670
rect 131740 544410 131760 544650
rect 131900 544410 131920 544650
rect 131740 544400 131920 544410
rect 131960 544650 132020 544670
rect 131960 544410 131970 544650
rect 132010 544410 132020 544650
rect 131960 544390 132020 544410
rect 132080 544650 132140 544670
rect 132080 544410 132090 544650
rect 132130 544410 132140 544650
rect 132080 544390 132140 544410
rect 132180 544650 132360 544670
rect 132180 544410 132200 544650
rect 132340 544410 132360 544650
rect 132180 544400 132360 544410
rect 132400 544650 132460 544670
rect 132400 544410 132410 544650
rect 132450 544410 132460 544650
rect 132400 544390 132460 544410
rect 132520 544650 132580 544670
rect 132520 544410 132530 544650
rect 132570 544410 132580 544650
rect 132520 544390 132580 544410
rect 132620 544650 132800 544670
rect 132620 544410 132640 544650
rect 132780 544410 132800 544650
rect 132620 544400 132800 544410
rect 132840 544650 132900 544670
rect 132840 544410 132850 544650
rect 132890 544410 132900 544650
rect 132840 544390 132900 544410
rect 132960 544650 133020 544670
rect 132960 544410 132970 544650
rect 133010 544410 133020 544650
rect 132960 544390 133020 544410
rect 133060 544650 133240 544670
rect 133060 544410 133080 544650
rect 133220 544410 133240 544650
rect 133060 544400 133240 544410
rect 133280 544650 133340 544670
rect 133280 544410 133290 544650
rect 133330 544410 133340 544650
rect 133280 544390 133340 544410
rect 133400 544650 133460 544670
rect 133400 544410 133410 544650
rect 133450 544410 133460 544650
rect 133400 544390 133460 544410
rect 133500 544650 133680 544670
rect 133500 544410 133520 544650
rect 133660 544410 133680 544650
rect 133500 544400 133680 544410
rect 133720 544650 133780 544670
rect 133720 544410 133730 544650
rect 133770 544410 133780 544650
rect 133720 544390 133780 544410
rect 125100 544070 125240 544160
rect 134030 544300 134040 544740
rect 134030 544120 134040 544170
rect 133900 544070 134040 544120
rect 125100 543940 125290 544070
rect 125430 543940 125890 544070
rect 126030 543940 126490 544070
rect 126730 543940 127190 544070
rect 127330 543940 127790 544070
rect 128030 543940 128490 544070
rect 128630 543940 129090 544070
rect 129330 543940 129790 544070
rect 129930 543940 130390 544070
rect 130630 543940 131090 544070
rect 131230 543940 131690 544070
rect 131930 543940 132390 544070
rect 132530 543940 132990 544070
rect 133230 543940 133690 544070
rect 133830 543940 134040 544070
rect 125120 538540 125180 538560
rect 125120 538500 125130 538540
rect 125170 538500 125180 538540
rect 125120 538480 125180 538500
rect 124960 538340 125020 538360
rect 119500 538320 119560 538330
rect 119490 538310 119570 538320
rect 119490 538250 119500 538310
rect 119560 538250 119570 538310
rect 124960 538300 124970 538340
rect 125010 538300 125020 538340
rect 124960 538280 125020 538300
rect 125060 538340 125140 538360
rect 125060 538300 125080 538340
rect 125120 538300 125140 538340
rect 125060 538290 125140 538300
rect 125180 538340 125240 538360
rect 125180 538300 125190 538340
rect 125230 538300 125240 538340
rect 125180 538280 125240 538300
rect 119490 538240 119570 538250
rect 119170 538200 119250 538210
rect 119170 538140 119180 538200
rect 119240 538140 119250 538200
rect 119500 538150 119560 538240
rect 119170 538130 119250 538140
rect 119330 538100 120320 538150
rect 119330 538000 119390 538100
rect 119610 538030 119650 538100
rect 119330 537950 119340 538000
rect 119380 537950 119390 538000
rect 119330 537930 119390 537950
rect 119440 538000 119500 538020
rect 119440 537950 119450 538000
rect 119490 537950 119500 538000
rect 119440 537800 119500 537950
rect 119610 537850 119650 537870
rect 119690 538030 119750 538050
rect 119690 537870 119700 538030
rect 119740 537870 119750 538030
rect 119540 537800 119620 537810
rect 119440 537790 119620 537800
rect 119440 537750 119560 537790
rect 119600 537750 119620 537790
rect 119330 537720 119390 537740
rect 119330 537670 119340 537720
rect 119380 537670 119390 537720
rect 119330 537650 119390 537670
rect 119440 537720 119500 537750
rect 119540 537730 119620 537750
rect 119440 537670 119450 537720
rect 119490 537670 119500 537720
rect 119440 537650 119500 537670
rect 119690 537640 119750 537870
rect 119610 537520 119650 537540
rect 119330 537290 119410 537300
rect 119610 537290 119650 537360
rect 119690 537520 119750 537580
rect 119690 537360 119700 537520
rect 119740 537360 119750 537520
rect 119690 537340 119750 537360
rect 119800 538030 119860 538050
rect 119800 537870 119810 538030
rect 119850 537870 119860 538030
rect 119800 537640 119860 537870
rect 120070 538030 120130 538050
rect 120070 537870 120080 538030
rect 120120 537870 120130 538030
rect 119920 537810 120000 537820
rect 119920 537750 119930 537810
rect 119990 537750 120000 537810
rect 119920 537740 120000 537750
rect 119920 537640 120000 537650
rect 120070 537640 120130 537870
rect 119800 537580 119930 537640
rect 119990 537580 120130 537640
rect 119800 537520 119860 537580
rect 119920 537570 120000 537580
rect 119800 537360 119810 537520
rect 119850 537360 119860 537520
rect 119800 537340 119860 537360
rect 120070 537520 120130 537580
rect 120070 537360 120080 537520
rect 120120 537360 120130 537520
rect 120070 537340 120130 537360
rect 120180 538030 120240 538050
rect 120180 537870 120190 538030
rect 120230 537870 120240 538030
rect 120180 537520 120240 537870
rect 120280 538030 120320 538100
rect 120280 537850 120320 537870
rect 120290 537800 120370 537810
rect 120290 537740 120300 537800
rect 120360 537740 120370 537800
rect 120290 537730 120370 537740
rect 120180 537360 120190 537520
rect 120230 537360 120240 537520
rect 120180 537290 120240 537360
rect 120280 537520 120320 537540
rect 120280 537290 120320 537360
rect 119320 537230 119340 537290
rect 119400 537230 120320 537290
rect 119330 537220 119410 537230
rect 125070 536880 125260 537010
rect 125400 536880 125860 537010
rect 126000 536880 126460 537010
rect 126700 536880 127160 537010
rect 127300 536880 127760 537010
rect 128000 536880 128460 537010
rect 128600 536880 129060 537010
rect 129300 536880 129760 537010
rect 129900 536880 130360 537010
rect 130600 536880 131060 537010
rect 131200 536880 131660 537010
rect 131900 536880 132360 537010
rect 132500 536880 132960 537010
rect 133200 536880 133660 537010
rect 133800 536880 134010 537010
rect 125070 536790 125210 536880
rect 133870 536830 134010 536880
rect 134000 536810 134010 536830
rect 125710 536790 125770 536810
rect 125710 536750 125720 536790
rect 125760 536750 125770 536790
rect 125710 536730 125770 536750
rect 126150 536790 126210 536810
rect 126150 536750 126160 536790
rect 126200 536750 126210 536790
rect 126150 536730 126210 536750
rect 126590 536790 126650 536810
rect 126590 536750 126600 536790
rect 126640 536750 126650 536790
rect 126590 536730 126650 536750
rect 127030 536790 127090 536810
rect 127030 536750 127040 536790
rect 127080 536750 127090 536790
rect 127030 536730 127090 536750
rect 127470 536790 127530 536810
rect 127470 536750 127480 536790
rect 127520 536750 127530 536790
rect 127470 536730 127530 536750
rect 127910 536790 127970 536810
rect 127910 536750 127920 536790
rect 127960 536750 127970 536790
rect 127910 536730 127970 536750
rect 128350 536790 128410 536810
rect 128350 536750 128360 536790
rect 128400 536750 128410 536790
rect 128350 536730 128410 536750
rect 128790 536790 128850 536810
rect 128790 536750 128800 536790
rect 128840 536750 128850 536790
rect 128790 536730 128850 536750
rect 129230 536790 129290 536810
rect 129230 536750 129240 536790
rect 129280 536750 129290 536790
rect 129230 536730 129290 536750
rect 129670 536790 129730 536810
rect 129670 536750 129680 536790
rect 129720 536750 129730 536790
rect 129670 536730 129730 536750
rect 130110 536790 130170 536810
rect 130110 536750 130120 536790
rect 130160 536750 130170 536790
rect 130110 536730 130170 536750
rect 130550 536790 130610 536810
rect 130550 536750 130560 536790
rect 130600 536750 130610 536790
rect 130550 536730 130610 536750
rect 130990 536790 131050 536810
rect 130990 536750 131000 536790
rect 131040 536750 131050 536790
rect 130990 536730 131050 536750
rect 131430 536790 131490 536810
rect 131430 536750 131440 536790
rect 131480 536750 131490 536790
rect 131430 536730 131490 536750
rect 131870 536790 131930 536810
rect 131870 536750 131880 536790
rect 131920 536750 131930 536790
rect 131870 536730 131930 536750
rect 132310 536790 132370 536810
rect 132310 536750 132320 536790
rect 132360 536750 132370 536790
rect 132310 536730 132370 536750
rect 132750 536790 132810 536810
rect 132750 536750 132760 536790
rect 132800 536750 132810 536790
rect 132750 536730 132810 536750
rect 133190 536790 133250 536810
rect 133190 536750 133200 536790
rect 133240 536750 133250 536790
rect 133190 536730 133250 536750
rect 133630 536790 133690 536810
rect 133630 536750 133640 536790
rect 133680 536750 133690 536790
rect 133630 536730 133690 536750
rect 125070 536030 125210 536660
rect 125450 536590 125510 536610
rect 125450 536150 125460 536590
rect 125500 536150 125510 536590
rect 125450 536130 125510 536150
rect 125550 536590 125730 536610
rect 125550 536150 125570 536590
rect 125710 536150 125730 536590
rect 125550 536140 125730 536150
rect 125770 536590 125830 536610
rect 125770 536150 125780 536590
rect 125820 536150 125830 536590
rect 125770 536130 125830 536150
rect 125890 536590 125950 536610
rect 125890 536150 125900 536590
rect 125940 536150 125950 536590
rect 125890 536130 125950 536150
rect 125990 536590 126170 536610
rect 125990 536150 126010 536590
rect 126150 536150 126170 536590
rect 125990 536140 126170 536150
rect 126210 536590 126270 536610
rect 126210 536150 126220 536590
rect 126260 536150 126270 536590
rect 126210 536130 126270 536150
rect 126330 536590 126390 536610
rect 126330 536150 126340 536590
rect 126380 536150 126390 536590
rect 126330 536130 126390 536150
rect 126430 536590 126610 536610
rect 126430 536150 126450 536590
rect 126590 536150 126610 536590
rect 126430 536140 126610 536150
rect 126650 536590 126710 536610
rect 126650 536150 126660 536590
rect 126700 536150 126710 536590
rect 126650 536130 126710 536150
rect 126770 536590 126830 536610
rect 126770 536150 126780 536590
rect 126820 536150 126830 536590
rect 126770 536130 126830 536150
rect 126870 536590 127050 536610
rect 126870 536150 126890 536590
rect 127030 536150 127050 536590
rect 126870 536140 127050 536150
rect 127090 536590 127150 536610
rect 127090 536150 127100 536590
rect 127140 536150 127150 536590
rect 127090 536130 127150 536150
rect 127210 536590 127270 536610
rect 127210 536150 127220 536590
rect 127260 536150 127270 536590
rect 127210 536130 127270 536150
rect 127310 536590 127490 536610
rect 127310 536150 127330 536590
rect 127470 536150 127490 536590
rect 127310 536140 127490 536150
rect 127530 536590 127590 536610
rect 127530 536150 127540 536590
rect 127580 536150 127590 536590
rect 127530 536130 127590 536150
rect 127650 536590 127710 536610
rect 127650 536150 127660 536590
rect 127700 536150 127710 536590
rect 127650 536130 127710 536150
rect 127750 536590 127930 536610
rect 127750 536150 127770 536590
rect 127910 536150 127930 536590
rect 127750 536140 127930 536150
rect 127970 536590 128030 536610
rect 127970 536150 127980 536590
rect 128020 536150 128030 536590
rect 127970 536130 128030 536150
rect 128090 536590 128150 536610
rect 128090 536150 128100 536590
rect 128140 536150 128150 536590
rect 128090 536130 128150 536150
rect 128190 536590 128370 536610
rect 128190 536150 128210 536590
rect 128350 536150 128370 536590
rect 128190 536140 128370 536150
rect 128410 536590 128470 536610
rect 128410 536150 128420 536590
rect 128460 536150 128470 536590
rect 128410 536130 128470 536150
rect 128530 536590 128590 536610
rect 128530 536150 128540 536590
rect 128580 536150 128590 536590
rect 128530 536130 128590 536150
rect 128630 536590 128810 536610
rect 128630 536150 128650 536590
rect 128790 536150 128810 536590
rect 128630 536140 128810 536150
rect 128850 536590 128910 536610
rect 128850 536150 128860 536590
rect 128900 536150 128910 536590
rect 128850 536130 128910 536150
rect 128970 536590 129030 536610
rect 128970 536150 128980 536590
rect 129020 536150 129030 536590
rect 128970 536130 129030 536150
rect 129070 536590 129250 536610
rect 129070 536150 129090 536590
rect 129230 536150 129250 536590
rect 129070 536140 129250 536150
rect 129290 536590 129350 536610
rect 129290 536150 129300 536590
rect 129340 536150 129350 536590
rect 129290 536130 129350 536150
rect 129410 536590 129470 536610
rect 129410 536150 129420 536590
rect 129460 536150 129470 536590
rect 129410 536130 129470 536150
rect 129510 536590 129690 536610
rect 129510 536150 129530 536590
rect 129670 536150 129690 536590
rect 129510 536140 129690 536150
rect 129730 536590 129790 536610
rect 129730 536150 129740 536590
rect 129780 536150 129790 536590
rect 129730 536130 129790 536150
rect 129850 536590 129910 536610
rect 129850 536150 129860 536590
rect 129900 536150 129910 536590
rect 129850 536130 129910 536150
rect 129950 536590 130130 536610
rect 129950 536150 129970 536590
rect 130110 536150 130130 536590
rect 129950 536140 130130 536150
rect 130170 536590 130230 536610
rect 130170 536150 130180 536590
rect 130220 536150 130230 536590
rect 130170 536130 130230 536150
rect 130290 536590 130350 536610
rect 130290 536150 130300 536590
rect 130340 536150 130350 536590
rect 130290 536130 130350 536150
rect 130390 536590 130570 536610
rect 130390 536150 130410 536590
rect 130550 536150 130570 536590
rect 130390 536140 130570 536150
rect 130610 536590 130670 536610
rect 130610 536150 130620 536590
rect 130660 536150 130670 536590
rect 130610 536130 130670 536150
rect 130730 536590 130790 536610
rect 130730 536150 130740 536590
rect 130780 536150 130790 536590
rect 130730 536130 130790 536150
rect 130830 536590 131010 536610
rect 130830 536150 130850 536590
rect 130990 536150 131010 536590
rect 130830 536140 131010 536150
rect 131050 536590 131110 536610
rect 131050 536150 131060 536590
rect 131100 536150 131110 536590
rect 131050 536130 131110 536150
rect 131170 536590 131230 536610
rect 131170 536150 131180 536590
rect 131220 536150 131230 536590
rect 131170 536130 131230 536150
rect 131270 536590 131450 536610
rect 131270 536150 131290 536590
rect 131430 536150 131450 536590
rect 131270 536140 131450 536150
rect 131490 536590 131550 536610
rect 131490 536150 131500 536590
rect 131540 536150 131550 536590
rect 131490 536130 131550 536150
rect 131610 536590 131670 536610
rect 131610 536150 131620 536590
rect 131660 536150 131670 536590
rect 131610 536130 131670 536150
rect 131710 536590 131890 536610
rect 131710 536150 131730 536590
rect 131870 536150 131890 536590
rect 131710 536140 131890 536150
rect 131930 536590 131990 536610
rect 131930 536150 131940 536590
rect 131980 536150 131990 536590
rect 131930 536130 131990 536150
rect 132050 536590 132110 536610
rect 132050 536150 132060 536590
rect 132100 536150 132110 536590
rect 132050 536130 132110 536150
rect 132150 536590 132330 536610
rect 132150 536150 132170 536590
rect 132310 536150 132330 536590
rect 132150 536140 132330 536150
rect 132370 536590 132430 536610
rect 132370 536150 132380 536590
rect 132420 536150 132430 536590
rect 132370 536130 132430 536150
rect 132490 536590 132550 536610
rect 132490 536150 132500 536590
rect 132540 536150 132550 536590
rect 132490 536130 132550 536150
rect 132590 536590 132770 536610
rect 132590 536150 132610 536590
rect 132750 536150 132770 536590
rect 132590 536140 132770 536150
rect 132810 536590 132870 536610
rect 132810 536150 132820 536590
rect 132860 536150 132870 536590
rect 132810 536130 132870 536150
rect 132930 536590 132990 536610
rect 132930 536150 132940 536590
rect 132980 536150 132990 536590
rect 132930 536130 132990 536150
rect 133030 536590 133210 536610
rect 133030 536150 133050 536590
rect 133190 536150 133210 536590
rect 133030 536140 133210 536150
rect 133250 536590 133310 536610
rect 133250 536150 133260 536590
rect 133300 536150 133310 536590
rect 133250 536130 133310 536150
rect 133370 536590 133430 536610
rect 133370 536150 133380 536590
rect 133420 536150 133430 536590
rect 133370 536130 133430 536150
rect 133470 536590 133650 536610
rect 133470 536150 133490 536590
rect 133630 536150 133650 536590
rect 133470 536140 133650 536150
rect 133690 536590 133750 536610
rect 133690 536150 133700 536590
rect 133740 536150 133750 536590
rect 133690 536130 133750 536150
rect 125070 535810 125210 535900
rect 134000 536040 134010 536680
rect 134000 535860 134010 535910
rect 133870 535810 134010 535860
rect 125070 535680 125260 535810
rect 125400 535680 125860 535810
rect 126000 535680 126460 535810
rect 126700 535680 127160 535810
rect 127300 535680 127760 535810
rect 128000 535680 128460 535810
rect 128600 535680 129060 535810
rect 129300 535680 129760 535810
rect 129900 535680 130360 535810
rect 130600 535680 131060 535810
rect 131200 535680 131660 535810
rect 131900 535680 132360 535810
rect 132500 535680 132960 535810
rect 133200 535680 133660 535810
rect 133800 535680 134010 535810
<< viali >>
rect 124040 642710 124080 642750
rect 123830 642040 123960 642610
rect 124170 642450 124220 642500
rect 124350 642450 124400 642500
rect 124530 642450 124580 642500
rect 124710 642450 124760 642500
rect 124890 642450 124940 642500
rect 125070 642450 125120 642500
rect 125250 642450 125300 642500
rect 125430 642450 125480 642500
rect 125610 642450 125660 642500
rect 125790 642450 125840 642500
rect 125970 642450 126020 642500
rect 126150 642450 126200 642500
rect 126330 642450 126380 642500
rect 126510 642450 126560 642500
rect 126690 642450 126740 642500
rect 126870 642450 126920 642500
rect 127050 642450 127100 642500
rect 127230 642450 127280 642500
rect 127410 642450 127460 642500
rect 127590 642450 127640 642500
rect 127770 642450 127820 642500
rect 127950 642450 128000 642500
rect 128130 642450 128180 642500
rect 128310 642450 128360 642500
rect 128490 642450 128540 642500
rect 128670 642450 128720 642500
rect 128850 642450 128900 642500
rect 129030 642450 129080 642500
rect 129210 642450 129260 642500
rect 129390 642450 129440 642500
rect 129570 642450 129620 642500
rect 129750 642450 129800 642500
rect 129930 642450 129980 642500
rect 130110 642450 130160 642500
rect 130290 642450 130340 642500
rect 130470 642450 130520 642500
rect 130650 642450 130700 642500
rect 130830 642450 130880 642500
rect 131010 642450 131060 642500
rect 131190 642450 131240 642500
rect 124170 642150 124220 642200
rect 124350 642150 124400 642200
rect 124530 642150 124580 642200
rect 124710 642150 124760 642200
rect 124890 642150 124940 642200
rect 125070 642150 125120 642200
rect 125250 642150 125300 642200
rect 125430 642150 125480 642200
rect 125610 642150 125660 642200
rect 125790 642150 125840 642200
rect 125970 642150 126020 642200
rect 126150 642150 126200 642200
rect 126330 642150 126380 642200
rect 126510 642150 126560 642200
rect 126690 642150 126740 642200
rect 126870 642150 126920 642200
rect 127050 642150 127100 642200
rect 127230 642150 127280 642200
rect 127410 642150 127460 642200
rect 127590 642150 127640 642200
rect 127770 642150 127820 642200
rect 127950 642150 128000 642200
rect 128130 642150 128180 642200
rect 128310 642150 128360 642200
rect 128490 642150 128540 642200
rect 128670 642150 128720 642200
rect 128850 642150 128900 642200
rect 129030 642150 129080 642200
rect 129210 642150 129260 642200
rect 129390 642150 129440 642200
rect 129570 642150 129620 642200
rect 129750 642150 129800 642200
rect 129930 642150 129980 642200
rect 130110 642150 130160 642200
rect 130290 642150 130340 642200
rect 130470 642150 130520 642200
rect 130650 642150 130700 642200
rect 130830 642150 130880 642200
rect 131010 642150 131060 642200
rect 131190 642150 131240 642200
rect 131500 642060 131630 642630
rect 124200 636280 124340 636330
rect 124440 636280 124580 636330
rect 124680 636280 124820 636330
rect 124920 636280 125060 636330
rect 125160 636280 125300 636330
rect 125400 636280 125540 636330
rect 125640 636280 125780 636330
rect 125880 636280 126020 636330
rect 126120 636280 126260 636330
rect 126360 636280 126500 636330
rect 126600 636280 126740 636330
rect 126840 636280 126980 636330
rect 127080 636280 127220 636330
rect 127320 636280 127460 636330
rect 127560 636280 127700 636330
rect 127800 636280 127940 636330
rect 128040 636280 128180 636330
rect 128280 636280 128420 636330
rect 128520 636280 128660 636330
rect 128760 636280 128900 636330
rect 124070 636130 124110 636170
rect 124200 635980 124340 636030
rect 124440 635980 124580 636030
rect 124680 635980 124820 636030
rect 124920 635980 125060 636030
rect 125160 635980 125300 636030
rect 125400 635980 125540 636030
rect 125640 635980 125780 636030
rect 125880 635980 126020 636030
rect 126120 635980 126260 636030
rect 126360 635980 126500 636030
rect 126600 635980 126740 636030
rect 126840 635980 126980 636030
rect 127080 635980 127220 636030
rect 127320 635980 127460 636030
rect 127560 635980 127700 636030
rect 127800 635980 127940 636030
rect 128040 635980 128180 636030
rect 128280 635980 128420 636030
rect 128520 635980 128660 636030
rect 128760 635980 128900 636030
rect 129100 635900 129230 636470
rect 124260 632690 124620 632740
rect 124260 632390 124620 632440
rect 124470 630250 124830 630300
rect 124930 630250 125290 630300
rect 125390 630250 125750 630300
rect 125850 630250 126210 630300
rect 126310 630250 126670 630300
rect 126770 630250 127130 630300
rect 127230 630250 127590 630300
rect 127690 630250 128050 630300
rect 128150 630250 128510 630300
rect 128610 630250 128970 630300
rect 124350 630100 124390 630140
rect 124470 629950 124830 630000
rect 124930 629950 125290 630000
rect 125390 629950 125750 630000
rect 125850 629950 126210 630000
rect 126310 629950 126670 630000
rect 126770 629950 127130 630000
rect 127230 629950 127590 630000
rect 127690 629950 128050 630000
rect 128150 629950 128510 630000
rect 128610 629950 128970 630000
rect 129170 629840 129300 630410
rect 124240 625020 124800 625070
rect 124240 624720 124800 624770
rect 124600 623970 124640 624010
rect 124800 623730 125360 623780
rect 125460 623730 126020 623780
rect 126120 623730 126680 623780
rect 126780 623730 127340 623780
rect 127440 623730 128000 623780
rect 128100 623730 128660 623780
rect 124800 623430 125360 623480
rect 125460 623430 126020 623480
rect 126120 623430 126680 623480
rect 126780 623430 127340 623480
rect 127440 623430 128000 623480
rect 128100 623430 128660 623480
rect 128820 623320 128950 623890
rect 125360 619310 125400 619350
rect 125470 619310 125510 619350
rect 125580 619310 125620 619350
rect 131940 618790 132070 618810
rect 125590 618730 125630 618770
rect 125930 618730 125970 618770
rect 126270 618730 126310 618770
rect 126610 618730 126650 618770
rect 126950 618730 126990 618770
rect 127290 618730 127330 618770
rect 127630 618730 127670 618770
rect 127970 618730 128010 618770
rect 128310 618730 128350 618770
rect 128650 618730 128690 618770
rect 128990 618730 129030 618770
rect 129330 618730 129370 618770
rect 129670 618730 129710 618770
rect 130010 618730 130050 618770
rect 130350 618730 130390 618770
rect 130690 618730 130730 618770
rect 131030 618730 131070 618770
rect 131370 618730 131410 618770
rect 131710 618730 131750 618770
rect 131940 618660 132070 618790
rect 125430 618530 125470 618570
rect 125540 618530 125580 618570
rect 125650 618530 125690 618570
rect 125770 618530 125810 618570
rect 125880 618530 125920 618570
rect 125990 618530 126030 618570
rect 126110 618530 126150 618570
rect 126220 618530 126260 618570
rect 126330 618530 126370 618570
rect 126450 618530 126490 618570
rect 126560 618530 126600 618570
rect 126670 618530 126710 618570
rect 126790 618530 126830 618570
rect 126900 618530 126940 618570
rect 127010 618530 127050 618570
rect 127130 618530 127170 618570
rect 127240 618530 127280 618570
rect 127350 618530 127390 618570
rect 127470 618530 127510 618570
rect 127580 618530 127620 618570
rect 127690 618530 127730 618570
rect 127810 618530 127850 618570
rect 127920 618530 127960 618570
rect 128030 618530 128070 618570
rect 128150 618530 128190 618570
rect 128260 618530 128300 618570
rect 128370 618530 128410 618570
rect 128490 618530 128530 618570
rect 128600 618530 128640 618570
rect 128710 618530 128750 618570
rect 128830 618530 128870 618570
rect 128940 618530 128980 618570
rect 129050 618530 129090 618570
rect 129170 618530 129210 618570
rect 129280 618530 129320 618570
rect 129390 618530 129430 618570
rect 129510 618530 129550 618570
rect 129620 618530 129660 618570
rect 129730 618530 129770 618570
rect 129850 618530 129890 618570
rect 129960 618530 130000 618570
rect 130070 618530 130110 618570
rect 130190 618530 130230 618570
rect 130300 618530 130340 618570
rect 130410 618530 130450 618570
rect 130530 618530 130570 618570
rect 130640 618530 130680 618570
rect 130750 618530 130790 618570
rect 130870 618530 130910 618570
rect 130980 618530 131020 618570
rect 131090 618530 131130 618570
rect 131210 618530 131250 618570
rect 131320 618530 131360 618570
rect 131430 618530 131470 618570
rect 131550 618530 131590 618570
rect 131660 618530 131700 618570
rect 131770 618530 131810 618570
rect 131940 618420 132070 618660
rect 131940 618290 132070 618420
rect 131940 618240 132070 618290
rect 125010 611860 125050 611900
rect 125120 611860 125160 611900
rect 125230 611860 125270 611900
rect 131590 611340 131720 611360
rect 125240 611280 125280 611320
rect 125580 611280 125620 611320
rect 125920 611280 125960 611320
rect 126260 611280 126300 611320
rect 126600 611280 126640 611320
rect 126940 611280 126980 611320
rect 127280 611280 127320 611320
rect 127620 611280 127660 611320
rect 127960 611280 128000 611320
rect 128300 611280 128340 611320
rect 128640 611280 128680 611320
rect 128980 611280 129020 611320
rect 129320 611280 129360 611320
rect 129660 611280 129700 611320
rect 130000 611280 130040 611320
rect 130340 611280 130380 611320
rect 130680 611280 130720 611320
rect 131020 611280 131060 611320
rect 131360 611280 131400 611320
rect 131590 611210 131720 611340
rect 125080 610930 125120 611120
rect 125190 610930 125230 611120
rect 125300 610930 125340 611120
rect 125420 610930 125460 611120
rect 125530 610930 125570 611120
rect 125640 610930 125680 611120
rect 125760 610930 125800 611120
rect 125870 610930 125910 611120
rect 125980 610930 126020 611120
rect 126100 610930 126140 611120
rect 126210 610930 126250 611120
rect 126320 610930 126360 611120
rect 126440 610930 126480 611120
rect 126550 610930 126590 611120
rect 126660 610930 126700 611120
rect 126780 610930 126820 611120
rect 126890 610930 126930 611120
rect 127000 610930 127040 611120
rect 127120 610930 127160 611120
rect 127230 610930 127270 611120
rect 127340 610930 127380 611120
rect 127460 610930 127500 611120
rect 127570 610930 127610 611120
rect 127680 610930 127720 611120
rect 127800 610930 127840 611120
rect 127910 610930 127950 611120
rect 128020 610930 128060 611120
rect 128140 610930 128180 611120
rect 128250 610930 128290 611120
rect 128360 610930 128400 611120
rect 128480 610930 128520 611120
rect 128590 610930 128630 611120
rect 128700 610930 128740 611120
rect 128820 610930 128860 611120
rect 128930 610930 128970 611120
rect 129040 610930 129080 611120
rect 129160 610930 129200 611120
rect 129270 610930 129310 611120
rect 129380 610930 129420 611120
rect 129500 610930 129540 611120
rect 129610 610930 129650 611120
rect 129720 610930 129760 611120
rect 129840 610930 129880 611120
rect 129950 610930 129990 611120
rect 130060 610930 130100 611120
rect 130180 610930 130220 611120
rect 130290 610930 130330 611120
rect 130400 610930 130440 611120
rect 130520 610930 130560 611120
rect 130630 610930 130670 611120
rect 130740 610930 130780 611120
rect 130860 610930 130900 611120
rect 130970 610930 131010 611120
rect 131080 610930 131120 611120
rect 131200 610930 131240 611120
rect 131310 610930 131350 611120
rect 131420 610930 131460 611120
rect 131590 610970 131720 611210
rect 131590 610840 131720 610970
rect 131590 610790 131720 610840
rect 125140 605810 125180 605850
rect 125250 605810 125290 605850
rect 125360 605810 125400 605850
rect 131720 605290 131850 605310
rect 125370 605230 125410 605270
rect 125710 605230 125750 605270
rect 126050 605230 126090 605270
rect 126390 605230 126430 605270
rect 126730 605230 126770 605270
rect 127070 605230 127110 605270
rect 127410 605230 127450 605270
rect 127750 605230 127790 605270
rect 128090 605230 128130 605270
rect 128430 605230 128470 605270
rect 128770 605230 128810 605270
rect 129110 605230 129150 605270
rect 129450 605230 129490 605270
rect 129790 605230 129830 605270
rect 130130 605230 130170 605270
rect 130470 605230 130510 605270
rect 130810 605230 130850 605270
rect 131150 605230 131190 605270
rect 131490 605230 131530 605270
rect 131720 605160 131850 605290
rect 125210 604780 125250 605070
rect 125320 604780 125360 605070
rect 125430 604780 125470 605070
rect 125550 604780 125590 605070
rect 125660 604780 125700 605070
rect 125770 604780 125810 605070
rect 125890 604780 125930 605070
rect 126000 604780 126040 605070
rect 126110 604780 126150 605070
rect 126230 604780 126270 605070
rect 126340 604780 126380 605070
rect 126450 604780 126490 605070
rect 126570 604780 126610 605070
rect 126680 604780 126720 605070
rect 126790 604780 126830 605070
rect 126910 604780 126950 605070
rect 127020 604780 127060 605070
rect 127130 604780 127170 605070
rect 127250 604780 127290 605070
rect 127360 604780 127400 605070
rect 127470 604780 127510 605070
rect 127590 604780 127630 605070
rect 127700 604780 127740 605070
rect 127810 604780 127850 605070
rect 127930 604780 127970 605070
rect 128040 604780 128080 605070
rect 128150 604780 128190 605070
rect 128270 604780 128310 605070
rect 128380 604780 128420 605070
rect 128490 604780 128530 605070
rect 128610 604780 128650 605070
rect 128720 604780 128760 605070
rect 128830 604780 128870 605070
rect 128950 604780 128990 605070
rect 129060 604780 129100 605070
rect 129170 604780 129210 605070
rect 129290 604780 129330 605070
rect 129400 604780 129440 605070
rect 129510 604780 129550 605070
rect 129630 604780 129670 605070
rect 129740 604780 129780 605070
rect 129850 604780 129890 605070
rect 129970 604780 130010 605070
rect 130080 604780 130120 605070
rect 130190 604780 130230 605070
rect 130310 604780 130350 605070
rect 130420 604780 130460 605070
rect 130530 604780 130570 605070
rect 130650 604780 130690 605070
rect 130760 604780 130800 605070
rect 130870 604780 130910 605070
rect 130990 604780 131030 605070
rect 131100 604780 131140 605070
rect 131210 604780 131250 605070
rect 131330 604780 131370 605070
rect 131440 604780 131480 605070
rect 131550 604780 131590 605070
rect 131720 604820 131850 605160
rect 131720 604690 131850 604820
rect 131720 604640 131850 604690
rect 124940 599550 124980 599590
rect 125050 599550 125090 599590
rect 125160 599550 125200 599590
rect 131520 599030 131650 599050
rect 125170 598970 125210 599010
rect 125510 598970 125550 599010
rect 125850 598970 125890 599010
rect 126190 598970 126230 599010
rect 126530 598970 126570 599010
rect 126870 598970 126910 599010
rect 127210 598970 127250 599010
rect 127550 598970 127590 599010
rect 127890 598970 127930 599010
rect 128230 598970 128270 599010
rect 128570 598970 128610 599010
rect 128910 598970 128950 599010
rect 129250 598970 129290 599010
rect 129590 598970 129630 599010
rect 129930 598970 129970 599010
rect 130270 598970 130310 599010
rect 130610 598970 130650 599010
rect 130950 598970 130990 599010
rect 131290 598970 131330 599010
rect 131520 598900 131650 599030
rect 125010 598420 125050 598810
rect 125120 598420 125160 598810
rect 125230 598420 125270 598810
rect 125350 598420 125390 598810
rect 125460 598420 125500 598810
rect 125570 598420 125610 598810
rect 125690 598420 125730 598810
rect 125800 598420 125840 598810
rect 125910 598420 125950 598810
rect 126030 598420 126070 598810
rect 126140 598420 126180 598810
rect 126250 598420 126290 598810
rect 126370 598420 126410 598810
rect 126480 598420 126520 598810
rect 126590 598420 126630 598810
rect 126710 598420 126750 598810
rect 126820 598420 126860 598810
rect 126930 598420 126970 598810
rect 127050 598420 127090 598810
rect 127160 598420 127200 598810
rect 127270 598420 127310 598810
rect 127390 598420 127430 598810
rect 127500 598420 127540 598810
rect 127610 598420 127650 598810
rect 127730 598420 127770 598810
rect 127840 598420 127880 598810
rect 127950 598420 127990 598810
rect 128070 598420 128110 598810
rect 128180 598420 128220 598810
rect 128290 598420 128330 598810
rect 128410 598420 128450 598810
rect 128520 598420 128560 598810
rect 128630 598420 128670 598810
rect 128750 598420 128790 598810
rect 128860 598420 128900 598810
rect 128970 598420 129010 598810
rect 129090 598420 129130 598810
rect 129200 598420 129240 598810
rect 129310 598420 129350 598810
rect 129430 598420 129470 598810
rect 129540 598420 129580 598810
rect 129650 598420 129690 598810
rect 129770 598420 129810 598810
rect 129880 598420 129920 598810
rect 129990 598420 130030 598810
rect 130110 598420 130150 598810
rect 130220 598420 130260 598810
rect 130330 598420 130370 598810
rect 130450 598420 130490 598810
rect 130560 598420 130600 598810
rect 130670 598420 130710 598810
rect 130790 598420 130830 598810
rect 130900 598420 130940 598810
rect 131010 598420 131050 598810
rect 131130 598420 131170 598810
rect 131240 598420 131280 598810
rect 131350 598420 131390 598810
rect 131520 598460 131650 598900
rect 131520 598330 131650 598460
rect 131520 598280 131650 598330
rect 119430 593480 119490 593540
rect 119110 593420 119170 593430
rect 119110 593380 119120 593420
rect 119120 593380 119160 593420
rect 119160 593380 119170 593420
rect 119110 593370 119170 593380
rect 119270 592900 119310 592950
rect 119620 592810 119680 592870
rect 119860 593030 119920 593040
rect 119860 592990 119870 593030
rect 119870 592990 119910 593030
rect 119910 592990 119920 593030
rect 119860 592980 119920 592990
rect 119860 592810 119920 592870
rect 120230 593020 120290 593030
rect 120230 592980 120240 593020
rect 120240 592980 120280 593020
rect 120280 592980 120290 593020
rect 120230 592970 120290 592980
rect 119270 592460 119330 592520
rect 124900 592000 124940 592040
rect 125010 592000 125050 592040
rect 125120 592000 125160 592040
rect 131480 591480 131610 591500
rect 125130 591420 125170 591460
rect 125470 591420 125510 591460
rect 125810 591420 125850 591460
rect 126150 591420 126190 591460
rect 126490 591420 126530 591460
rect 126830 591420 126870 591460
rect 127170 591420 127210 591460
rect 127510 591420 127550 591460
rect 127850 591420 127890 591460
rect 128190 591420 128230 591460
rect 128530 591420 128570 591460
rect 128870 591420 128910 591460
rect 129210 591420 129250 591460
rect 129550 591420 129590 591460
rect 129890 591420 129930 591460
rect 130230 591420 130270 591460
rect 130570 591420 130610 591460
rect 130910 591420 130950 591460
rect 131250 591420 131290 591460
rect 131480 591350 131610 591480
rect 124970 590770 125010 591260
rect 125080 590770 125120 591260
rect 125190 590770 125230 591260
rect 125310 590770 125350 591260
rect 125420 590770 125460 591260
rect 125530 590770 125570 591260
rect 125650 590770 125690 591260
rect 125760 590770 125800 591260
rect 125870 590770 125910 591260
rect 125990 590770 126030 591260
rect 126100 590770 126140 591260
rect 126210 590770 126250 591260
rect 126330 590770 126370 591260
rect 126440 590770 126480 591260
rect 126550 590770 126590 591260
rect 126670 590770 126710 591260
rect 126780 590770 126820 591260
rect 126890 590770 126930 591260
rect 127010 590770 127050 591260
rect 127120 590770 127160 591260
rect 127230 590770 127270 591260
rect 127350 590770 127390 591260
rect 127460 590770 127500 591260
rect 127570 590770 127610 591260
rect 127690 590770 127730 591260
rect 127800 590770 127840 591260
rect 127910 590770 127950 591260
rect 128030 590770 128070 591260
rect 128140 590770 128180 591260
rect 128250 590770 128290 591260
rect 128370 590770 128410 591260
rect 128480 590770 128520 591260
rect 128590 590770 128630 591260
rect 128710 590770 128750 591260
rect 128820 590770 128860 591260
rect 128930 590770 128970 591260
rect 129050 590770 129090 591260
rect 129160 590770 129200 591260
rect 129270 590770 129310 591260
rect 129390 590770 129430 591260
rect 129500 590770 129540 591260
rect 129610 590770 129650 591260
rect 129730 590770 129770 591260
rect 129840 590770 129880 591260
rect 129950 590770 129990 591260
rect 130070 590770 130110 591260
rect 130180 590770 130220 591260
rect 130290 590770 130330 591260
rect 130410 590770 130450 591260
rect 130520 590770 130560 591260
rect 130630 590770 130670 591260
rect 130750 590770 130790 591260
rect 130860 590770 130900 591260
rect 130970 590770 131010 591260
rect 131090 590770 131130 591260
rect 131200 590770 131240 591260
rect 131310 590770 131350 591260
rect 131480 590810 131610 591350
rect 131480 590680 131610 590810
rect 131480 590630 131610 590680
rect 119470 583940 119530 584000
rect 119150 583880 119210 583890
rect 119150 583840 119160 583880
rect 119160 583840 119200 583880
rect 119200 583840 119210 583880
rect 119150 583830 119210 583840
rect 119310 583360 119350 583410
rect 119660 583270 119720 583330
rect 119900 583490 119960 583500
rect 119900 583450 119910 583490
rect 119910 583450 119950 583490
rect 119950 583450 119960 583490
rect 119900 583440 119960 583450
rect 119900 583270 119960 583330
rect 120270 583480 120330 583490
rect 120270 583440 120280 583480
rect 120280 583440 120320 583480
rect 120320 583440 120330 583480
rect 120270 583430 120330 583440
rect 125360 583020 125400 583060
rect 125470 583020 125510 583060
rect 125580 583020 125620 583060
rect 119310 582920 119370 582980
rect 132890 582500 133020 582520
rect 125640 582440 125680 582480
rect 126030 582440 126070 582480
rect 126420 582440 126460 582480
rect 126810 582440 126850 582480
rect 127200 582440 127240 582480
rect 127590 582440 127630 582480
rect 127980 582440 128020 582480
rect 128370 582440 128410 582480
rect 128760 582440 128800 582480
rect 129150 582440 129190 582480
rect 129540 582440 129580 582480
rect 129930 582440 129970 582480
rect 130320 582440 130360 582480
rect 130710 582440 130750 582480
rect 131100 582440 131140 582480
rect 131490 582440 131530 582480
rect 131880 582440 131920 582480
rect 132270 582440 132310 582480
rect 132660 582440 132700 582480
rect 132890 582370 133020 582500
rect 125430 582240 125470 582280
rect 125540 582240 125630 582280
rect 125700 582240 125740 582280
rect 125820 582240 125860 582280
rect 125930 582240 126020 582280
rect 126090 582240 126130 582280
rect 126210 582240 126250 582280
rect 126320 582240 126410 582280
rect 126480 582240 126520 582280
rect 126600 582240 126640 582280
rect 126710 582240 126800 582280
rect 126870 582240 126910 582280
rect 126990 582240 127030 582280
rect 127100 582240 127190 582280
rect 127260 582240 127300 582280
rect 127380 582240 127420 582280
rect 127490 582240 127580 582280
rect 127650 582240 127690 582280
rect 127770 582240 127810 582280
rect 127880 582240 127970 582280
rect 128040 582240 128080 582280
rect 128160 582240 128200 582280
rect 128270 582240 128360 582280
rect 128430 582240 128470 582280
rect 128550 582240 128590 582280
rect 128660 582240 128750 582280
rect 128820 582240 128860 582280
rect 128940 582240 128980 582280
rect 129050 582240 129140 582280
rect 129210 582240 129250 582280
rect 129330 582240 129370 582280
rect 129440 582240 129530 582280
rect 129600 582240 129640 582280
rect 129720 582240 129760 582280
rect 129830 582240 129920 582280
rect 129990 582240 130030 582280
rect 130110 582240 130150 582280
rect 130220 582240 130310 582280
rect 130380 582240 130420 582280
rect 130500 582240 130540 582280
rect 130610 582240 130700 582280
rect 130770 582240 130810 582280
rect 130890 582240 130930 582280
rect 131000 582240 131090 582280
rect 131160 582240 131200 582280
rect 131280 582240 131320 582280
rect 131390 582240 131480 582280
rect 131550 582240 131590 582280
rect 131670 582240 131710 582280
rect 131780 582240 131870 582280
rect 131940 582240 131980 582280
rect 132060 582240 132100 582280
rect 132170 582240 132260 582280
rect 132330 582240 132370 582280
rect 132450 582240 132490 582280
rect 132560 582240 132650 582280
rect 132720 582240 132760 582280
rect 132890 582130 133020 582370
rect 132890 582000 133020 582130
rect 132890 581950 133020 582000
rect 119510 574920 119570 574980
rect 119190 574860 119250 574870
rect 119190 574820 119200 574860
rect 119200 574820 119240 574860
rect 119240 574820 119250 574860
rect 119190 574810 119250 574820
rect 119350 574340 119390 574390
rect 119700 574250 119760 574310
rect 119940 574470 120000 574480
rect 119940 574430 119950 574470
rect 119950 574430 119990 574470
rect 119990 574430 120000 574470
rect 119940 574420 120000 574430
rect 119940 574250 120000 574310
rect 120310 574460 120370 574470
rect 120310 574420 120320 574460
rect 120320 574420 120360 574460
rect 120360 574420 120370 574460
rect 120310 574410 120370 574420
rect 125400 574000 125440 574040
rect 125510 574000 125550 574040
rect 125620 574000 125660 574040
rect 119350 573900 119410 573960
rect 132930 573480 133060 573500
rect 125680 573420 125720 573460
rect 126070 573420 126110 573460
rect 126460 573420 126500 573460
rect 126850 573420 126890 573460
rect 127240 573420 127280 573460
rect 127630 573420 127670 573460
rect 128020 573420 128060 573460
rect 128410 573420 128450 573460
rect 128800 573420 128840 573460
rect 129190 573420 129230 573460
rect 129580 573420 129620 573460
rect 129970 573420 130010 573460
rect 130360 573420 130400 573460
rect 130750 573420 130790 573460
rect 131140 573420 131180 573460
rect 131530 573420 131570 573460
rect 131920 573420 131960 573460
rect 132310 573420 132350 573460
rect 132700 573420 132740 573460
rect 132930 573350 133060 573480
rect 125470 573120 125510 573260
rect 125580 573120 125670 573260
rect 125740 573120 125780 573260
rect 125860 573120 125900 573260
rect 125970 573120 126060 573260
rect 126130 573120 126170 573260
rect 126250 573120 126290 573260
rect 126360 573120 126450 573260
rect 126520 573120 126560 573260
rect 126640 573120 126680 573260
rect 126750 573120 126840 573260
rect 126910 573120 126950 573260
rect 127030 573120 127070 573260
rect 127140 573120 127230 573260
rect 127300 573120 127340 573260
rect 127420 573120 127460 573260
rect 127530 573120 127620 573260
rect 127690 573120 127730 573260
rect 127810 573120 127850 573260
rect 127920 573120 128010 573260
rect 128080 573120 128120 573260
rect 128200 573120 128240 573260
rect 128310 573120 128400 573260
rect 128470 573120 128510 573260
rect 128590 573120 128630 573260
rect 128700 573120 128790 573260
rect 128860 573120 128900 573260
rect 128980 573120 129020 573260
rect 129090 573120 129180 573260
rect 129250 573120 129290 573260
rect 129370 573120 129410 573260
rect 129480 573120 129570 573260
rect 129640 573120 129680 573260
rect 129760 573120 129800 573260
rect 129870 573120 129960 573260
rect 130030 573120 130070 573260
rect 130150 573120 130190 573260
rect 130260 573120 130350 573260
rect 130420 573120 130460 573260
rect 130540 573120 130580 573260
rect 130650 573120 130740 573260
rect 130810 573120 130850 573260
rect 130930 573120 130970 573260
rect 131040 573120 131130 573260
rect 131200 573120 131240 573260
rect 131320 573120 131360 573260
rect 131430 573120 131520 573260
rect 131590 573120 131630 573260
rect 131710 573120 131750 573260
rect 131820 573120 131910 573260
rect 131980 573120 132020 573260
rect 132100 573120 132140 573260
rect 132210 573120 132300 573260
rect 132370 573120 132410 573260
rect 132490 573120 132530 573260
rect 132600 573120 132690 573260
rect 132760 573120 132800 573260
rect 132930 573010 133060 573350
rect 132930 572880 133060 573010
rect 132930 572830 133060 572880
rect 119460 567250 119520 567310
rect 119140 567190 119200 567200
rect 119140 567150 119150 567190
rect 119150 567150 119190 567190
rect 119190 567150 119200 567190
rect 119140 567140 119200 567150
rect 119300 566670 119340 566720
rect 119650 566580 119710 566640
rect 119890 566800 119950 566810
rect 119890 566760 119900 566800
rect 119900 566760 119940 566800
rect 119940 566760 119950 566800
rect 119890 566750 119950 566760
rect 119890 566580 119950 566640
rect 120260 566790 120320 566800
rect 120260 566750 120270 566790
rect 120270 566750 120310 566790
rect 120310 566750 120320 566790
rect 120260 566740 120320 566750
rect 125350 566330 125390 566370
rect 125460 566330 125500 566370
rect 125570 566330 125610 566370
rect 119300 566230 119360 566290
rect 132880 565810 133010 565830
rect 125630 565750 125670 565790
rect 126020 565750 126060 565790
rect 126410 565750 126450 565790
rect 126800 565750 126840 565790
rect 127190 565750 127230 565790
rect 127580 565750 127620 565790
rect 127970 565750 128010 565790
rect 128360 565750 128400 565790
rect 128750 565750 128790 565790
rect 129140 565750 129180 565790
rect 129530 565750 129570 565790
rect 129920 565750 129960 565790
rect 130310 565750 130350 565790
rect 130700 565750 130740 565790
rect 131090 565750 131130 565790
rect 131480 565750 131520 565790
rect 131870 565750 131910 565790
rect 132260 565750 132300 565790
rect 132650 565750 132690 565790
rect 132880 565680 133010 565810
rect 125420 565350 125460 565590
rect 125530 565350 125620 565590
rect 125690 565350 125730 565590
rect 125810 565350 125850 565590
rect 125920 565350 126010 565590
rect 126080 565350 126120 565590
rect 126200 565350 126240 565590
rect 126310 565350 126400 565590
rect 126470 565350 126510 565590
rect 126590 565350 126630 565590
rect 126700 565350 126790 565590
rect 126860 565350 126900 565590
rect 126980 565350 127020 565590
rect 127090 565350 127180 565590
rect 127250 565350 127290 565590
rect 127370 565350 127410 565590
rect 127480 565350 127570 565590
rect 127640 565350 127680 565590
rect 127760 565350 127800 565590
rect 127870 565350 127960 565590
rect 128030 565350 128070 565590
rect 128150 565350 128190 565590
rect 128260 565350 128350 565590
rect 128420 565350 128460 565590
rect 128540 565350 128580 565590
rect 128650 565350 128740 565590
rect 128810 565350 128850 565590
rect 128930 565350 128970 565590
rect 129040 565350 129130 565590
rect 129200 565350 129240 565590
rect 129320 565350 129360 565590
rect 129430 565350 129520 565590
rect 129590 565350 129630 565590
rect 129710 565350 129750 565590
rect 129820 565350 129910 565590
rect 129980 565350 130020 565590
rect 130100 565350 130140 565590
rect 130210 565350 130300 565590
rect 130370 565350 130410 565590
rect 130490 565350 130530 565590
rect 130600 565350 130690 565590
rect 130760 565350 130800 565590
rect 130880 565350 130920 565590
rect 130990 565350 131080 565590
rect 131150 565350 131190 565590
rect 131270 565350 131310 565590
rect 131380 565350 131470 565590
rect 131540 565350 131580 565590
rect 131660 565350 131700 565590
rect 131770 565350 131860 565590
rect 131930 565350 131970 565590
rect 132050 565350 132090 565590
rect 132160 565350 132250 565590
rect 132320 565350 132360 565590
rect 132440 565350 132480 565590
rect 132550 565350 132640 565590
rect 132710 565350 132750 565590
rect 132880 565240 133010 565680
rect 132880 565110 133010 565240
rect 132880 565060 133010 565110
rect 119460 560710 119520 560770
rect 119140 560650 119200 560660
rect 119140 560610 119150 560650
rect 119150 560610 119190 560650
rect 119190 560610 119200 560650
rect 119140 560600 119200 560610
rect 119300 560130 119340 560180
rect 119650 560040 119710 560100
rect 119890 560260 119950 560270
rect 119890 560220 119900 560260
rect 119900 560220 119940 560260
rect 119940 560220 119950 560260
rect 119890 560210 119950 560220
rect 119890 560040 119950 560100
rect 120260 560250 120320 560260
rect 120260 560210 120270 560250
rect 120270 560210 120310 560250
rect 120310 560210 120320 560250
rect 120260 560200 120320 560210
rect 125350 559790 125390 559830
rect 125460 559790 125500 559830
rect 125570 559790 125610 559830
rect 119300 559690 119360 559750
rect 132880 559270 133010 559290
rect 125630 559210 125670 559250
rect 126020 559210 126060 559250
rect 126410 559210 126450 559250
rect 126800 559210 126840 559250
rect 127190 559210 127230 559250
rect 127580 559210 127620 559250
rect 127970 559210 128010 559250
rect 128360 559210 128400 559250
rect 128750 559210 128790 559250
rect 129140 559210 129180 559250
rect 129530 559210 129570 559250
rect 129920 559210 129960 559250
rect 130310 559210 130350 559250
rect 130700 559210 130740 559250
rect 131090 559210 131130 559250
rect 131480 559210 131520 559250
rect 131870 559210 131910 559250
rect 132260 559210 132300 559250
rect 132650 559210 132690 559250
rect 132880 559140 133010 559270
rect 125420 558710 125460 559050
rect 125530 558710 125620 559050
rect 125690 558710 125730 559050
rect 125810 558710 125850 559050
rect 125920 558710 126010 559050
rect 126080 558710 126120 559050
rect 126200 558710 126240 559050
rect 126310 558710 126400 559050
rect 126470 558710 126510 559050
rect 126590 558710 126630 559050
rect 126700 558710 126790 559050
rect 126860 558710 126900 559050
rect 126980 558710 127020 559050
rect 127090 558710 127180 559050
rect 127250 558710 127290 559050
rect 127370 558710 127410 559050
rect 127480 558710 127570 559050
rect 127640 558710 127680 559050
rect 127760 558710 127800 559050
rect 127870 558710 127960 559050
rect 128030 558710 128070 559050
rect 128150 558710 128190 559050
rect 128260 558710 128350 559050
rect 128420 558710 128460 559050
rect 128540 558710 128580 559050
rect 128650 558710 128740 559050
rect 128810 558710 128850 559050
rect 128930 558710 128970 559050
rect 129040 558710 129130 559050
rect 129200 558710 129240 559050
rect 129320 558710 129360 559050
rect 129430 558710 129520 559050
rect 129590 558710 129630 559050
rect 129710 558710 129750 559050
rect 129820 558710 129910 559050
rect 129980 558710 130020 559050
rect 130100 558710 130140 559050
rect 130210 558710 130300 559050
rect 130370 558710 130410 559050
rect 130490 558710 130530 559050
rect 130600 558710 130690 559050
rect 130760 558710 130800 559050
rect 130880 558710 130920 559050
rect 130990 558710 131080 559050
rect 131150 558710 131190 559050
rect 131270 558710 131310 559050
rect 131380 558710 131470 559050
rect 131540 558710 131580 559050
rect 131660 558710 131700 559050
rect 131770 558710 131860 559050
rect 131930 558710 131970 559050
rect 132050 558710 132090 559050
rect 132160 558710 132250 559050
rect 132320 558710 132360 559050
rect 132440 558710 132480 559050
rect 132550 558710 132640 559050
rect 132710 558710 132750 559050
rect 132880 558600 133010 559140
rect 132880 558470 133010 558600
rect 132880 558420 133010 558470
rect 119530 553880 119590 553940
rect 125000 553930 125040 553970
rect 125110 553930 125150 553970
rect 125220 553930 125260 553970
rect 119210 553820 119270 553830
rect 119210 553780 119220 553820
rect 119220 553780 119260 553820
rect 119260 553780 119270 553820
rect 119210 553770 119270 553780
rect 119370 553300 119410 553350
rect 119720 553210 119780 553270
rect 119960 553430 120020 553440
rect 119960 553390 119970 553430
rect 119970 553390 120010 553430
rect 120010 553390 120020 553430
rect 119960 553380 120020 553390
rect 119960 553210 120020 553270
rect 120330 553420 120390 553430
rect 120330 553380 120340 553420
rect 120340 553380 120380 553420
rect 120380 553380 120390 553420
rect 120330 553370 120390 553380
rect 119370 552860 119430 552920
rect 133900 552440 134030 552460
rect 125750 552380 125790 552420
rect 126190 552380 126230 552420
rect 126630 552380 126670 552420
rect 127070 552380 127110 552420
rect 127510 552380 127550 552420
rect 127950 552380 127990 552420
rect 128390 552380 128430 552420
rect 128830 552380 128870 552420
rect 129270 552380 129310 552420
rect 129710 552380 129750 552420
rect 130150 552380 130190 552420
rect 130590 552380 130630 552420
rect 131030 552380 131070 552420
rect 131470 552380 131510 552420
rect 131910 552380 131950 552420
rect 132350 552380 132390 552420
rect 132790 552380 132830 552420
rect 133230 552380 133270 552420
rect 133670 552380 133710 552420
rect 133900 552310 134030 552440
rect 125490 552180 125530 552220
rect 125600 552180 125740 552220
rect 125810 552180 125850 552220
rect 125930 552180 125970 552220
rect 126040 552180 126180 552220
rect 126250 552180 126290 552220
rect 126370 552180 126410 552220
rect 126480 552180 126620 552220
rect 126690 552180 126730 552220
rect 126810 552180 126850 552220
rect 126920 552180 127060 552220
rect 127130 552180 127170 552220
rect 127250 552180 127290 552220
rect 127360 552180 127500 552220
rect 127570 552180 127610 552220
rect 127690 552180 127730 552220
rect 127800 552180 127940 552220
rect 128010 552180 128050 552220
rect 128130 552180 128170 552220
rect 128240 552180 128380 552220
rect 128450 552180 128490 552220
rect 128570 552180 128610 552220
rect 128680 552180 128820 552220
rect 128890 552180 128930 552220
rect 129010 552180 129050 552220
rect 129120 552180 129260 552220
rect 129330 552180 129370 552220
rect 129450 552180 129490 552220
rect 129560 552180 129700 552220
rect 129770 552180 129810 552220
rect 129890 552180 129930 552220
rect 130000 552180 130140 552220
rect 130210 552180 130250 552220
rect 130330 552180 130370 552220
rect 130440 552180 130580 552220
rect 130650 552180 130690 552220
rect 130770 552180 130810 552220
rect 130880 552180 131020 552220
rect 131090 552180 131130 552220
rect 131210 552180 131250 552220
rect 131320 552180 131460 552220
rect 131530 552180 131570 552220
rect 131650 552180 131690 552220
rect 131760 552180 131900 552220
rect 131970 552180 132010 552220
rect 132090 552180 132130 552220
rect 132200 552180 132340 552220
rect 132410 552180 132450 552220
rect 132530 552180 132570 552220
rect 132640 552180 132780 552220
rect 132850 552180 132890 552220
rect 132970 552180 133010 552220
rect 133080 552180 133220 552220
rect 133290 552180 133330 552220
rect 133410 552180 133450 552220
rect 133520 552180 133660 552220
rect 133730 552180 133770 552220
rect 133900 552070 134030 552310
rect 133900 551940 134030 552070
rect 133900 551890 134030 551940
rect 119530 546310 119590 546370
rect 125000 546360 125040 546400
rect 125110 546360 125150 546400
rect 125220 546360 125260 546400
rect 119210 546250 119270 546260
rect 119210 546210 119220 546250
rect 119220 546210 119260 546250
rect 119260 546210 119270 546250
rect 119210 546200 119270 546210
rect 119370 545730 119410 545780
rect 119720 545640 119780 545700
rect 119960 545860 120020 545870
rect 119960 545820 119970 545860
rect 119970 545820 120010 545860
rect 120010 545820 120020 545860
rect 119960 545810 120020 545820
rect 119960 545640 120020 545700
rect 120330 545850 120390 545860
rect 120330 545810 120340 545850
rect 120340 545810 120380 545850
rect 120380 545810 120390 545850
rect 120330 545800 120390 545810
rect 119370 545290 119430 545350
rect 133900 544870 134030 544890
rect 125750 544810 125790 544850
rect 126190 544810 126230 544850
rect 126630 544810 126670 544850
rect 127070 544810 127110 544850
rect 127510 544810 127550 544850
rect 127950 544810 127990 544850
rect 128390 544810 128430 544850
rect 128830 544810 128870 544850
rect 129270 544810 129310 544850
rect 129710 544810 129750 544850
rect 130150 544810 130190 544850
rect 130590 544810 130630 544850
rect 131030 544810 131070 544850
rect 131470 544810 131510 544850
rect 131910 544810 131950 544850
rect 132350 544810 132390 544850
rect 132790 544810 132830 544850
rect 133230 544810 133270 544850
rect 133670 544810 133710 544850
rect 133900 544740 134030 544870
rect 125490 544410 125530 544650
rect 125600 544410 125740 544650
rect 125810 544410 125850 544650
rect 125930 544410 125970 544650
rect 126040 544410 126180 544650
rect 126250 544410 126290 544650
rect 126370 544410 126410 544650
rect 126480 544410 126620 544650
rect 126690 544410 126730 544650
rect 126810 544410 126850 544650
rect 126920 544410 127060 544650
rect 127130 544410 127170 544650
rect 127250 544410 127290 544650
rect 127360 544410 127500 544650
rect 127570 544410 127610 544650
rect 127690 544410 127730 544650
rect 127800 544410 127940 544650
rect 128010 544410 128050 544650
rect 128130 544410 128170 544650
rect 128240 544410 128380 544650
rect 128450 544410 128490 544650
rect 128570 544410 128610 544650
rect 128680 544410 128820 544650
rect 128890 544410 128930 544650
rect 129010 544410 129050 544650
rect 129120 544410 129260 544650
rect 129330 544410 129370 544650
rect 129450 544410 129490 544650
rect 129560 544410 129700 544650
rect 129770 544410 129810 544650
rect 129890 544410 129930 544650
rect 130000 544410 130140 544650
rect 130210 544410 130250 544650
rect 130330 544410 130370 544650
rect 130440 544410 130580 544650
rect 130650 544410 130690 544650
rect 130770 544410 130810 544650
rect 130880 544410 131020 544650
rect 131090 544410 131130 544650
rect 131210 544410 131250 544650
rect 131320 544410 131460 544650
rect 131530 544410 131570 544650
rect 131650 544410 131690 544650
rect 131760 544410 131900 544650
rect 131970 544410 132010 544650
rect 132090 544410 132130 544650
rect 132200 544410 132340 544650
rect 132410 544410 132450 544650
rect 132530 544410 132570 544650
rect 132640 544410 132780 544650
rect 132850 544410 132890 544650
rect 132970 544410 133010 544650
rect 133080 544410 133220 544650
rect 133290 544410 133330 544650
rect 133410 544410 133450 544650
rect 133520 544410 133660 544650
rect 133730 544410 133770 544650
rect 133900 544300 134030 544740
rect 133900 544170 134030 544300
rect 133900 544120 134030 544170
rect 119500 538250 119560 538310
rect 124970 538300 125010 538340
rect 125080 538300 125120 538340
rect 125190 538300 125230 538340
rect 119180 538190 119240 538200
rect 119180 538150 119190 538190
rect 119190 538150 119230 538190
rect 119230 538150 119240 538190
rect 119180 538140 119240 538150
rect 119340 537670 119380 537720
rect 119690 537580 119750 537640
rect 119930 537800 119990 537810
rect 119930 537760 119940 537800
rect 119940 537760 119980 537800
rect 119980 537760 119990 537800
rect 119930 537750 119990 537760
rect 119930 537580 119990 537640
rect 120300 537790 120360 537800
rect 120300 537750 120310 537790
rect 120310 537750 120350 537790
rect 120350 537750 120360 537790
rect 120300 537740 120360 537750
rect 119340 537230 119400 537290
rect 133870 536810 134000 536830
rect 125720 536750 125760 536790
rect 126160 536750 126200 536790
rect 126600 536750 126640 536790
rect 127040 536750 127080 536790
rect 127480 536750 127520 536790
rect 127920 536750 127960 536790
rect 128360 536750 128400 536790
rect 128800 536750 128840 536790
rect 129240 536750 129280 536790
rect 129680 536750 129720 536790
rect 130120 536750 130160 536790
rect 130560 536750 130600 536790
rect 131000 536750 131040 536790
rect 131440 536750 131480 536790
rect 131880 536750 131920 536790
rect 132320 536750 132360 536790
rect 132760 536750 132800 536790
rect 133200 536750 133240 536790
rect 133640 536750 133680 536790
rect 133870 536680 134000 536810
rect 125460 536150 125500 536590
rect 125570 536150 125710 536590
rect 125780 536150 125820 536590
rect 125900 536150 125940 536590
rect 126010 536150 126150 536590
rect 126220 536150 126260 536590
rect 126340 536150 126380 536590
rect 126450 536150 126590 536590
rect 126660 536150 126700 536590
rect 126780 536150 126820 536590
rect 126890 536150 127030 536590
rect 127100 536150 127140 536590
rect 127220 536150 127260 536590
rect 127330 536150 127470 536590
rect 127540 536150 127580 536590
rect 127660 536150 127700 536590
rect 127770 536150 127910 536590
rect 127980 536150 128020 536590
rect 128100 536150 128140 536590
rect 128210 536150 128350 536590
rect 128420 536150 128460 536590
rect 128540 536150 128580 536590
rect 128650 536150 128790 536590
rect 128860 536150 128900 536590
rect 128980 536150 129020 536590
rect 129090 536150 129230 536590
rect 129300 536150 129340 536590
rect 129420 536150 129460 536590
rect 129530 536150 129670 536590
rect 129740 536150 129780 536590
rect 129860 536150 129900 536590
rect 129970 536150 130110 536590
rect 130180 536150 130220 536590
rect 130300 536150 130340 536590
rect 130410 536150 130550 536590
rect 130620 536150 130660 536590
rect 130740 536150 130780 536590
rect 130850 536150 130990 536590
rect 131060 536150 131100 536590
rect 131180 536150 131220 536590
rect 131290 536150 131430 536590
rect 131500 536150 131540 536590
rect 131620 536150 131660 536590
rect 131730 536150 131870 536590
rect 131940 536150 131980 536590
rect 132060 536150 132100 536590
rect 132170 536150 132310 536590
rect 132380 536150 132420 536590
rect 132500 536150 132540 536590
rect 132610 536150 132750 536590
rect 132820 536150 132860 536590
rect 132940 536150 132980 536590
rect 133050 536150 133190 536590
rect 133260 536150 133300 536590
rect 133380 536150 133420 536590
rect 133490 536150 133630 536590
rect 133700 536150 133740 536590
rect 133870 536040 134000 536680
rect 133870 535910 134000 536040
rect 133870 535860 134000 535910
<< metal1 >>
rect 82716 687251 85076 687282
rect 82712 687217 85076 687251
rect 82716 687192 85076 687217
rect 82696 686707 85056 686732
rect 82696 686673 85079 686707
rect 82696 686642 85056 686673
rect 102326 651972 102426 651978
rect 102326 651962 102332 651972
rect 102041 651892 102332 651962
rect 102424 651892 102426 651972
rect 102041 651866 102426 651892
rect 102041 651546 102137 651866
rect 102326 651856 102426 651866
rect 102041 651450 102550 651546
rect 102041 650461 102137 651450
rect 115242 650993 115661 651002
rect 115242 650906 115700 650993
rect 102041 650365 102506 650461
rect 102041 649372 102137 650365
rect 115622 649914 115700 650906
rect 115242 649818 115700 649914
rect 102041 649276 102514 649372
rect 102041 648273 102137 649276
rect 115622 648826 115700 649818
rect 115242 648730 115700 648826
rect 102041 648177 102534 648273
rect 102041 647198 102137 648177
rect 115622 647738 115700 648730
rect 115242 647642 115700 647738
rect 102041 647102 102516 647198
rect 95499 646722 96634 646815
rect 95499 644429 95870 646722
rect 96526 645904 96634 646722
rect 102041 646099 102137 647102
rect 115622 646650 115700 647642
rect 115242 646554 115700 646650
rect 102041 646003 102546 646099
rect 102041 645904 102137 646003
rect 96526 645263 102137 645904
rect 115622 645562 115700 646554
rect 119290 646200 119390 646206
rect 119290 646120 119296 646200
rect 119388 646120 119390 646200
rect 119112 646006 119242 646020
rect 119112 645916 119128 646006
rect 119228 645916 119242 646006
rect 119112 645902 119242 645916
rect 119290 645910 119390 646120
rect 119962 646018 120062 646024
rect 119962 646010 119968 646018
rect 119450 645938 119968 646010
rect 120060 645938 120062 646018
rect 119450 645910 120062 645938
rect 119962 645902 120062 645910
rect 115242 645466 115700 645562
rect 96526 644429 96634 645263
rect 95499 644298 96634 644429
rect 102041 645014 102137 645263
rect 102041 644918 102549 645014
rect 102041 643933 102137 644918
rect 115622 644474 115700 645466
rect 115242 644378 115700 644474
rect 102041 643837 102490 643933
rect 102041 642842 102137 643837
rect 115622 643386 115700 644378
rect 115242 643290 115700 643386
rect 102041 642746 102568 642842
rect 102041 641737 102137 642746
rect 115622 642298 115700 643290
rect 120760 642790 120860 645240
rect 120760 642750 124100 642790
rect 120760 642710 124040 642750
rect 124080 642710 124100 642750
rect 120760 642690 124100 642710
rect 127460 642780 128360 642790
rect 127460 642700 127470 642780
rect 128350 642700 128360 642780
rect 115242 642202 115700 642298
rect 102041 641641 102501 641737
rect 102041 640653 102137 641641
rect 115622 641210 115700 642202
rect 123800 642610 123990 642630
rect 127460 642610 128360 642700
rect 131470 642630 131660 642650
rect 123800 642040 123830 642610
rect 123960 642040 123990 642610
rect 124150 642530 131350 642610
rect 124150 642500 124240 642530
rect 124150 642450 124170 642500
rect 124220 642450 124240 642500
rect 124150 642430 124240 642450
rect 124330 642500 124420 642530
rect 124330 642450 124350 642500
rect 124400 642450 124420 642500
rect 124330 642430 124420 642450
rect 124510 642500 124600 642530
rect 124510 642450 124530 642500
rect 124580 642450 124600 642500
rect 124510 642430 124600 642450
rect 124690 642500 124780 642530
rect 124690 642450 124710 642500
rect 124760 642450 124780 642500
rect 124690 642430 124780 642450
rect 124870 642500 124960 642530
rect 124870 642450 124890 642500
rect 124940 642450 124960 642500
rect 124870 642430 124960 642450
rect 125050 642500 125140 642530
rect 125050 642450 125070 642500
rect 125120 642450 125140 642500
rect 125050 642430 125140 642450
rect 125230 642500 125320 642530
rect 125230 642450 125250 642500
rect 125300 642450 125320 642500
rect 125230 642430 125320 642450
rect 125410 642500 125500 642530
rect 125410 642450 125430 642500
rect 125480 642450 125500 642500
rect 125410 642430 125500 642450
rect 125590 642500 125680 642530
rect 125590 642450 125610 642500
rect 125660 642450 125680 642500
rect 125590 642430 125680 642450
rect 125770 642500 125860 642530
rect 125770 642450 125790 642500
rect 125840 642450 125860 642500
rect 125770 642430 125860 642450
rect 125950 642500 126040 642530
rect 125950 642450 125970 642500
rect 126020 642450 126040 642500
rect 125950 642430 126040 642450
rect 126130 642500 126220 642530
rect 126130 642450 126150 642500
rect 126200 642450 126220 642500
rect 126130 642430 126220 642450
rect 126310 642500 126400 642530
rect 126310 642450 126330 642500
rect 126380 642450 126400 642500
rect 126310 642430 126400 642450
rect 126490 642500 126580 642530
rect 126490 642450 126510 642500
rect 126560 642450 126580 642500
rect 126490 642430 126580 642450
rect 126670 642500 126760 642530
rect 126670 642450 126690 642500
rect 126740 642450 126760 642500
rect 126670 642430 126760 642450
rect 126850 642500 126940 642530
rect 126850 642450 126870 642500
rect 126920 642450 126940 642500
rect 126850 642430 126940 642450
rect 127030 642500 127120 642530
rect 127030 642450 127050 642500
rect 127100 642450 127120 642500
rect 127030 642430 127120 642450
rect 127210 642500 127300 642530
rect 127210 642450 127230 642500
rect 127280 642450 127300 642500
rect 127210 642430 127300 642450
rect 127390 642500 127480 642530
rect 127390 642450 127410 642500
rect 127460 642450 127480 642500
rect 127390 642430 127480 642450
rect 127570 642500 127660 642530
rect 127570 642450 127590 642500
rect 127640 642450 127660 642500
rect 127570 642430 127660 642450
rect 127750 642500 127840 642530
rect 127750 642450 127770 642500
rect 127820 642450 127840 642500
rect 127750 642430 127840 642450
rect 127930 642500 128020 642530
rect 127930 642450 127950 642500
rect 128000 642450 128020 642500
rect 127930 642430 128020 642450
rect 128110 642500 128200 642530
rect 128110 642450 128130 642500
rect 128180 642450 128200 642500
rect 128110 642430 128200 642450
rect 128290 642500 128380 642530
rect 128290 642450 128310 642500
rect 128360 642450 128380 642500
rect 128290 642430 128380 642450
rect 128470 642500 128560 642530
rect 128470 642450 128490 642500
rect 128540 642450 128560 642500
rect 128470 642430 128560 642450
rect 128650 642500 128740 642530
rect 128650 642450 128670 642500
rect 128720 642450 128740 642500
rect 128650 642430 128740 642450
rect 128830 642500 128920 642530
rect 128830 642450 128850 642500
rect 128900 642450 128920 642500
rect 128830 642430 128920 642450
rect 129010 642500 129100 642530
rect 129010 642450 129030 642500
rect 129080 642450 129100 642500
rect 129010 642430 129100 642450
rect 129190 642500 129280 642530
rect 129190 642450 129210 642500
rect 129260 642450 129280 642500
rect 129190 642430 129280 642450
rect 129370 642500 129460 642530
rect 129370 642450 129390 642500
rect 129440 642450 129460 642500
rect 129370 642430 129460 642450
rect 129550 642500 129640 642530
rect 129550 642450 129570 642500
rect 129620 642450 129640 642500
rect 129550 642430 129640 642450
rect 129730 642500 129820 642530
rect 129730 642450 129750 642500
rect 129800 642450 129820 642500
rect 129730 642430 129820 642450
rect 129910 642500 130000 642530
rect 129910 642450 129930 642500
rect 129980 642450 130000 642500
rect 129910 642430 130000 642450
rect 130090 642500 130180 642530
rect 130090 642450 130110 642500
rect 130160 642450 130180 642500
rect 130090 642430 130180 642450
rect 130270 642500 130360 642530
rect 130270 642450 130290 642500
rect 130340 642450 130360 642500
rect 130270 642430 130360 642450
rect 130450 642500 130540 642530
rect 130450 642450 130470 642500
rect 130520 642450 130540 642500
rect 130450 642430 130540 642450
rect 130630 642500 130720 642530
rect 130630 642450 130650 642500
rect 130700 642450 130720 642500
rect 130630 642430 130720 642450
rect 130810 642500 130900 642530
rect 130810 642450 130830 642500
rect 130880 642450 130900 642500
rect 130810 642430 130900 642450
rect 130990 642500 131080 642530
rect 130990 642450 131010 642500
rect 131060 642450 131080 642500
rect 130990 642430 131080 642450
rect 131170 642500 131260 642530
rect 131170 642450 131190 642500
rect 131240 642450 131260 642500
rect 131170 642430 131260 642450
rect 124150 642200 124240 642220
rect 124150 642150 124170 642200
rect 124220 642150 124240 642200
rect 124150 642120 124240 642150
rect 124330 642200 124420 642220
rect 124330 642150 124350 642200
rect 124400 642150 124420 642200
rect 124330 642120 124420 642150
rect 124510 642200 124600 642220
rect 124510 642150 124530 642200
rect 124580 642150 124600 642200
rect 124510 642120 124600 642150
rect 124690 642200 124780 642220
rect 124690 642150 124710 642200
rect 124760 642150 124780 642200
rect 124690 642120 124780 642150
rect 124870 642200 124960 642220
rect 124870 642150 124890 642200
rect 124940 642150 124960 642200
rect 124870 642120 124960 642150
rect 125050 642200 125140 642220
rect 125050 642150 125070 642200
rect 125120 642150 125140 642200
rect 125050 642120 125140 642150
rect 125230 642200 125320 642220
rect 125230 642150 125250 642200
rect 125300 642150 125320 642200
rect 125230 642120 125320 642150
rect 125410 642200 125500 642220
rect 125410 642150 125430 642200
rect 125480 642150 125500 642200
rect 125410 642120 125500 642150
rect 125590 642200 125680 642220
rect 125590 642150 125610 642200
rect 125660 642150 125680 642200
rect 125590 642120 125680 642150
rect 125770 642200 125860 642220
rect 125770 642150 125790 642200
rect 125840 642150 125860 642200
rect 125770 642120 125860 642150
rect 125950 642200 126040 642220
rect 125950 642150 125970 642200
rect 126020 642150 126040 642200
rect 125950 642120 126040 642150
rect 126130 642200 126220 642220
rect 126130 642150 126150 642200
rect 126200 642150 126220 642200
rect 126130 642120 126220 642150
rect 126310 642200 126400 642220
rect 126310 642150 126330 642200
rect 126380 642150 126400 642200
rect 126310 642120 126400 642150
rect 126490 642200 126580 642220
rect 126490 642150 126510 642200
rect 126560 642150 126580 642200
rect 126490 642120 126580 642150
rect 126670 642200 126760 642220
rect 126670 642150 126690 642200
rect 126740 642150 126760 642200
rect 126670 642120 126760 642150
rect 126850 642200 126940 642220
rect 126850 642150 126870 642200
rect 126920 642150 126940 642200
rect 126850 642120 126940 642150
rect 127030 642200 127120 642220
rect 127030 642150 127050 642200
rect 127100 642150 127120 642200
rect 127030 642120 127120 642150
rect 127210 642200 127300 642220
rect 127210 642150 127230 642200
rect 127280 642150 127300 642200
rect 127210 642120 127300 642150
rect 127390 642200 127480 642220
rect 127390 642150 127410 642200
rect 127460 642150 127480 642200
rect 127390 642120 127480 642150
rect 127570 642200 127660 642220
rect 127570 642150 127590 642200
rect 127640 642150 127660 642200
rect 127570 642120 127660 642150
rect 127750 642200 127840 642220
rect 127750 642150 127770 642200
rect 127820 642150 127840 642200
rect 127750 642120 127840 642150
rect 127930 642200 128020 642220
rect 127930 642150 127950 642200
rect 128000 642150 128020 642200
rect 127930 642120 128020 642150
rect 128110 642200 128200 642220
rect 128110 642150 128130 642200
rect 128180 642150 128200 642200
rect 128110 642120 128200 642150
rect 128290 642200 128380 642220
rect 128290 642150 128310 642200
rect 128360 642150 128380 642200
rect 128290 642120 128380 642150
rect 128470 642200 128560 642220
rect 128470 642150 128490 642200
rect 128540 642150 128560 642200
rect 128470 642120 128560 642150
rect 128650 642200 128740 642220
rect 128650 642150 128670 642200
rect 128720 642150 128740 642200
rect 128650 642120 128740 642150
rect 128830 642200 128920 642220
rect 128830 642150 128850 642200
rect 128900 642150 128920 642200
rect 128830 642120 128920 642150
rect 129010 642200 129100 642220
rect 129010 642150 129030 642200
rect 129080 642150 129100 642200
rect 129010 642120 129100 642150
rect 129190 642200 129280 642220
rect 129190 642150 129210 642200
rect 129260 642150 129280 642200
rect 129190 642120 129280 642150
rect 129370 642200 129460 642220
rect 129370 642150 129390 642200
rect 129440 642150 129460 642200
rect 129370 642120 129460 642150
rect 129550 642200 129640 642220
rect 129550 642150 129570 642200
rect 129620 642150 129640 642200
rect 129550 642120 129640 642150
rect 129730 642200 129820 642220
rect 129730 642150 129750 642200
rect 129800 642150 129820 642200
rect 129730 642120 129820 642150
rect 129910 642200 130000 642220
rect 129910 642150 129930 642200
rect 129980 642150 130000 642200
rect 129910 642120 130000 642150
rect 130090 642200 130180 642220
rect 130090 642150 130110 642200
rect 130160 642150 130180 642200
rect 130090 642120 130180 642150
rect 130270 642200 130360 642220
rect 130270 642150 130290 642200
rect 130340 642150 130360 642200
rect 130270 642120 130360 642150
rect 130450 642200 130540 642220
rect 130450 642150 130470 642200
rect 130520 642150 130540 642200
rect 130450 642120 130540 642150
rect 130630 642200 130720 642220
rect 130630 642150 130650 642200
rect 130700 642150 130720 642200
rect 130630 642120 130720 642150
rect 130810 642200 130900 642220
rect 130810 642150 130830 642200
rect 130880 642150 130900 642200
rect 130810 642120 130900 642150
rect 130990 642200 131080 642220
rect 130990 642150 131010 642200
rect 131060 642150 131080 642200
rect 130990 642120 131080 642150
rect 131170 642200 131260 642220
rect 131170 642150 131190 642200
rect 131240 642150 131260 642200
rect 131170 642120 131260 642150
rect 124150 642040 131350 642120
rect 131470 642060 131500 642630
rect 131630 642060 131660 642630
rect 131470 642040 131660 642060
rect 123800 642020 123990 642040
rect 127450 641960 128350 642040
rect 127450 641880 127460 641960
rect 128340 641880 128350 641960
rect 127450 641870 128350 641880
rect 115242 641114 115700 641210
rect 102041 640557 102500 640653
rect 102041 639582 102137 640557
rect 115622 640122 115700 641114
rect 115242 640026 115700 640122
rect 102041 639486 102553 639582
rect 102041 639203 102137 639486
rect 102455 638949 102491 639045
rect 115622 639034 115700 640026
rect 119284 640140 119384 640146
rect 119284 640060 119290 640140
rect 119382 640066 119384 640140
rect 119382 640060 119390 640066
rect 119284 640022 119390 640060
rect 119112 639672 119242 639686
rect 119112 639582 119128 639672
rect 119228 639582 119242 639672
rect 119112 639568 119242 639582
rect 119130 639562 119230 639568
rect 119290 639510 119390 640022
rect 120004 639656 120104 639662
rect 120004 639608 120010 639656
rect 119450 639576 120010 639608
rect 120102 639608 120104 639656
rect 120102 639576 120114 639608
rect 119450 639508 120114 639576
rect 115242 638938 115700 639034
rect 115622 638833 115700 638938
rect 115587 638812 115700 638833
rect 115587 638220 115692 638812
rect 120760 638740 121860 638840
rect 115410 638189 115692 638220
rect 115410 638077 115696 638189
rect 115410 637499 115455 638077
rect 115663 637499 115696 638077
rect 115410 637416 115696 637499
rect 121760 636210 121860 638740
rect 126060 636660 126960 636670
rect 126060 636580 126070 636660
rect 126950 636580 126960 636660
rect 126060 636490 126960 636580
rect 124180 636350 128920 636490
rect 124180 636330 124360 636350
rect 124180 636280 124200 636330
rect 124340 636280 124360 636330
rect 124180 636260 124360 636280
rect 124420 636330 124600 636350
rect 124420 636280 124440 636330
rect 124580 636280 124600 636330
rect 124420 636260 124600 636280
rect 124660 636330 124840 636350
rect 124660 636280 124680 636330
rect 124820 636280 124840 636330
rect 124660 636260 124840 636280
rect 124900 636330 125080 636350
rect 124900 636280 124920 636330
rect 125060 636280 125080 636330
rect 124900 636260 125080 636280
rect 125140 636330 125320 636350
rect 125140 636280 125160 636330
rect 125300 636280 125320 636330
rect 125140 636260 125320 636280
rect 125380 636330 125560 636350
rect 125380 636280 125400 636330
rect 125540 636280 125560 636330
rect 125380 636260 125560 636280
rect 125620 636330 125800 636350
rect 125620 636280 125640 636330
rect 125780 636280 125800 636330
rect 125620 636260 125800 636280
rect 125860 636330 126040 636350
rect 125860 636280 125880 636330
rect 126020 636280 126040 636330
rect 125860 636260 126040 636280
rect 126100 636330 126280 636350
rect 126100 636280 126120 636330
rect 126260 636280 126280 636330
rect 126100 636260 126280 636280
rect 126340 636330 126520 636350
rect 126340 636280 126360 636330
rect 126500 636280 126520 636330
rect 126340 636260 126520 636280
rect 126580 636330 126760 636350
rect 126580 636280 126600 636330
rect 126740 636280 126760 636330
rect 126580 636260 126760 636280
rect 126820 636330 127000 636350
rect 126820 636280 126840 636330
rect 126980 636280 127000 636330
rect 126820 636260 127000 636280
rect 127060 636330 127240 636350
rect 127060 636280 127080 636330
rect 127220 636280 127240 636330
rect 127060 636260 127240 636280
rect 127300 636330 127480 636350
rect 127300 636280 127320 636330
rect 127460 636280 127480 636330
rect 127300 636260 127480 636280
rect 127540 636330 127720 636350
rect 127540 636280 127560 636330
rect 127700 636280 127720 636330
rect 127540 636260 127720 636280
rect 127780 636330 127960 636350
rect 127780 636280 127800 636330
rect 127940 636280 127960 636330
rect 127780 636260 127960 636280
rect 128020 636330 128200 636350
rect 128020 636280 128040 636330
rect 128180 636280 128200 636330
rect 128020 636260 128200 636280
rect 128260 636330 128440 636350
rect 128260 636280 128280 636330
rect 128420 636280 128440 636330
rect 128260 636260 128440 636280
rect 128500 636330 128680 636350
rect 128500 636280 128520 636330
rect 128660 636280 128680 636330
rect 128500 636260 128680 636280
rect 128740 636330 128920 636350
rect 128740 636280 128760 636330
rect 128900 636280 128920 636330
rect 128740 636260 128920 636280
rect 129070 636470 129260 636490
rect 121760 636170 124130 636210
rect 121760 636130 124070 636170
rect 124110 636130 124130 636170
rect 121760 636110 124130 636130
rect 124180 636030 124360 636050
rect 124180 635980 124200 636030
rect 124340 635980 124360 636030
rect 124180 635960 124360 635980
rect 124420 636030 124600 636050
rect 124420 635980 124440 636030
rect 124580 635980 124600 636030
rect 124420 635960 124600 635980
rect 124660 636030 124840 636050
rect 124660 635980 124680 636030
rect 124820 635980 124840 636030
rect 124660 635960 124840 635980
rect 124900 636030 125080 636050
rect 124900 635980 124920 636030
rect 125060 635980 125080 636030
rect 124900 635960 125080 635980
rect 125140 636030 125320 636050
rect 125140 635980 125160 636030
rect 125300 635980 125320 636030
rect 125140 635960 125320 635980
rect 125380 636030 125560 636050
rect 125380 635980 125400 636030
rect 125540 635980 125560 636030
rect 125380 635960 125560 635980
rect 125620 636030 125800 636050
rect 125620 635980 125640 636030
rect 125780 635980 125800 636030
rect 125620 635960 125800 635980
rect 125860 636030 126040 636050
rect 125860 635980 125880 636030
rect 126020 635980 126040 636030
rect 125860 635960 126040 635980
rect 126100 636030 126280 636050
rect 126100 635980 126120 636030
rect 126260 635980 126280 636030
rect 126100 635960 126280 635980
rect 126340 636030 126520 636050
rect 126340 635980 126360 636030
rect 126500 635980 126520 636030
rect 126340 635960 126520 635980
rect 126580 636030 126760 636050
rect 126580 635980 126600 636030
rect 126740 635980 126760 636030
rect 126580 635960 126760 635980
rect 126820 636030 127000 636050
rect 126820 635980 126840 636030
rect 126980 635980 127000 636030
rect 126820 635960 127000 635980
rect 127060 636030 127240 636050
rect 127060 635980 127080 636030
rect 127220 635980 127240 636030
rect 127060 635960 127240 635980
rect 127300 636030 127480 636050
rect 127300 635980 127320 636030
rect 127460 635980 127480 636030
rect 127300 635960 127480 635980
rect 127540 636030 127720 636050
rect 127540 635980 127560 636030
rect 127700 635980 127720 636030
rect 127540 635960 127720 635980
rect 127780 636030 127960 636050
rect 127780 635980 127800 636030
rect 127940 635980 127960 636030
rect 127780 635960 127960 635980
rect 128020 636030 128200 636050
rect 128020 635980 128040 636030
rect 128180 635980 128200 636030
rect 128020 635960 128200 635980
rect 128260 636030 128440 636050
rect 128260 635980 128280 636030
rect 128420 635980 128440 636030
rect 128260 635960 128440 635980
rect 128500 636030 128680 636050
rect 128500 635980 128520 636030
rect 128660 635980 128680 636030
rect 128500 635960 128680 635980
rect 128740 636030 128920 636050
rect 128740 635980 128760 636030
rect 128900 635980 128920 636030
rect 128740 635960 128920 635980
rect 124180 635820 128920 635960
rect 129070 635900 129100 636470
rect 129230 635900 129260 636470
rect 129070 635880 129260 635900
rect 126070 635760 126970 635820
rect 126070 635680 126080 635760
rect 126960 635680 126970 635760
rect 126070 635670 126970 635680
rect 119286 633758 119386 633764
rect 119286 633678 119292 633758
rect 119384 633708 119386 633758
rect 119384 633678 119390 633708
rect 119286 633640 119390 633678
rect 119130 633388 119230 633396
rect 119130 633304 119138 633388
rect 119220 633304 119230 633388
rect 119130 633110 119230 633304
rect 119290 633102 119390 633640
rect 119930 633222 120030 633228
rect 119930 633210 119936 633222
rect 119450 633142 119936 633210
rect 120028 633142 120030 633222
rect 119450 633110 120030 633142
rect 119930 633104 120030 633110
rect 124240 632740 124640 632850
rect 124240 632690 124260 632740
rect 124620 632690 124640 632740
rect 124240 632670 124640 632690
rect 124240 632440 124640 632460
rect 120732 632340 123548 632440
rect 123448 630180 123548 632340
rect 124240 632390 124260 632440
rect 124620 632390 124640 632440
rect 124240 632280 124640 632390
rect 126280 630580 127180 630590
rect 126280 630500 126290 630580
rect 127170 630500 127180 630580
rect 126280 630410 127180 630500
rect 129140 630410 129330 630430
rect 124450 630320 128990 630410
rect 124450 630300 124850 630320
rect 124450 630250 124470 630300
rect 124830 630250 124850 630300
rect 124450 630230 124850 630250
rect 124910 630300 125310 630320
rect 124910 630250 124930 630300
rect 125290 630250 125310 630300
rect 124910 630230 125310 630250
rect 125370 630300 125770 630320
rect 125370 630250 125390 630300
rect 125750 630250 125770 630300
rect 125370 630230 125770 630250
rect 125830 630300 126230 630320
rect 125830 630250 125850 630300
rect 126210 630250 126230 630300
rect 125830 630230 126230 630250
rect 126290 630300 126690 630320
rect 126290 630250 126310 630300
rect 126670 630250 126690 630300
rect 126290 630230 126690 630250
rect 126750 630300 127150 630320
rect 126750 630250 126770 630300
rect 127130 630250 127150 630300
rect 126750 630230 127150 630250
rect 127210 630300 127610 630320
rect 127210 630250 127230 630300
rect 127590 630250 127610 630300
rect 127210 630230 127610 630250
rect 127670 630300 128070 630320
rect 127670 630250 127690 630300
rect 128050 630250 128070 630300
rect 127670 630230 128070 630250
rect 128130 630300 128530 630320
rect 128130 630250 128150 630300
rect 128510 630250 128530 630300
rect 128130 630230 128530 630250
rect 128590 630300 128990 630320
rect 128590 630250 128610 630300
rect 128970 630250 128990 630300
rect 128590 630230 128990 630250
rect 123448 630140 124410 630180
rect 123448 630100 124350 630140
rect 124390 630100 124410 630140
rect 123448 630080 124410 630100
rect 124450 630000 124850 630020
rect 124450 629950 124470 630000
rect 124830 629950 124850 630000
rect 124450 629930 124850 629950
rect 124910 630000 125310 630020
rect 124910 629950 124930 630000
rect 125290 629950 125310 630000
rect 124910 629930 125310 629950
rect 125370 630000 125770 630020
rect 125370 629950 125390 630000
rect 125750 629950 125770 630000
rect 125370 629930 125770 629950
rect 125830 630000 126230 630020
rect 125830 629950 125850 630000
rect 126210 629950 126230 630000
rect 125830 629930 126230 629950
rect 126290 630000 126690 630020
rect 126290 629950 126310 630000
rect 126670 629950 126690 630000
rect 126290 629930 126690 629950
rect 126750 630000 127150 630020
rect 126750 629950 126770 630000
rect 127130 629950 127150 630000
rect 126750 629930 127150 629950
rect 127210 630000 127610 630020
rect 127210 629950 127230 630000
rect 127590 629950 127610 630000
rect 127210 629930 127610 629950
rect 127670 630000 128070 630020
rect 127670 629950 127690 630000
rect 128050 629950 128070 630000
rect 127670 629930 128070 629950
rect 128130 630000 128530 630020
rect 128130 629950 128150 630000
rect 128510 629950 128530 630000
rect 128130 629930 128530 629950
rect 128590 630000 128990 630020
rect 128590 629950 128610 630000
rect 128970 629950 128990 630000
rect 128590 629930 128990 629950
rect 124450 629840 128990 629930
rect 129140 629840 129170 630410
rect 129300 629840 129330 630410
rect 126210 629830 127250 629840
rect 126280 629770 127180 629830
rect 129140 629820 129330 629840
rect 126280 629690 126290 629770
rect 127170 629690 127180 629770
rect 126280 629680 127180 629690
rect 119302 627220 119402 627226
rect 119302 627186 119308 627220
rect 119290 627140 119308 627186
rect 119400 627140 119402 627220
rect 119290 627102 119402 627140
rect 119128 626890 119228 626898
rect 119128 626806 119136 626890
rect 119218 626806 119228 626890
rect 119128 626792 119228 626806
rect 119290 626710 119390 627102
rect 119450 626788 120006 626810
rect 119450 626782 120012 626788
rect 119450 626710 119918 626782
rect 119912 626702 119918 626710
rect 120010 626702 120012 626782
rect 119912 626664 120012 626702
rect 120740 625940 123478 626040
rect 123378 624042 123478 625940
rect 124220 625070 124820 625180
rect 124220 625020 124240 625070
rect 124800 625020 124820 625070
rect 124220 625000 124820 625020
rect 124220 624770 124820 624790
rect 124220 624720 124240 624770
rect 124800 624720 124820 624770
rect 124220 624610 124820 624720
rect 126530 624060 127430 624070
rect 123378 624040 124256 624042
rect 123378 624010 124660 624040
rect 123378 623970 124600 624010
rect 124640 623970 124660 624010
rect 123378 623942 124660 623970
rect 124250 623940 124660 623942
rect 126530 623980 126540 624060
rect 127420 623980 127430 624060
rect 126530 623890 127430 623980
rect 128790 623890 128980 623910
rect 124780 623780 128680 623890
rect 124780 623730 124800 623780
rect 125360 623730 125460 623780
rect 126020 623730 126120 623780
rect 126680 623730 126780 623780
rect 127340 623730 127440 623780
rect 128000 623730 128100 623780
rect 128660 623730 128680 623780
rect 124780 623710 128680 623730
rect 124780 623480 128680 623500
rect 124780 623430 124800 623480
rect 125360 623430 125460 623480
rect 126020 623430 126120 623480
rect 126680 623430 126780 623480
rect 127340 623430 127440 623480
rect 128000 623430 128100 623480
rect 128660 623430 128680 623480
rect 124780 623320 128680 623430
rect 128790 623320 128820 623890
rect 128950 623320 128980 623890
rect 126530 623250 127430 623320
rect 128790 623300 128980 623320
rect 126530 623170 126540 623250
rect 127420 623170 127430 623250
rect 126530 623160 127430 623170
rect 119290 620844 119390 620850
rect 119290 620764 119296 620844
rect 119388 620764 119390 620844
rect 119134 620484 119234 620492
rect 119134 620400 119142 620484
rect 119224 620400 119234 620484
rect 119134 620386 119234 620400
rect 119290 620304 119390 620764
rect 119450 620380 120010 620400
rect 119450 620374 120044 620380
rect 119450 620300 119950 620374
rect 119944 620294 119950 620300
rect 120042 620294 120044 620374
rect 119944 620256 120044 620294
rect 120760 619540 124342 619640
rect 124242 618834 124342 619540
rect 125300 619400 125720 619460
rect 125460 619370 125520 619400
rect 125350 619350 125410 619370
rect 125350 619310 125360 619350
rect 125400 619310 125410 619350
rect 125350 619180 125410 619310
rect 125450 619350 125530 619370
rect 125450 619310 125470 619350
rect 125510 619310 125530 619350
rect 125450 619290 125530 619310
rect 125570 619350 125630 619370
rect 125570 619310 125580 619350
rect 125620 619310 125630 619350
rect 125570 619180 125630 619310
rect 124242 618770 131768 618834
rect 124242 618734 125590 618770
rect 125580 618730 125590 618734
rect 125630 618734 125930 618770
rect 125630 618730 125640 618734
rect 125580 618710 125640 618730
rect 125920 618730 125930 618734
rect 125970 618734 126270 618770
rect 125970 618730 125980 618734
rect 125920 618710 125980 618730
rect 126260 618730 126270 618734
rect 126310 618734 126610 618770
rect 126310 618730 126320 618734
rect 126260 618710 126320 618730
rect 126600 618730 126610 618734
rect 126650 618734 126950 618770
rect 126650 618730 126660 618734
rect 126600 618710 126660 618730
rect 126940 618730 126950 618734
rect 126990 618734 127290 618770
rect 126990 618730 127000 618734
rect 126940 618710 127000 618730
rect 127280 618730 127290 618734
rect 127330 618734 127630 618770
rect 127330 618730 127340 618734
rect 127280 618710 127340 618730
rect 127620 618730 127630 618734
rect 127670 618734 127970 618770
rect 127670 618730 127680 618734
rect 127620 618710 127680 618730
rect 127960 618730 127970 618734
rect 128010 618734 128310 618770
rect 128010 618730 128020 618734
rect 127960 618710 128020 618730
rect 128300 618730 128310 618734
rect 128350 618734 128650 618770
rect 128350 618730 128360 618734
rect 128300 618710 128360 618730
rect 128640 618730 128650 618734
rect 128690 618734 128990 618770
rect 128690 618730 128700 618734
rect 128640 618710 128700 618730
rect 128980 618730 128990 618734
rect 129030 618734 129330 618770
rect 129030 618730 129040 618734
rect 128980 618710 129040 618730
rect 129320 618730 129330 618734
rect 129370 618734 129670 618770
rect 129370 618730 129380 618734
rect 129320 618710 129380 618730
rect 129660 618730 129670 618734
rect 129710 618734 130010 618770
rect 129710 618730 129720 618734
rect 129660 618710 129720 618730
rect 130000 618730 130010 618734
rect 130050 618734 130350 618770
rect 130050 618730 130060 618734
rect 130000 618710 130060 618730
rect 130340 618730 130350 618734
rect 130390 618734 130690 618770
rect 130390 618730 130400 618734
rect 130340 618710 130400 618730
rect 130680 618730 130690 618734
rect 130730 618734 131030 618770
rect 130730 618730 130740 618734
rect 130680 618710 130740 618730
rect 131020 618730 131030 618734
rect 131070 618734 131370 618770
rect 131070 618730 131080 618734
rect 131020 618710 131080 618730
rect 131360 618730 131370 618734
rect 131410 618734 131710 618770
rect 131410 618730 131420 618734
rect 131360 618710 131420 618730
rect 131700 618730 131710 618734
rect 131750 618734 131768 618770
rect 131910 618810 132100 618830
rect 131750 618730 131760 618734
rect 131700 618710 131760 618730
rect 125360 618620 128380 618680
rect 128860 618620 131820 618680
rect 125530 618590 125590 618620
rect 125870 618590 125930 618620
rect 126210 618590 126270 618620
rect 126550 618590 126610 618620
rect 126890 618590 126950 618620
rect 127230 618590 127290 618620
rect 127570 618590 127630 618620
rect 127910 618590 127970 618620
rect 128250 618590 128310 618620
rect 128590 618590 128650 618620
rect 128930 618590 128990 618620
rect 129270 618590 129330 618620
rect 129610 618590 129670 618620
rect 129950 618590 130010 618620
rect 130290 618590 130350 618620
rect 130630 618590 130690 618620
rect 130970 618590 131030 618620
rect 131310 618590 131370 618620
rect 131650 618590 131710 618620
rect 125420 618570 125480 618590
rect 125420 618530 125430 618570
rect 125470 618530 125480 618570
rect 125420 618460 125480 618530
rect 125520 618570 125600 618590
rect 125520 618530 125540 618570
rect 125580 618530 125600 618570
rect 125520 618510 125600 618530
rect 125640 618570 125700 618590
rect 125640 618530 125650 618570
rect 125690 618530 125700 618570
rect 125640 618460 125700 618530
rect 125760 618570 125820 618590
rect 125760 618530 125770 618570
rect 125810 618530 125820 618570
rect 125760 618460 125820 618530
rect 125860 618570 125940 618590
rect 125860 618530 125880 618570
rect 125920 618530 125940 618570
rect 125860 618510 125940 618530
rect 125980 618570 126040 618590
rect 125980 618530 125990 618570
rect 126030 618530 126040 618570
rect 125980 618460 126040 618530
rect 126100 618570 126160 618590
rect 126100 618530 126110 618570
rect 126150 618530 126160 618570
rect 126100 618460 126160 618530
rect 126200 618570 126280 618590
rect 126200 618530 126220 618570
rect 126260 618530 126280 618570
rect 126200 618510 126280 618530
rect 126320 618570 126380 618590
rect 126320 618530 126330 618570
rect 126370 618530 126380 618570
rect 126320 618460 126380 618530
rect 126440 618570 126500 618590
rect 126440 618530 126450 618570
rect 126490 618530 126500 618570
rect 126440 618460 126500 618530
rect 126540 618570 126620 618590
rect 126540 618530 126560 618570
rect 126600 618530 126620 618570
rect 126540 618510 126620 618530
rect 126660 618570 126720 618590
rect 126660 618530 126670 618570
rect 126710 618530 126720 618570
rect 126660 618460 126720 618530
rect 126780 618570 126840 618590
rect 126780 618530 126790 618570
rect 126830 618530 126840 618570
rect 126780 618460 126840 618530
rect 126880 618570 126960 618590
rect 126880 618530 126900 618570
rect 126940 618530 126960 618570
rect 126880 618510 126960 618530
rect 127000 618570 127060 618590
rect 127000 618530 127010 618570
rect 127050 618530 127060 618570
rect 127000 618460 127060 618530
rect 127120 618570 127180 618590
rect 127120 618530 127130 618570
rect 127170 618530 127180 618570
rect 127120 618460 127180 618530
rect 127220 618570 127300 618590
rect 127220 618530 127240 618570
rect 127280 618530 127300 618570
rect 127220 618510 127300 618530
rect 127340 618570 127400 618590
rect 127340 618530 127350 618570
rect 127390 618530 127400 618570
rect 127340 618460 127400 618530
rect 127460 618570 127520 618590
rect 127460 618530 127470 618570
rect 127510 618530 127520 618570
rect 127460 618460 127520 618530
rect 127560 618570 127640 618590
rect 127560 618530 127580 618570
rect 127620 618530 127640 618570
rect 127560 618510 127640 618530
rect 127680 618570 127740 618590
rect 127680 618530 127690 618570
rect 127730 618530 127740 618570
rect 127680 618460 127740 618530
rect 127800 618570 127860 618590
rect 127800 618530 127810 618570
rect 127850 618530 127860 618570
rect 127800 618460 127860 618530
rect 127900 618570 127980 618590
rect 127900 618530 127920 618570
rect 127960 618530 127980 618570
rect 127900 618510 127980 618530
rect 128020 618570 128080 618590
rect 128020 618530 128030 618570
rect 128070 618530 128080 618570
rect 128020 618460 128080 618530
rect 128140 618570 128200 618590
rect 128140 618530 128150 618570
rect 128190 618530 128200 618570
rect 128140 618460 128200 618530
rect 128240 618570 128320 618590
rect 128240 618530 128260 618570
rect 128300 618530 128320 618570
rect 128240 618510 128320 618530
rect 128360 618570 128420 618590
rect 128360 618530 128370 618570
rect 128410 618530 128420 618570
rect 128360 618460 128420 618530
rect 128480 618570 128540 618590
rect 128480 618530 128490 618570
rect 128530 618530 128540 618570
rect 128480 618460 128540 618530
rect 128580 618570 128660 618590
rect 128580 618530 128600 618570
rect 128640 618530 128660 618570
rect 128580 618510 128660 618530
rect 128700 618570 128760 618590
rect 128700 618530 128710 618570
rect 128750 618530 128760 618570
rect 128700 618460 128760 618530
rect 128820 618570 128880 618590
rect 128820 618530 128830 618570
rect 128870 618530 128880 618570
rect 128820 618460 128880 618530
rect 128920 618570 129000 618590
rect 128920 618530 128940 618570
rect 128980 618530 129000 618570
rect 128920 618510 129000 618530
rect 129040 618570 129100 618590
rect 129040 618530 129050 618570
rect 129090 618530 129100 618570
rect 129040 618460 129100 618530
rect 129160 618570 129220 618590
rect 129160 618530 129170 618570
rect 129210 618530 129220 618570
rect 129160 618460 129220 618530
rect 129260 618570 129340 618590
rect 129260 618530 129280 618570
rect 129320 618530 129340 618570
rect 129260 618510 129340 618530
rect 129380 618570 129440 618590
rect 129380 618530 129390 618570
rect 129430 618530 129440 618570
rect 129380 618460 129440 618530
rect 129500 618570 129560 618590
rect 129500 618530 129510 618570
rect 129550 618530 129560 618570
rect 129500 618460 129560 618530
rect 129600 618570 129680 618590
rect 129600 618530 129620 618570
rect 129660 618530 129680 618570
rect 129600 618510 129680 618530
rect 129720 618570 129780 618590
rect 129720 618530 129730 618570
rect 129770 618530 129780 618570
rect 129720 618460 129780 618530
rect 129840 618570 129900 618590
rect 129840 618530 129850 618570
rect 129890 618530 129900 618570
rect 129840 618460 129900 618530
rect 129940 618570 130020 618590
rect 129940 618530 129960 618570
rect 130000 618530 130020 618570
rect 129940 618510 130020 618530
rect 130060 618570 130120 618590
rect 130060 618530 130070 618570
rect 130110 618530 130120 618570
rect 130060 618460 130120 618530
rect 130180 618570 130240 618590
rect 130180 618530 130190 618570
rect 130230 618530 130240 618570
rect 130180 618460 130240 618530
rect 130280 618570 130360 618590
rect 130280 618530 130300 618570
rect 130340 618530 130360 618570
rect 130280 618510 130360 618530
rect 130400 618570 130460 618590
rect 130400 618530 130410 618570
rect 130450 618530 130460 618570
rect 130400 618460 130460 618530
rect 130520 618570 130580 618590
rect 130520 618530 130530 618570
rect 130570 618530 130580 618570
rect 130520 618460 130580 618530
rect 130620 618570 130700 618590
rect 130620 618530 130640 618570
rect 130680 618530 130700 618570
rect 130620 618510 130700 618530
rect 130740 618570 130800 618590
rect 130740 618530 130750 618570
rect 130790 618530 130800 618570
rect 130740 618460 130800 618530
rect 130860 618570 130920 618590
rect 130860 618530 130870 618570
rect 130910 618530 130920 618570
rect 130860 618460 130920 618530
rect 130960 618570 131040 618590
rect 130960 618530 130980 618570
rect 131020 618530 131040 618570
rect 130960 618510 131040 618530
rect 131080 618570 131140 618590
rect 131080 618530 131090 618570
rect 131130 618530 131140 618570
rect 131080 618460 131140 618530
rect 131200 618570 131260 618590
rect 131200 618530 131210 618570
rect 131250 618530 131260 618570
rect 131200 618460 131260 618530
rect 131300 618570 131380 618590
rect 131300 618530 131320 618570
rect 131360 618530 131380 618570
rect 131300 618510 131380 618530
rect 131420 618570 131480 618590
rect 131420 618530 131430 618570
rect 131470 618530 131480 618570
rect 131420 618460 131480 618530
rect 131540 618570 131600 618590
rect 131540 618530 131550 618570
rect 131590 618530 131600 618570
rect 131540 618460 131600 618530
rect 131640 618570 131720 618590
rect 131640 618530 131660 618570
rect 131700 618530 131720 618570
rect 131640 618510 131720 618530
rect 131760 618570 131820 618590
rect 131760 618530 131770 618570
rect 131810 618530 131820 618570
rect 131760 618460 131820 618530
rect 125420 618400 128380 618460
rect 128860 618400 131820 618460
rect 131910 618240 131940 618810
rect 132070 618240 132100 618810
rect 131910 618220 132100 618240
rect 119298 614364 119398 614370
rect 119298 614324 119304 614364
rect 119290 614284 119304 614324
rect 119396 614284 119398 614364
rect 119290 614246 119398 614284
rect 119134 614058 119234 614066
rect 119134 613974 119142 614058
rect 119224 613974 119234 614058
rect 119134 613960 119234 613974
rect 119290 613902 119390 614246
rect 119450 613974 120012 614002
rect 119450 613968 120072 613974
rect 119450 613902 119978 613968
rect 119972 613888 119978 613902
rect 120070 613888 120072 613968
rect 119972 613850 120072 613888
rect 120578 613140 123992 613240
rect 123892 611384 123992 613140
rect 124950 611950 125370 612010
rect 125110 611920 125170 611950
rect 125000 611900 125060 611920
rect 125000 611860 125010 611900
rect 125050 611860 125060 611900
rect 125000 611730 125060 611860
rect 125100 611900 125180 611920
rect 125100 611860 125120 611900
rect 125160 611860 125180 611900
rect 125100 611840 125180 611860
rect 125220 611900 125280 611920
rect 125220 611860 125230 611900
rect 125270 611860 125280 611900
rect 125220 611730 125280 611860
rect 123892 611320 131418 611384
rect 123892 611284 125240 611320
rect 125230 611280 125240 611284
rect 125280 611284 125580 611320
rect 125280 611280 125290 611284
rect 125230 611260 125290 611280
rect 125570 611280 125580 611284
rect 125620 611284 125920 611320
rect 125620 611280 125630 611284
rect 125570 611260 125630 611280
rect 125910 611280 125920 611284
rect 125960 611284 126260 611320
rect 125960 611280 125970 611284
rect 125910 611260 125970 611280
rect 126250 611280 126260 611284
rect 126300 611284 126600 611320
rect 126300 611280 126310 611284
rect 126250 611260 126310 611280
rect 126590 611280 126600 611284
rect 126640 611284 126940 611320
rect 126640 611280 126650 611284
rect 126590 611260 126650 611280
rect 126930 611280 126940 611284
rect 126980 611284 127280 611320
rect 126980 611280 126990 611284
rect 126930 611260 126990 611280
rect 127270 611280 127280 611284
rect 127320 611284 127620 611320
rect 127320 611280 127330 611284
rect 127270 611260 127330 611280
rect 127610 611280 127620 611284
rect 127660 611284 127960 611320
rect 127660 611280 127670 611284
rect 127610 611260 127670 611280
rect 127950 611280 127960 611284
rect 128000 611284 128300 611320
rect 128000 611280 128010 611284
rect 127950 611260 128010 611280
rect 128290 611280 128300 611284
rect 128340 611284 128640 611320
rect 128340 611280 128350 611284
rect 128290 611260 128350 611280
rect 128630 611280 128640 611284
rect 128680 611284 128980 611320
rect 128680 611280 128690 611284
rect 128630 611260 128690 611280
rect 128970 611280 128980 611284
rect 129020 611284 129320 611320
rect 129020 611280 129030 611284
rect 128970 611260 129030 611280
rect 129310 611280 129320 611284
rect 129360 611284 129660 611320
rect 129360 611280 129370 611284
rect 129310 611260 129370 611280
rect 129650 611280 129660 611284
rect 129700 611284 130000 611320
rect 129700 611280 129710 611284
rect 129650 611260 129710 611280
rect 129990 611280 130000 611284
rect 130040 611284 130340 611320
rect 130040 611280 130050 611284
rect 129990 611260 130050 611280
rect 130330 611280 130340 611284
rect 130380 611284 130680 611320
rect 130380 611280 130390 611284
rect 130330 611260 130390 611280
rect 130670 611280 130680 611284
rect 130720 611284 131020 611320
rect 130720 611280 130730 611284
rect 130670 611260 130730 611280
rect 131010 611280 131020 611284
rect 131060 611284 131360 611320
rect 131060 611280 131070 611284
rect 131010 611260 131070 611280
rect 131350 611280 131360 611284
rect 131400 611284 131418 611320
rect 131560 611360 131750 611380
rect 131400 611280 131410 611284
rect 131350 611260 131410 611280
rect 125010 611170 128030 611230
rect 128510 611170 131470 611230
rect 125180 611140 125240 611170
rect 125520 611140 125580 611170
rect 125860 611140 125920 611170
rect 126200 611140 126260 611170
rect 126540 611140 126600 611170
rect 126880 611140 126940 611170
rect 127220 611140 127280 611170
rect 127560 611140 127620 611170
rect 127900 611140 127960 611170
rect 128240 611140 128300 611170
rect 128580 611140 128640 611170
rect 128920 611140 128980 611170
rect 129260 611140 129320 611170
rect 129600 611140 129660 611170
rect 129940 611140 130000 611170
rect 130280 611140 130340 611170
rect 130620 611140 130680 611170
rect 130960 611140 131020 611170
rect 131300 611140 131360 611170
rect 125070 611120 125130 611140
rect 125070 610930 125080 611120
rect 125120 610930 125130 611120
rect 125070 610860 125130 610930
rect 125170 611120 125250 611140
rect 125170 610930 125190 611120
rect 125230 610930 125250 611120
rect 125170 610910 125250 610930
rect 125290 611120 125350 611140
rect 125290 610930 125300 611120
rect 125340 610930 125350 611120
rect 125290 610860 125350 610930
rect 125410 611120 125470 611140
rect 125410 610930 125420 611120
rect 125460 610930 125470 611120
rect 125410 610860 125470 610930
rect 125510 611120 125590 611140
rect 125510 610930 125530 611120
rect 125570 610930 125590 611120
rect 125510 610910 125590 610930
rect 125630 611120 125690 611140
rect 125630 610930 125640 611120
rect 125680 610930 125690 611120
rect 125630 610860 125690 610930
rect 125750 611120 125810 611140
rect 125750 610930 125760 611120
rect 125800 610930 125810 611120
rect 125750 610860 125810 610930
rect 125850 611120 125930 611140
rect 125850 610930 125870 611120
rect 125910 610930 125930 611120
rect 125850 610910 125930 610930
rect 125970 611120 126030 611140
rect 125970 610930 125980 611120
rect 126020 610930 126030 611120
rect 125970 610860 126030 610930
rect 126090 611120 126150 611140
rect 126090 610930 126100 611120
rect 126140 610930 126150 611120
rect 126090 610860 126150 610930
rect 126190 611120 126270 611140
rect 126190 610930 126210 611120
rect 126250 610930 126270 611120
rect 126190 610910 126270 610930
rect 126310 611120 126370 611140
rect 126310 610930 126320 611120
rect 126360 610930 126370 611120
rect 126310 610860 126370 610930
rect 126430 611120 126490 611140
rect 126430 610930 126440 611120
rect 126480 610930 126490 611120
rect 126430 610860 126490 610930
rect 126530 611120 126610 611140
rect 126530 610930 126550 611120
rect 126590 610930 126610 611120
rect 126530 610910 126610 610930
rect 126650 611120 126710 611140
rect 126650 610930 126660 611120
rect 126700 610930 126710 611120
rect 126650 610860 126710 610930
rect 126770 611120 126830 611140
rect 126770 610930 126780 611120
rect 126820 610930 126830 611120
rect 126770 610860 126830 610930
rect 126870 611120 126950 611140
rect 126870 610930 126890 611120
rect 126930 610930 126950 611120
rect 126870 610910 126950 610930
rect 126990 611120 127050 611140
rect 126990 610930 127000 611120
rect 127040 610930 127050 611120
rect 126990 610860 127050 610930
rect 127110 611120 127170 611140
rect 127110 610930 127120 611120
rect 127160 610930 127170 611120
rect 127110 610860 127170 610930
rect 127210 611120 127290 611140
rect 127210 610930 127230 611120
rect 127270 610930 127290 611120
rect 127210 610910 127290 610930
rect 127330 611120 127390 611140
rect 127330 610930 127340 611120
rect 127380 610930 127390 611120
rect 127330 610860 127390 610930
rect 127450 611120 127510 611140
rect 127450 610930 127460 611120
rect 127500 610930 127510 611120
rect 127450 610860 127510 610930
rect 127550 611120 127630 611140
rect 127550 610930 127570 611120
rect 127610 610930 127630 611120
rect 127550 610910 127630 610930
rect 127670 611120 127730 611140
rect 127670 610930 127680 611120
rect 127720 610930 127730 611120
rect 127670 610860 127730 610930
rect 127790 611120 127850 611140
rect 127790 610930 127800 611120
rect 127840 610930 127850 611120
rect 127790 610860 127850 610930
rect 127890 611120 127970 611140
rect 127890 610930 127910 611120
rect 127950 610930 127970 611120
rect 127890 610910 127970 610930
rect 128010 611120 128070 611140
rect 128010 610930 128020 611120
rect 128060 610930 128070 611120
rect 128010 610860 128070 610930
rect 128130 611120 128190 611140
rect 128130 610930 128140 611120
rect 128180 610930 128190 611120
rect 128130 610860 128190 610930
rect 128230 611120 128310 611140
rect 128230 610930 128250 611120
rect 128290 610930 128310 611120
rect 128230 610910 128310 610930
rect 128350 611120 128410 611140
rect 128350 610930 128360 611120
rect 128400 610930 128410 611120
rect 128350 610860 128410 610930
rect 128470 611120 128530 611140
rect 128470 610930 128480 611120
rect 128520 610930 128530 611120
rect 128470 610860 128530 610930
rect 128570 611120 128650 611140
rect 128570 610930 128590 611120
rect 128630 610930 128650 611120
rect 128570 610910 128650 610930
rect 128690 611120 128750 611140
rect 128690 610930 128700 611120
rect 128740 610930 128750 611120
rect 128690 610860 128750 610930
rect 128810 611120 128870 611140
rect 128810 610930 128820 611120
rect 128860 610930 128870 611120
rect 128810 610860 128870 610930
rect 128910 611120 128990 611140
rect 128910 610930 128930 611120
rect 128970 610930 128990 611120
rect 128910 610910 128990 610930
rect 129030 611120 129090 611140
rect 129030 610930 129040 611120
rect 129080 610930 129090 611120
rect 129030 610860 129090 610930
rect 129150 611120 129210 611140
rect 129150 610930 129160 611120
rect 129200 610930 129210 611120
rect 129150 610860 129210 610930
rect 129250 611120 129330 611140
rect 129250 610930 129270 611120
rect 129310 610930 129330 611120
rect 129250 610910 129330 610930
rect 129370 611120 129430 611140
rect 129370 610930 129380 611120
rect 129420 610930 129430 611120
rect 129370 610860 129430 610930
rect 129490 611120 129550 611140
rect 129490 610930 129500 611120
rect 129540 610930 129550 611120
rect 129490 610860 129550 610930
rect 129590 611120 129670 611140
rect 129590 610930 129610 611120
rect 129650 610930 129670 611120
rect 129590 610910 129670 610930
rect 129710 611120 129770 611140
rect 129710 610930 129720 611120
rect 129760 610930 129770 611120
rect 129710 610860 129770 610930
rect 129830 611120 129890 611140
rect 129830 610930 129840 611120
rect 129880 610930 129890 611120
rect 129830 610860 129890 610930
rect 129930 611120 130010 611140
rect 129930 610930 129950 611120
rect 129990 610930 130010 611120
rect 129930 610910 130010 610930
rect 130050 611120 130110 611140
rect 130050 610930 130060 611120
rect 130100 610930 130110 611120
rect 130050 610860 130110 610930
rect 130170 611120 130230 611140
rect 130170 610930 130180 611120
rect 130220 610930 130230 611120
rect 130170 610860 130230 610930
rect 130270 611120 130350 611140
rect 130270 610930 130290 611120
rect 130330 610930 130350 611120
rect 130270 610910 130350 610930
rect 130390 611120 130450 611140
rect 130390 610930 130400 611120
rect 130440 610930 130450 611120
rect 130390 610860 130450 610930
rect 130510 611120 130570 611140
rect 130510 610930 130520 611120
rect 130560 610930 130570 611120
rect 130510 610860 130570 610930
rect 130610 611120 130690 611140
rect 130610 610930 130630 611120
rect 130670 610930 130690 611120
rect 130610 610910 130690 610930
rect 130730 611120 130790 611140
rect 130730 610930 130740 611120
rect 130780 610930 130790 611120
rect 130730 610860 130790 610930
rect 130850 611120 130910 611140
rect 130850 610930 130860 611120
rect 130900 610930 130910 611120
rect 130850 610860 130910 610930
rect 130950 611120 131030 611140
rect 130950 610930 130970 611120
rect 131010 610930 131030 611120
rect 130950 610910 131030 610930
rect 131070 611120 131130 611140
rect 131070 610930 131080 611120
rect 131120 610930 131130 611120
rect 131070 610860 131130 610930
rect 131190 611120 131250 611140
rect 131190 610930 131200 611120
rect 131240 610930 131250 611120
rect 131190 610860 131250 610930
rect 131290 611120 131370 611140
rect 131290 610930 131310 611120
rect 131350 610930 131370 611120
rect 131290 610910 131370 610930
rect 131410 611120 131470 611140
rect 131410 610930 131420 611120
rect 131460 610930 131470 611120
rect 131410 610860 131470 610930
rect 125070 610800 128030 610860
rect 128510 610800 131470 610860
rect 131560 610790 131590 611360
rect 131720 610790 131750 611360
rect 131560 610770 131750 610790
rect 119302 608058 119402 608064
rect 119302 608002 119308 608058
rect 119290 607978 119308 608002
rect 119400 607978 119402 608058
rect 119290 607940 119402 607978
rect 119130 607676 119230 607684
rect 119130 607592 119138 607676
rect 119220 607592 119230 607676
rect 119130 607578 119230 607592
rect 119290 607502 119390 607940
rect 119450 607566 119974 607610
rect 119450 607560 120008 607566
rect 119450 607510 119914 607560
rect 119908 607480 119914 607510
rect 120006 607480 120008 607560
rect 119908 607442 120008 607480
rect 120626 606740 124122 606840
rect 124022 606140 124122 606740
rect 124020 606040 124122 606140
rect 124022 605334 124122 606040
rect 125080 605900 125500 605960
rect 125240 605870 125300 605900
rect 125130 605850 125190 605870
rect 125130 605810 125140 605850
rect 125180 605810 125190 605850
rect 125130 605680 125190 605810
rect 125230 605850 125310 605870
rect 125230 605810 125250 605850
rect 125290 605810 125310 605850
rect 125230 605790 125310 605810
rect 125350 605850 125410 605870
rect 125350 605810 125360 605850
rect 125400 605810 125410 605850
rect 125350 605680 125410 605810
rect 124022 605270 131548 605334
rect 124022 605234 125370 605270
rect 125360 605230 125370 605234
rect 125410 605234 125710 605270
rect 125410 605230 125420 605234
rect 125360 605210 125420 605230
rect 125700 605230 125710 605234
rect 125750 605234 126050 605270
rect 125750 605230 125760 605234
rect 125700 605210 125760 605230
rect 126040 605230 126050 605234
rect 126090 605234 126390 605270
rect 126090 605230 126100 605234
rect 126040 605210 126100 605230
rect 126380 605230 126390 605234
rect 126430 605234 126730 605270
rect 126430 605230 126440 605234
rect 126380 605210 126440 605230
rect 126720 605230 126730 605234
rect 126770 605234 127070 605270
rect 126770 605230 126780 605234
rect 126720 605210 126780 605230
rect 127060 605230 127070 605234
rect 127110 605234 127410 605270
rect 127110 605230 127120 605234
rect 127060 605210 127120 605230
rect 127400 605230 127410 605234
rect 127450 605234 127750 605270
rect 127450 605230 127460 605234
rect 127400 605210 127460 605230
rect 127740 605230 127750 605234
rect 127790 605234 128090 605270
rect 127790 605230 127800 605234
rect 127740 605210 127800 605230
rect 128080 605230 128090 605234
rect 128130 605234 128430 605270
rect 128130 605230 128140 605234
rect 128080 605210 128140 605230
rect 128420 605230 128430 605234
rect 128470 605234 128770 605270
rect 128470 605230 128480 605234
rect 128420 605210 128480 605230
rect 128760 605230 128770 605234
rect 128810 605234 129110 605270
rect 128810 605230 128820 605234
rect 128760 605210 128820 605230
rect 129100 605230 129110 605234
rect 129150 605234 129450 605270
rect 129150 605230 129160 605234
rect 129100 605210 129160 605230
rect 129440 605230 129450 605234
rect 129490 605234 129790 605270
rect 129490 605230 129500 605234
rect 129440 605210 129500 605230
rect 129780 605230 129790 605234
rect 129830 605234 130130 605270
rect 129830 605230 129840 605234
rect 129780 605210 129840 605230
rect 130120 605230 130130 605234
rect 130170 605234 130470 605270
rect 130170 605230 130180 605234
rect 130120 605210 130180 605230
rect 130460 605230 130470 605234
rect 130510 605234 130810 605270
rect 130510 605230 130520 605234
rect 130460 605210 130520 605230
rect 130800 605230 130810 605234
rect 130850 605234 131150 605270
rect 130850 605230 130860 605234
rect 130800 605210 130860 605230
rect 131140 605230 131150 605234
rect 131190 605234 131490 605270
rect 131190 605230 131200 605234
rect 131140 605210 131200 605230
rect 131480 605230 131490 605234
rect 131530 605234 131548 605270
rect 131690 605310 131880 605330
rect 131530 605230 131540 605234
rect 131480 605210 131540 605230
rect 125140 605120 128160 605180
rect 128640 605120 131600 605180
rect 125310 605090 125370 605120
rect 125650 605090 125710 605120
rect 125990 605090 126050 605120
rect 126330 605090 126390 605120
rect 126670 605090 126730 605120
rect 127010 605090 127070 605120
rect 127350 605090 127410 605120
rect 127690 605090 127750 605120
rect 128030 605090 128090 605120
rect 128370 605090 128430 605120
rect 128710 605090 128770 605120
rect 129050 605090 129110 605120
rect 129390 605090 129450 605120
rect 129730 605090 129790 605120
rect 130070 605090 130130 605120
rect 130410 605090 130470 605120
rect 130750 605090 130810 605120
rect 131090 605090 131150 605120
rect 131430 605090 131490 605120
rect 125200 605070 125260 605090
rect 125200 604780 125210 605070
rect 125250 604780 125260 605070
rect 125200 604710 125260 604780
rect 125300 605070 125380 605090
rect 125300 604780 125320 605070
rect 125360 604780 125380 605070
rect 125300 604760 125380 604780
rect 125420 605070 125480 605090
rect 125420 604780 125430 605070
rect 125470 604780 125480 605070
rect 125420 604710 125480 604780
rect 125540 605070 125600 605090
rect 125540 604780 125550 605070
rect 125590 604780 125600 605070
rect 125540 604710 125600 604780
rect 125640 605070 125720 605090
rect 125640 604780 125660 605070
rect 125700 604780 125720 605070
rect 125640 604760 125720 604780
rect 125760 605070 125820 605090
rect 125760 604780 125770 605070
rect 125810 604780 125820 605070
rect 125760 604710 125820 604780
rect 125880 605070 125940 605090
rect 125880 604780 125890 605070
rect 125930 604780 125940 605070
rect 125880 604710 125940 604780
rect 125980 605070 126060 605090
rect 125980 604780 126000 605070
rect 126040 604780 126060 605070
rect 125980 604760 126060 604780
rect 126100 605070 126160 605090
rect 126100 604780 126110 605070
rect 126150 604780 126160 605070
rect 126100 604710 126160 604780
rect 126220 605070 126280 605090
rect 126220 604780 126230 605070
rect 126270 604780 126280 605070
rect 126220 604710 126280 604780
rect 126320 605070 126400 605090
rect 126320 604780 126340 605070
rect 126380 604780 126400 605070
rect 126320 604760 126400 604780
rect 126440 605070 126500 605090
rect 126440 604780 126450 605070
rect 126490 604780 126500 605070
rect 126440 604710 126500 604780
rect 126560 605070 126620 605090
rect 126560 604780 126570 605070
rect 126610 604780 126620 605070
rect 126560 604710 126620 604780
rect 126660 605070 126740 605090
rect 126660 604780 126680 605070
rect 126720 604780 126740 605070
rect 126660 604760 126740 604780
rect 126780 605070 126840 605090
rect 126780 604780 126790 605070
rect 126830 604780 126840 605070
rect 126780 604710 126840 604780
rect 126900 605070 126960 605090
rect 126900 604780 126910 605070
rect 126950 604780 126960 605070
rect 126900 604710 126960 604780
rect 127000 605070 127080 605090
rect 127000 604780 127020 605070
rect 127060 604780 127080 605070
rect 127000 604760 127080 604780
rect 127120 605070 127180 605090
rect 127120 604780 127130 605070
rect 127170 604780 127180 605070
rect 127120 604710 127180 604780
rect 127240 605070 127300 605090
rect 127240 604780 127250 605070
rect 127290 604780 127300 605070
rect 127240 604710 127300 604780
rect 127340 605070 127420 605090
rect 127340 604780 127360 605070
rect 127400 604780 127420 605070
rect 127340 604760 127420 604780
rect 127460 605070 127520 605090
rect 127460 604780 127470 605070
rect 127510 604780 127520 605070
rect 127460 604710 127520 604780
rect 127580 605070 127640 605090
rect 127580 604780 127590 605070
rect 127630 604780 127640 605070
rect 127580 604710 127640 604780
rect 127680 605070 127760 605090
rect 127680 604780 127700 605070
rect 127740 604780 127760 605070
rect 127680 604760 127760 604780
rect 127800 605070 127860 605090
rect 127800 604780 127810 605070
rect 127850 604780 127860 605070
rect 127800 604710 127860 604780
rect 127920 605070 127980 605090
rect 127920 604780 127930 605070
rect 127970 604780 127980 605070
rect 127920 604710 127980 604780
rect 128020 605070 128100 605090
rect 128020 604780 128040 605070
rect 128080 604780 128100 605070
rect 128020 604760 128100 604780
rect 128140 605070 128200 605090
rect 128140 604780 128150 605070
rect 128190 604780 128200 605070
rect 128140 604710 128200 604780
rect 128260 605070 128320 605090
rect 128260 604780 128270 605070
rect 128310 604780 128320 605070
rect 128260 604710 128320 604780
rect 128360 605070 128440 605090
rect 128360 604780 128380 605070
rect 128420 604780 128440 605070
rect 128360 604760 128440 604780
rect 128480 605070 128540 605090
rect 128480 604780 128490 605070
rect 128530 604780 128540 605070
rect 128480 604710 128540 604780
rect 128600 605070 128660 605090
rect 128600 604780 128610 605070
rect 128650 604780 128660 605070
rect 128600 604710 128660 604780
rect 128700 605070 128780 605090
rect 128700 604780 128720 605070
rect 128760 604780 128780 605070
rect 128700 604760 128780 604780
rect 128820 605070 128880 605090
rect 128820 604780 128830 605070
rect 128870 604780 128880 605070
rect 128820 604710 128880 604780
rect 128940 605070 129000 605090
rect 128940 604780 128950 605070
rect 128990 604780 129000 605070
rect 128940 604710 129000 604780
rect 129040 605070 129120 605090
rect 129040 604780 129060 605070
rect 129100 604780 129120 605070
rect 129040 604760 129120 604780
rect 129160 605070 129220 605090
rect 129160 604780 129170 605070
rect 129210 604780 129220 605070
rect 129160 604710 129220 604780
rect 129280 605070 129340 605090
rect 129280 604780 129290 605070
rect 129330 604780 129340 605070
rect 129280 604710 129340 604780
rect 129380 605070 129460 605090
rect 129380 604780 129400 605070
rect 129440 604780 129460 605070
rect 129380 604760 129460 604780
rect 129500 605070 129560 605090
rect 129500 604780 129510 605070
rect 129550 604780 129560 605070
rect 129500 604710 129560 604780
rect 129620 605070 129680 605090
rect 129620 604780 129630 605070
rect 129670 604780 129680 605070
rect 129620 604710 129680 604780
rect 129720 605070 129800 605090
rect 129720 604780 129740 605070
rect 129780 604780 129800 605070
rect 129720 604760 129800 604780
rect 129840 605070 129900 605090
rect 129840 604780 129850 605070
rect 129890 604780 129900 605070
rect 129840 604710 129900 604780
rect 129960 605070 130020 605090
rect 129960 604780 129970 605070
rect 130010 604780 130020 605070
rect 129960 604710 130020 604780
rect 130060 605070 130140 605090
rect 130060 604780 130080 605070
rect 130120 604780 130140 605070
rect 130060 604760 130140 604780
rect 130180 605070 130240 605090
rect 130180 604780 130190 605070
rect 130230 604780 130240 605070
rect 130180 604710 130240 604780
rect 130300 605070 130360 605090
rect 130300 604780 130310 605070
rect 130350 604780 130360 605070
rect 130300 604710 130360 604780
rect 130400 605070 130480 605090
rect 130400 604780 130420 605070
rect 130460 604780 130480 605070
rect 130400 604760 130480 604780
rect 130520 605070 130580 605090
rect 130520 604780 130530 605070
rect 130570 604780 130580 605070
rect 130520 604710 130580 604780
rect 130640 605070 130700 605090
rect 130640 604780 130650 605070
rect 130690 604780 130700 605070
rect 130640 604710 130700 604780
rect 130740 605070 130820 605090
rect 130740 604780 130760 605070
rect 130800 604780 130820 605070
rect 130740 604760 130820 604780
rect 130860 605070 130920 605090
rect 130860 604780 130870 605070
rect 130910 604780 130920 605070
rect 130860 604710 130920 604780
rect 130980 605070 131040 605090
rect 130980 604780 130990 605070
rect 131030 604780 131040 605070
rect 130980 604710 131040 604780
rect 131080 605070 131160 605090
rect 131080 604780 131100 605070
rect 131140 604780 131160 605070
rect 131080 604760 131160 604780
rect 131200 605070 131260 605090
rect 131200 604780 131210 605070
rect 131250 604780 131260 605070
rect 131200 604710 131260 604780
rect 131320 605070 131380 605090
rect 131320 604780 131330 605070
rect 131370 604780 131380 605070
rect 131320 604710 131380 604780
rect 131420 605070 131500 605090
rect 131420 604780 131440 605070
rect 131480 604780 131500 605070
rect 131420 604760 131500 604780
rect 131540 605070 131600 605090
rect 131540 604780 131550 605070
rect 131590 604780 131600 605070
rect 131540 604710 131600 604780
rect 125200 604650 128160 604710
rect 128640 604650 131600 604710
rect 131690 604640 131720 605310
rect 131850 604640 131880 605310
rect 131690 604620 131880 604640
rect 119290 601766 119390 601772
rect 119290 601686 119296 601766
rect 119388 601686 119390 601766
rect 119136 601306 119236 601314
rect 119136 601222 119144 601306
rect 119226 601222 119236 601306
rect 119136 601208 119236 601222
rect 119290 601104 119390 601686
rect 119450 601190 120048 601210
rect 119450 601184 120052 601190
rect 119450 601110 119958 601184
rect 119952 601104 119958 601110
rect 120050 601104 120052 601184
rect 119952 601066 120052 601104
rect 120618 600340 123930 600440
rect 123822 599880 123922 600340
rect 123816 599780 123922 599880
rect 123822 599070 123922 599780
rect 124880 599640 125300 599700
rect 125040 599610 125100 599640
rect 124930 599590 124990 599610
rect 124930 599550 124940 599590
rect 124980 599550 124990 599590
rect 124930 599420 124990 599550
rect 125030 599590 125110 599610
rect 125030 599550 125050 599590
rect 125090 599550 125110 599590
rect 125030 599530 125110 599550
rect 125150 599590 125210 599610
rect 125150 599550 125160 599590
rect 125200 599550 125210 599590
rect 125150 599420 125210 599550
rect 125170 599070 131348 599074
rect 123820 599010 131348 599070
rect 123820 598970 125170 599010
rect 125210 598974 125510 599010
rect 125210 598970 125220 598974
rect 125160 598950 125220 598970
rect 125500 598970 125510 598974
rect 125550 598974 125850 599010
rect 125550 598970 125560 598974
rect 125500 598950 125560 598970
rect 125840 598970 125850 598974
rect 125890 598974 126190 599010
rect 125890 598970 125900 598974
rect 125840 598950 125900 598970
rect 126180 598970 126190 598974
rect 126230 598974 126530 599010
rect 126230 598970 126240 598974
rect 126180 598950 126240 598970
rect 126520 598970 126530 598974
rect 126570 598974 126870 599010
rect 126570 598970 126580 598974
rect 126520 598950 126580 598970
rect 126860 598970 126870 598974
rect 126910 598974 127210 599010
rect 126910 598970 126920 598974
rect 126860 598950 126920 598970
rect 127200 598970 127210 598974
rect 127250 598974 127550 599010
rect 127250 598970 127260 598974
rect 127200 598950 127260 598970
rect 127540 598970 127550 598974
rect 127590 598974 127890 599010
rect 127590 598970 127600 598974
rect 127540 598950 127600 598970
rect 127880 598970 127890 598974
rect 127930 598974 128230 599010
rect 127930 598970 127940 598974
rect 127880 598950 127940 598970
rect 128220 598970 128230 598974
rect 128270 598974 128570 599010
rect 128270 598970 128280 598974
rect 128220 598950 128280 598970
rect 128560 598970 128570 598974
rect 128610 598974 128910 599010
rect 128610 598970 128620 598974
rect 128560 598950 128620 598970
rect 128900 598970 128910 598974
rect 128950 598974 129250 599010
rect 128950 598970 128960 598974
rect 128900 598950 128960 598970
rect 129240 598970 129250 598974
rect 129290 598974 129590 599010
rect 129290 598970 129300 598974
rect 129240 598950 129300 598970
rect 129580 598970 129590 598974
rect 129630 598974 129930 599010
rect 129630 598970 129640 598974
rect 129580 598950 129640 598970
rect 129920 598970 129930 598974
rect 129970 598974 130270 599010
rect 129970 598970 129980 598974
rect 129920 598950 129980 598970
rect 130260 598970 130270 598974
rect 130310 598974 130610 599010
rect 130310 598970 130320 598974
rect 130260 598950 130320 598970
rect 130600 598970 130610 598974
rect 130650 598974 130950 599010
rect 130650 598970 130660 598974
rect 130600 598950 130660 598970
rect 130940 598970 130950 598974
rect 130990 598974 131290 599010
rect 130990 598970 131000 598974
rect 130940 598950 131000 598970
rect 131280 598970 131290 598974
rect 131330 598974 131348 599010
rect 131490 599050 131680 599070
rect 131330 598970 131340 598974
rect 131280 598950 131340 598970
rect 124940 598860 127960 598920
rect 128440 598860 131400 598920
rect 125110 598830 125170 598860
rect 125450 598830 125510 598860
rect 125790 598830 125850 598860
rect 126130 598830 126190 598860
rect 126470 598830 126530 598860
rect 126810 598830 126870 598860
rect 127150 598830 127210 598860
rect 127490 598830 127550 598860
rect 127830 598830 127890 598860
rect 128170 598830 128230 598860
rect 128510 598830 128570 598860
rect 128850 598830 128910 598860
rect 129190 598830 129250 598860
rect 129530 598830 129590 598860
rect 129870 598830 129930 598860
rect 130210 598830 130270 598860
rect 130550 598830 130610 598860
rect 130890 598830 130950 598860
rect 131230 598830 131290 598860
rect 125000 598810 125060 598830
rect 125000 598420 125010 598810
rect 125050 598420 125060 598810
rect 125000 598350 125060 598420
rect 125100 598810 125180 598830
rect 125100 598420 125120 598810
rect 125160 598420 125180 598810
rect 125100 598400 125180 598420
rect 125220 598810 125280 598830
rect 125220 598420 125230 598810
rect 125270 598420 125280 598810
rect 125220 598350 125280 598420
rect 125340 598810 125400 598830
rect 125340 598420 125350 598810
rect 125390 598420 125400 598810
rect 125340 598350 125400 598420
rect 125440 598810 125520 598830
rect 125440 598420 125460 598810
rect 125500 598420 125520 598810
rect 125440 598400 125520 598420
rect 125560 598810 125620 598830
rect 125560 598420 125570 598810
rect 125610 598420 125620 598810
rect 125560 598350 125620 598420
rect 125680 598810 125740 598830
rect 125680 598420 125690 598810
rect 125730 598420 125740 598810
rect 125680 598350 125740 598420
rect 125780 598810 125860 598830
rect 125780 598420 125800 598810
rect 125840 598420 125860 598810
rect 125780 598400 125860 598420
rect 125900 598810 125960 598830
rect 125900 598420 125910 598810
rect 125950 598420 125960 598810
rect 125900 598350 125960 598420
rect 126020 598810 126080 598830
rect 126020 598420 126030 598810
rect 126070 598420 126080 598810
rect 126020 598350 126080 598420
rect 126120 598810 126200 598830
rect 126120 598420 126140 598810
rect 126180 598420 126200 598810
rect 126120 598400 126200 598420
rect 126240 598810 126300 598830
rect 126240 598420 126250 598810
rect 126290 598420 126300 598810
rect 126240 598350 126300 598420
rect 126360 598810 126420 598830
rect 126360 598420 126370 598810
rect 126410 598420 126420 598810
rect 126360 598350 126420 598420
rect 126460 598810 126540 598830
rect 126460 598420 126480 598810
rect 126520 598420 126540 598810
rect 126460 598400 126540 598420
rect 126580 598810 126640 598830
rect 126580 598420 126590 598810
rect 126630 598420 126640 598810
rect 126580 598350 126640 598420
rect 126700 598810 126760 598830
rect 126700 598420 126710 598810
rect 126750 598420 126760 598810
rect 126700 598350 126760 598420
rect 126800 598810 126880 598830
rect 126800 598420 126820 598810
rect 126860 598420 126880 598810
rect 126800 598400 126880 598420
rect 126920 598810 126980 598830
rect 126920 598420 126930 598810
rect 126970 598420 126980 598810
rect 126920 598350 126980 598420
rect 127040 598810 127100 598830
rect 127040 598420 127050 598810
rect 127090 598420 127100 598810
rect 127040 598350 127100 598420
rect 127140 598810 127220 598830
rect 127140 598420 127160 598810
rect 127200 598420 127220 598810
rect 127140 598400 127220 598420
rect 127260 598810 127320 598830
rect 127260 598420 127270 598810
rect 127310 598420 127320 598810
rect 127260 598350 127320 598420
rect 127380 598810 127440 598830
rect 127380 598420 127390 598810
rect 127430 598420 127440 598810
rect 127380 598350 127440 598420
rect 127480 598810 127560 598830
rect 127480 598420 127500 598810
rect 127540 598420 127560 598810
rect 127480 598400 127560 598420
rect 127600 598810 127660 598830
rect 127600 598420 127610 598810
rect 127650 598420 127660 598810
rect 127600 598350 127660 598420
rect 127720 598810 127780 598830
rect 127720 598420 127730 598810
rect 127770 598420 127780 598810
rect 127720 598350 127780 598420
rect 127820 598810 127900 598830
rect 127820 598420 127840 598810
rect 127880 598420 127900 598810
rect 127820 598400 127900 598420
rect 127940 598810 128000 598830
rect 127940 598420 127950 598810
rect 127990 598420 128000 598810
rect 127940 598350 128000 598420
rect 128060 598810 128120 598830
rect 128060 598420 128070 598810
rect 128110 598420 128120 598810
rect 128060 598350 128120 598420
rect 128160 598810 128240 598830
rect 128160 598420 128180 598810
rect 128220 598420 128240 598810
rect 128160 598400 128240 598420
rect 128280 598810 128340 598830
rect 128280 598420 128290 598810
rect 128330 598420 128340 598810
rect 128280 598350 128340 598420
rect 128400 598810 128460 598830
rect 128400 598420 128410 598810
rect 128450 598420 128460 598810
rect 128400 598350 128460 598420
rect 128500 598810 128580 598830
rect 128500 598420 128520 598810
rect 128560 598420 128580 598810
rect 128500 598400 128580 598420
rect 128620 598810 128680 598830
rect 128620 598420 128630 598810
rect 128670 598420 128680 598810
rect 128620 598350 128680 598420
rect 128740 598810 128800 598830
rect 128740 598420 128750 598810
rect 128790 598420 128800 598810
rect 128740 598350 128800 598420
rect 128840 598810 128920 598830
rect 128840 598420 128860 598810
rect 128900 598420 128920 598810
rect 128840 598400 128920 598420
rect 128960 598810 129020 598830
rect 128960 598420 128970 598810
rect 129010 598420 129020 598810
rect 128960 598350 129020 598420
rect 129080 598810 129140 598830
rect 129080 598420 129090 598810
rect 129130 598420 129140 598810
rect 129080 598350 129140 598420
rect 129180 598810 129260 598830
rect 129180 598420 129200 598810
rect 129240 598420 129260 598810
rect 129180 598400 129260 598420
rect 129300 598810 129360 598830
rect 129300 598420 129310 598810
rect 129350 598420 129360 598810
rect 129300 598350 129360 598420
rect 129420 598810 129480 598830
rect 129420 598420 129430 598810
rect 129470 598420 129480 598810
rect 129420 598350 129480 598420
rect 129520 598810 129600 598830
rect 129520 598420 129540 598810
rect 129580 598420 129600 598810
rect 129520 598400 129600 598420
rect 129640 598810 129700 598830
rect 129640 598420 129650 598810
rect 129690 598420 129700 598810
rect 129640 598350 129700 598420
rect 129760 598810 129820 598830
rect 129760 598420 129770 598810
rect 129810 598420 129820 598810
rect 129760 598350 129820 598420
rect 129860 598810 129940 598830
rect 129860 598420 129880 598810
rect 129920 598420 129940 598810
rect 129860 598400 129940 598420
rect 129980 598810 130040 598830
rect 129980 598420 129990 598810
rect 130030 598420 130040 598810
rect 129980 598350 130040 598420
rect 130100 598810 130160 598830
rect 130100 598420 130110 598810
rect 130150 598420 130160 598810
rect 130100 598350 130160 598420
rect 130200 598810 130280 598830
rect 130200 598420 130220 598810
rect 130260 598420 130280 598810
rect 130200 598400 130280 598420
rect 130320 598810 130380 598830
rect 130320 598420 130330 598810
rect 130370 598420 130380 598810
rect 130320 598350 130380 598420
rect 130440 598810 130500 598830
rect 130440 598420 130450 598810
rect 130490 598420 130500 598810
rect 130440 598350 130500 598420
rect 130540 598810 130620 598830
rect 130540 598420 130560 598810
rect 130600 598420 130620 598810
rect 130540 598400 130620 598420
rect 130660 598810 130720 598830
rect 130660 598420 130670 598810
rect 130710 598420 130720 598810
rect 130660 598350 130720 598420
rect 130780 598810 130840 598830
rect 130780 598420 130790 598810
rect 130830 598420 130840 598810
rect 130780 598350 130840 598420
rect 130880 598810 130960 598830
rect 130880 598420 130900 598810
rect 130940 598420 130960 598810
rect 130880 598400 130960 598420
rect 131000 598810 131060 598830
rect 131000 598420 131010 598810
rect 131050 598420 131060 598810
rect 131000 598350 131060 598420
rect 131120 598810 131180 598830
rect 131120 598420 131130 598810
rect 131170 598420 131180 598810
rect 131120 598350 131180 598420
rect 131220 598810 131300 598830
rect 131220 598420 131240 598810
rect 131280 598420 131300 598810
rect 131220 598400 131300 598420
rect 131340 598810 131400 598830
rect 131340 598420 131350 598810
rect 131390 598420 131400 598810
rect 131340 598350 131400 598420
rect 125000 598290 127960 598350
rect 128440 598290 131400 598350
rect 131490 598280 131520 599050
rect 131650 598280 131680 599050
rect 131490 598260 131680 598280
rect 119250 594240 119350 594244
rect 119250 594234 119430 594240
rect 119250 594154 119336 594234
rect 119428 594154 119430 594234
rect 119250 594116 119430 594154
rect 119096 593756 119196 593764
rect 119096 593672 119104 593756
rect 119186 593672 119196 593756
rect 119096 593660 119196 593672
rect 119090 593658 119196 593660
rect 119090 593430 119190 593658
rect 119090 593370 119110 593430
rect 119170 593370 119190 593430
rect 119090 593350 119190 593370
rect 119250 592950 119350 594116
rect 119410 593632 120018 593660
rect 119410 593626 120020 593632
rect 119410 593560 119926 593626
rect 119410 593540 119510 593560
rect 119410 593480 119430 593540
rect 119490 593480 119510 593540
rect 119920 593546 119926 593560
rect 120018 593546 120020 593626
rect 119920 593508 120020 593546
rect 119410 593460 119510 593480
rect 119840 593040 119940 593060
rect 120210 593040 120310 593050
rect 119840 592980 119860 593040
rect 119920 593030 120310 593040
rect 119920 592980 120230 593030
rect 119840 592960 119940 592980
rect 120210 592970 120230 592980
rect 120290 592970 120310 593030
rect 120210 592950 120310 592970
rect 119250 592900 119270 592950
rect 119310 592900 119350 592950
rect 119250 592520 119350 592900
rect 119600 592880 119700 592890
rect 119600 592800 119610 592880
rect 119690 592800 119700 592880
rect 119600 592790 119700 592800
rect 119840 592870 123878 592890
rect 119840 592810 119860 592870
rect 119920 592854 123878 592870
rect 119920 592810 123882 592854
rect 119840 592790 123882 592810
rect 119250 592460 119270 592520
rect 119330 592460 119350 592520
rect 119250 592450 119350 592460
rect 123782 592330 123882 592790
rect 123774 592230 123882 592330
rect 123782 591520 123882 592230
rect 124840 592090 125260 592150
rect 125000 592060 125060 592090
rect 124890 592040 124950 592060
rect 124890 592000 124900 592040
rect 124940 592000 124950 592040
rect 124890 591870 124950 592000
rect 124990 592040 125070 592060
rect 124990 592000 125010 592040
rect 125050 592000 125070 592040
rect 124990 591980 125070 592000
rect 125110 592040 125170 592060
rect 125110 592000 125120 592040
rect 125160 592000 125170 592040
rect 125110 591870 125170 592000
rect 125130 591520 131308 591524
rect 123780 591460 131308 591520
rect 123780 591420 125130 591460
rect 125170 591424 125470 591460
rect 125170 591420 125180 591424
rect 125120 591400 125180 591420
rect 125460 591420 125470 591424
rect 125510 591424 125810 591460
rect 125510 591420 125520 591424
rect 125460 591400 125520 591420
rect 125800 591420 125810 591424
rect 125850 591424 126150 591460
rect 125850 591420 125860 591424
rect 125800 591400 125860 591420
rect 126140 591420 126150 591424
rect 126190 591424 126490 591460
rect 126190 591420 126200 591424
rect 126140 591400 126200 591420
rect 126480 591420 126490 591424
rect 126530 591424 126830 591460
rect 126530 591420 126540 591424
rect 126480 591400 126540 591420
rect 126820 591420 126830 591424
rect 126870 591424 127170 591460
rect 126870 591420 126880 591424
rect 126820 591400 126880 591420
rect 127160 591420 127170 591424
rect 127210 591424 127510 591460
rect 127210 591420 127220 591424
rect 127160 591400 127220 591420
rect 127500 591420 127510 591424
rect 127550 591424 127850 591460
rect 127550 591420 127560 591424
rect 127500 591400 127560 591420
rect 127840 591420 127850 591424
rect 127890 591424 128190 591460
rect 127890 591420 127900 591424
rect 127840 591400 127900 591420
rect 128180 591420 128190 591424
rect 128230 591424 128530 591460
rect 128230 591420 128240 591424
rect 128180 591400 128240 591420
rect 128520 591420 128530 591424
rect 128570 591424 128870 591460
rect 128570 591420 128580 591424
rect 128520 591400 128580 591420
rect 128860 591420 128870 591424
rect 128910 591424 129210 591460
rect 128910 591420 128920 591424
rect 128860 591400 128920 591420
rect 129200 591420 129210 591424
rect 129250 591424 129550 591460
rect 129250 591420 129260 591424
rect 129200 591400 129260 591420
rect 129540 591420 129550 591424
rect 129590 591424 129890 591460
rect 129590 591420 129600 591424
rect 129540 591400 129600 591420
rect 129880 591420 129890 591424
rect 129930 591424 130230 591460
rect 129930 591420 129940 591424
rect 129880 591400 129940 591420
rect 130220 591420 130230 591424
rect 130270 591424 130570 591460
rect 130270 591420 130280 591424
rect 130220 591400 130280 591420
rect 130560 591420 130570 591424
rect 130610 591424 130910 591460
rect 130610 591420 130620 591424
rect 130560 591400 130620 591420
rect 130900 591420 130910 591424
rect 130950 591424 131250 591460
rect 130950 591420 130960 591424
rect 130900 591400 130960 591420
rect 131240 591420 131250 591424
rect 131290 591424 131308 591460
rect 131450 591500 131640 591520
rect 131290 591420 131300 591424
rect 131240 591400 131300 591420
rect 124900 591310 127920 591370
rect 128400 591310 131360 591370
rect 125070 591280 125130 591310
rect 125410 591280 125470 591310
rect 125750 591280 125810 591310
rect 126090 591280 126150 591310
rect 126430 591280 126490 591310
rect 126770 591280 126830 591310
rect 127110 591280 127170 591310
rect 127450 591280 127510 591310
rect 127790 591280 127850 591310
rect 128130 591280 128190 591310
rect 128470 591280 128530 591310
rect 128810 591280 128870 591310
rect 129150 591280 129210 591310
rect 129490 591280 129550 591310
rect 129830 591280 129890 591310
rect 130170 591280 130230 591310
rect 130510 591280 130570 591310
rect 130850 591280 130910 591310
rect 131190 591280 131250 591310
rect 124960 591260 125020 591280
rect 124960 590770 124970 591260
rect 125010 590770 125020 591260
rect 124960 590700 125020 590770
rect 125060 591260 125140 591280
rect 125060 590770 125080 591260
rect 125120 590770 125140 591260
rect 125060 590750 125140 590770
rect 125180 591260 125240 591280
rect 125180 590770 125190 591260
rect 125230 590770 125240 591260
rect 125180 590700 125240 590770
rect 125300 591260 125360 591280
rect 125300 590770 125310 591260
rect 125350 590770 125360 591260
rect 125300 590700 125360 590770
rect 125400 591260 125480 591280
rect 125400 590770 125420 591260
rect 125460 590770 125480 591260
rect 125400 590750 125480 590770
rect 125520 591260 125580 591280
rect 125520 590770 125530 591260
rect 125570 590770 125580 591260
rect 125520 590700 125580 590770
rect 125640 591260 125700 591280
rect 125640 590770 125650 591260
rect 125690 590770 125700 591260
rect 125640 590700 125700 590770
rect 125740 591260 125820 591280
rect 125740 590770 125760 591260
rect 125800 590770 125820 591260
rect 125740 590750 125820 590770
rect 125860 591260 125920 591280
rect 125860 590770 125870 591260
rect 125910 590770 125920 591260
rect 125860 590700 125920 590770
rect 125980 591260 126040 591280
rect 125980 590770 125990 591260
rect 126030 590770 126040 591260
rect 125980 590700 126040 590770
rect 126080 591260 126160 591280
rect 126080 590770 126100 591260
rect 126140 590770 126160 591260
rect 126080 590750 126160 590770
rect 126200 591260 126260 591280
rect 126200 590770 126210 591260
rect 126250 590770 126260 591260
rect 126200 590700 126260 590770
rect 126320 591260 126380 591280
rect 126320 590770 126330 591260
rect 126370 590770 126380 591260
rect 126320 590700 126380 590770
rect 126420 591260 126500 591280
rect 126420 590770 126440 591260
rect 126480 590770 126500 591260
rect 126420 590750 126500 590770
rect 126540 591260 126600 591280
rect 126540 590770 126550 591260
rect 126590 590770 126600 591260
rect 126540 590700 126600 590770
rect 126660 591260 126720 591280
rect 126660 590770 126670 591260
rect 126710 590770 126720 591260
rect 126660 590700 126720 590770
rect 126760 591260 126840 591280
rect 126760 590770 126780 591260
rect 126820 590770 126840 591260
rect 126760 590750 126840 590770
rect 126880 591260 126940 591280
rect 126880 590770 126890 591260
rect 126930 590770 126940 591260
rect 126880 590700 126940 590770
rect 127000 591260 127060 591280
rect 127000 590770 127010 591260
rect 127050 590770 127060 591260
rect 127000 590700 127060 590770
rect 127100 591260 127180 591280
rect 127100 590770 127120 591260
rect 127160 590770 127180 591260
rect 127100 590750 127180 590770
rect 127220 591260 127280 591280
rect 127220 590770 127230 591260
rect 127270 590770 127280 591260
rect 127220 590700 127280 590770
rect 127340 591260 127400 591280
rect 127340 590770 127350 591260
rect 127390 590770 127400 591260
rect 127340 590700 127400 590770
rect 127440 591260 127520 591280
rect 127440 590770 127460 591260
rect 127500 590770 127520 591260
rect 127440 590750 127520 590770
rect 127560 591260 127620 591280
rect 127560 590770 127570 591260
rect 127610 590770 127620 591260
rect 127560 590700 127620 590770
rect 127680 591260 127740 591280
rect 127680 590770 127690 591260
rect 127730 590770 127740 591260
rect 127680 590700 127740 590770
rect 127780 591260 127860 591280
rect 127780 590770 127800 591260
rect 127840 590770 127860 591260
rect 127780 590750 127860 590770
rect 127900 591260 127960 591280
rect 127900 590770 127910 591260
rect 127950 590770 127960 591260
rect 127900 590700 127960 590770
rect 128020 591260 128080 591280
rect 128020 590770 128030 591260
rect 128070 590770 128080 591260
rect 128020 590700 128080 590770
rect 128120 591260 128200 591280
rect 128120 590770 128140 591260
rect 128180 590770 128200 591260
rect 128120 590750 128200 590770
rect 128240 591260 128300 591280
rect 128240 590770 128250 591260
rect 128290 590770 128300 591260
rect 128240 590700 128300 590770
rect 128360 591260 128420 591280
rect 128360 590770 128370 591260
rect 128410 590770 128420 591260
rect 128360 590700 128420 590770
rect 128460 591260 128540 591280
rect 128460 590770 128480 591260
rect 128520 590770 128540 591260
rect 128460 590750 128540 590770
rect 128580 591260 128640 591280
rect 128580 590770 128590 591260
rect 128630 590770 128640 591260
rect 128580 590700 128640 590770
rect 128700 591260 128760 591280
rect 128700 590770 128710 591260
rect 128750 590770 128760 591260
rect 128700 590700 128760 590770
rect 128800 591260 128880 591280
rect 128800 590770 128820 591260
rect 128860 590770 128880 591260
rect 128800 590750 128880 590770
rect 128920 591260 128980 591280
rect 128920 590770 128930 591260
rect 128970 590770 128980 591260
rect 128920 590700 128980 590770
rect 129040 591260 129100 591280
rect 129040 590770 129050 591260
rect 129090 590770 129100 591260
rect 129040 590700 129100 590770
rect 129140 591260 129220 591280
rect 129140 590770 129160 591260
rect 129200 590770 129220 591260
rect 129140 590750 129220 590770
rect 129260 591260 129320 591280
rect 129260 590770 129270 591260
rect 129310 590770 129320 591260
rect 129260 590700 129320 590770
rect 129380 591260 129440 591280
rect 129380 590770 129390 591260
rect 129430 590770 129440 591260
rect 129380 590700 129440 590770
rect 129480 591260 129560 591280
rect 129480 590770 129500 591260
rect 129540 590770 129560 591260
rect 129480 590750 129560 590770
rect 129600 591260 129660 591280
rect 129600 590770 129610 591260
rect 129650 590770 129660 591260
rect 129600 590700 129660 590770
rect 129720 591260 129780 591280
rect 129720 590770 129730 591260
rect 129770 590770 129780 591260
rect 129720 590700 129780 590770
rect 129820 591260 129900 591280
rect 129820 590770 129840 591260
rect 129880 590770 129900 591260
rect 129820 590750 129900 590770
rect 129940 591260 130000 591280
rect 129940 590770 129950 591260
rect 129990 590770 130000 591260
rect 129940 590700 130000 590770
rect 130060 591260 130120 591280
rect 130060 590770 130070 591260
rect 130110 590770 130120 591260
rect 130060 590700 130120 590770
rect 130160 591260 130240 591280
rect 130160 590770 130180 591260
rect 130220 590770 130240 591260
rect 130160 590750 130240 590770
rect 130280 591260 130340 591280
rect 130280 590770 130290 591260
rect 130330 590770 130340 591260
rect 130280 590700 130340 590770
rect 130400 591260 130460 591280
rect 130400 590770 130410 591260
rect 130450 590770 130460 591260
rect 130400 590700 130460 590770
rect 130500 591260 130580 591280
rect 130500 590770 130520 591260
rect 130560 590770 130580 591260
rect 130500 590750 130580 590770
rect 130620 591260 130680 591280
rect 130620 590770 130630 591260
rect 130670 590770 130680 591260
rect 130620 590700 130680 590770
rect 130740 591260 130800 591280
rect 130740 590770 130750 591260
rect 130790 590770 130800 591260
rect 130740 590700 130800 590770
rect 130840 591260 130920 591280
rect 130840 590770 130860 591260
rect 130900 590770 130920 591260
rect 130840 590750 130920 590770
rect 130960 591260 131020 591280
rect 130960 590770 130970 591260
rect 131010 590770 131020 591260
rect 130960 590700 131020 590770
rect 131080 591260 131140 591280
rect 131080 590770 131090 591260
rect 131130 590770 131140 591260
rect 131080 590700 131140 590770
rect 131180 591260 131260 591280
rect 131180 590770 131200 591260
rect 131240 590770 131260 591260
rect 131180 590750 131260 590770
rect 131300 591260 131360 591280
rect 131300 590770 131310 591260
rect 131350 590770 131360 591260
rect 131300 590700 131360 590770
rect 124960 590640 127920 590700
rect 128400 590640 131360 590700
rect 131450 590630 131480 591500
rect 131610 590630 131640 591500
rect 131450 590610 131640 590630
rect 119300 584682 119400 584688
rect 119300 584668 119306 584682
rect 119290 584602 119306 584668
rect 119398 584602 119400 584682
rect 119290 584564 119400 584602
rect 119136 584214 119236 584222
rect 119136 584130 119144 584214
rect 119226 584130 119236 584214
rect 119136 584120 119236 584130
rect 119130 584116 119236 584120
rect 119130 583890 119230 584116
rect 119130 583830 119150 583890
rect 119210 583830 119230 583890
rect 119130 583810 119230 583830
rect 119290 583410 119390 584564
rect 119450 584114 120216 584120
rect 119450 584108 120222 584114
rect 119450 584028 120128 584108
rect 120220 584028 120222 584108
rect 119450 584020 120222 584028
rect 119450 584000 119550 584020
rect 119450 583940 119470 584000
rect 119530 583940 119550 584000
rect 120122 583990 120222 584020
rect 119450 583920 119550 583940
rect 119880 583500 119980 583520
rect 120250 583500 120350 583510
rect 119880 583440 119900 583500
rect 119960 583490 120350 583500
rect 119960 583440 120270 583490
rect 119880 583420 119980 583440
rect 120250 583430 120270 583440
rect 120330 583430 120350 583490
rect 120250 583410 120350 583430
rect 119290 583360 119310 583410
rect 119350 583360 119390 583410
rect 119290 582980 119390 583360
rect 119640 583340 119740 583350
rect 119640 583260 119650 583340
rect 119730 583260 119740 583340
rect 119640 583250 119740 583260
rect 119880 583330 124342 583350
rect 119880 583270 119900 583330
rect 119960 583270 124342 583330
rect 119880 583250 124342 583270
rect 119290 582920 119310 582980
rect 119370 582920 119390 582980
rect 119290 582910 119390 582920
rect 124242 582544 124342 583250
rect 125300 583110 125720 583170
rect 125460 583080 125520 583110
rect 125350 583060 125410 583080
rect 125350 583020 125360 583060
rect 125400 583020 125410 583060
rect 125350 582890 125410 583020
rect 125450 583060 125530 583080
rect 125450 583020 125470 583060
rect 125510 583020 125530 583060
rect 125450 583000 125530 583020
rect 125570 583060 125630 583080
rect 125570 583020 125580 583060
rect 125620 583020 125630 583060
rect 125570 582890 125630 583020
rect 124242 582480 132718 582544
rect 124242 582444 125640 582480
rect 125630 582440 125640 582444
rect 125680 582444 126030 582480
rect 125680 582440 125690 582444
rect 125630 582420 125690 582440
rect 126020 582440 126030 582444
rect 126070 582444 126420 582480
rect 126070 582440 126080 582444
rect 126020 582420 126080 582440
rect 126410 582440 126420 582444
rect 126460 582444 126810 582480
rect 126460 582440 126470 582444
rect 126410 582420 126470 582440
rect 126800 582440 126810 582444
rect 126850 582444 127200 582480
rect 126850 582440 126860 582444
rect 126800 582420 126860 582440
rect 127190 582440 127200 582444
rect 127240 582444 127590 582480
rect 127240 582440 127250 582444
rect 127190 582420 127250 582440
rect 127580 582440 127590 582444
rect 127630 582444 127980 582480
rect 127630 582440 127640 582444
rect 127580 582420 127640 582440
rect 127970 582440 127980 582444
rect 128020 582444 128370 582480
rect 128020 582440 128030 582444
rect 127970 582420 128030 582440
rect 128360 582440 128370 582444
rect 128410 582444 128760 582480
rect 128410 582440 128420 582444
rect 128360 582420 128420 582440
rect 128750 582440 128760 582444
rect 128800 582444 129150 582480
rect 128800 582440 128810 582444
rect 128750 582420 128810 582440
rect 129140 582440 129150 582444
rect 129190 582444 129540 582480
rect 129190 582440 129200 582444
rect 129140 582420 129200 582440
rect 129530 582440 129540 582444
rect 129580 582444 129930 582480
rect 129580 582440 129590 582444
rect 129530 582420 129590 582440
rect 129920 582440 129930 582444
rect 129970 582444 130320 582480
rect 129970 582440 129980 582444
rect 129920 582420 129980 582440
rect 130310 582440 130320 582444
rect 130360 582444 130710 582480
rect 130360 582440 130370 582444
rect 130310 582420 130370 582440
rect 130700 582440 130710 582444
rect 130750 582444 131100 582480
rect 130750 582440 130760 582444
rect 130700 582420 130760 582440
rect 131090 582440 131100 582444
rect 131140 582444 131490 582480
rect 131140 582440 131150 582444
rect 131090 582420 131150 582440
rect 131480 582440 131490 582444
rect 131530 582444 131880 582480
rect 131530 582440 131540 582444
rect 131480 582420 131540 582440
rect 131870 582440 131880 582444
rect 131920 582444 132270 582480
rect 131920 582440 131930 582444
rect 131870 582420 131930 582440
rect 132260 582440 132270 582444
rect 132310 582444 132660 582480
rect 132310 582440 132320 582444
rect 132260 582420 132320 582440
rect 132650 582440 132660 582444
rect 132700 582444 132718 582480
rect 132860 582520 133050 582540
rect 132700 582440 132710 582444
rect 132650 582420 132710 582440
rect 125360 582330 128370 582390
rect 128870 582330 132770 582390
rect 125530 582300 125640 582330
rect 125920 582300 126030 582330
rect 126310 582300 126420 582330
rect 126700 582300 126810 582330
rect 127090 582300 127200 582330
rect 127480 582300 127590 582330
rect 127870 582300 127980 582330
rect 128260 582300 128370 582330
rect 128650 582300 128760 582330
rect 129040 582300 129150 582330
rect 129430 582300 129540 582330
rect 129820 582300 129930 582330
rect 130210 582300 130320 582330
rect 130600 582300 130710 582330
rect 130990 582300 131100 582330
rect 131380 582300 131490 582330
rect 131770 582300 131880 582330
rect 132160 582300 132270 582330
rect 132550 582300 132660 582330
rect 125420 582280 125480 582300
rect 125420 582240 125430 582280
rect 125470 582240 125480 582280
rect 125420 582170 125480 582240
rect 125520 582280 125650 582300
rect 125520 582240 125540 582280
rect 125630 582240 125650 582280
rect 125520 582220 125650 582240
rect 125690 582280 125750 582300
rect 125690 582240 125700 582280
rect 125740 582240 125750 582280
rect 125690 582170 125750 582240
rect 125810 582280 125870 582300
rect 125810 582240 125820 582280
rect 125860 582240 125870 582280
rect 125810 582170 125870 582240
rect 125910 582280 126040 582300
rect 125910 582240 125930 582280
rect 126020 582240 126040 582280
rect 125910 582220 126040 582240
rect 126080 582280 126140 582300
rect 126080 582240 126090 582280
rect 126130 582240 126140 582280
rect 126080 582170 126140 582240
rect 126200 582280 126260 582300
rect 126200 582240 126210 582280
rect 126250 582240 126260 582280
rect 126200 582170 126260 582240
rect 126300 582280 126430 582300
rect 126300 582240 126320 582280
rect 126410 582240 126430 582280
rect 126300 582220 126430 582240
rect 126470 582280 126530 582300
rect 126470 582240 126480 582280
rect 126520 582240 126530 582280
rect 126470 582170 126530 582240
rect 126590 582280 126650 582300
rect 126590 582240 126600 582280
rect 126640 582240 126650 582280
rect 126590 582170 126650 582240
rect 126690 582280 126820 582300
rect 126690 582240 126710 582280
rect 126800 582240 126820 582280
rect 126690 582220 126820 582240
rect 126860 582280 126920 582300
rect 126860 582240 126870 582280
rect 126910 582240 126920 582280
rect 126860 582170 126920 582240
rect 126980 582280 127040 582300
rect 126980 582240 126990 582280
rect 127030 582240 127040 582280
rect 126980 582170 127040 582240
rect 127080 582280 127210 582300
rect 127080 582240 127100 582280
rect 127190 582240 127210 582280
rect 127080 582220 127210 582240
rect 127250 582280 127310 582300
rect 127250 582240 127260 582280
rect 127300 582240 127310 582280
rect 127250 582170 127310 582240
rect 127370 582280 127430 582300
rect 127370 582240 127380 582280
rect 127420 582240 127430 582280
rect 127370 582170 127430 582240
rect 127470 582280 127600 582300
rect 127470 582240 127490 582280
rect 127580 582240 127600 582280
rect 127470 582220 127600 582240
rect 127640 582280 127700 582300
rect 127640 582240 127650 582280
rect 127690 582240 127700 582280
rect 127640 582170 127700 582240
rect 127760 582280 127820 582300
rect 127760 582240 127770 582280
rect 127810 582240 127820 582280
rect 127760 582170 127820 582240
rect 127860 582280 127990 582300
rect 127860 582240 127880 582280
rect 127970 582240 127990 582280
rect 127860 582220 127990 582240
rect 128030 582280 128090 582300
rect 128030 582240 128040 582280
rect 128080 582240 128090 582280
rect 128030 582170 128090 582240
rect 128150 582280 128210 582300
rect 128150 582240 128160 582280
rect 128200 582240 128210 582280
rect 128150 582170 128210 582240
rect 128250 582280 128380 582300
rect 128250 582240 128270 582280
rect 128360 582240 128380 582280
rect 128250 582220 128380 582240
rect 128420 582280 128480 582300
rect 128420 582240 128430 582280
rect 128470 582240 128480 582280
rect 128420 582170 128480 582240
rect 128540 582280 128600 582300
rect 128540 582240 128550 582280
rect 128590 582240 128600 582280
rect 128540 582170 128600 582240
rect 128640 582280 128770 582300
rect 128640 582240 128660 582280
rect 128750 582240 128770 582280
rect 128640 582220 128770 582240
rect 128810 582280 128870 582300
rect 128810 582240 128820 582280
rect 128860 582240 128870 582280
rect 128810 582170 128870 582240
rect 128930 582280 128990 582300
rect 128930 582240 128940 582280
rect 128980 582240 128990 582280
rect 128930 582170 128990 582240
rect 129030 582280 129160 582300
rect 129030 582240 129050 582280
rect 129140 582240 129160 582280
rect 129030 582220 129160 582240
rect 129200 582280 129260 582300
rect 129200 582240 129210 582280
rect 129250 582240 129260 582280
rect 129200 582170 129260 582240
rect 129320 582280 129380 582300
rect 129320 582240 129330 582280
rect 129370 582240 129380 582280
rect 129320 582170 129380 582240
rect 129420 582280 129550 582300
rect 129420 582240 129440 582280
rect 129530 582240 129550 582280
rect 129420 582220 129550 582240
rect 129590 582280 129650 582300
rect 129590 582240 129600 582280
rect 129640 582240 129650 582280
rect 129590 582170 129650 582240
rect 129710 582280 129770 582300
rect 129710 582240 129720 582280
rect 129760 582240 129770 582280
rect 129710 582170 129770 582240
rect 129810 582280 129940 582300
rect 129810 582240 129830 582280
rect 129920 582240 129940 582280
rect 129810 582220 129940 582240
rect 129980 582280 130040 582300
rect 129980 582240 129990 582280
rect 130030 582240 130040 582280
rect 129980 582170 130040 582240
rect 130100 582280 130160 582300
rect 130100 582240 130110 582280
rect 130150 582240 130160 582280
rect 130100 582170 130160 582240
rect 130200 582280 130330 582300
rect 130200 582240 130220 582280
rect 130310 582240 130330 582280
rect 130200 582220 130330 582240
rect 130370 582280 130430 582300
rect 130370 582240 130380 582280
rect 130420 582240 130430 582280
rect 130370 582170 130430 582240
rect 130490 582280 130550 582300
rect 130490 582240 130500 582280
rect 130540 582240 130550 582280
rect 130490 582170 130550 582240
rect 130590 582280 130720 582300
rect 130590 582240 130610 582280
rect 130700 582240 130720 582280
rect 130590 582220 130720 582240
rect 130760 582280 130820 582300
rect 130760 582240 130770 582280
rect 130810 582240 130820 582280
rect 130760 582170 130820 582240
rect 130880 582280 130940 582300
rect 130880 582240 130890 582280
rect 130930 582240 130940 582280
rect 130880 582170 130940 582240
rect 130980 582280 131110 582300
rect 130980 582240 131000 582280
rect 131090 582240 131110 582280
rect 130980 582220 131110 582240
rect 131150 582280 131210 582300
rect 131150 582240 131160 582280
rect 131200 582240 131210 582280
rect 131150 582170 131210 582240
rect 131270 582280 131330 582300
rect 131270 582240 131280 582280
rect 131320 582240 131330 582280
rect 131270 582170 131330 582240
rect 131370 582280 131500 582300
rect 131370 582240 131390 582280
rect 131480 582240 131500 582280
rect 131370 582220 131500 582240
rect 131540 582280 131600 582300
rect 131540 582240 131550 582280
rect 131590 582240 131600 582280
rect 131540 582170 131600 582240
rect 131660 582280 131720 582300
rect 131660 582240 131670 582280
rect 131710 582240 131720 582280
rect 131660 582170 131720 582240
rect 131760 582280 131890 582300
rect 131760 582240 131780 582280
rect 131870 582240 131890 582280
rect 131760 582220 131890 582240
rect 131930 582280 131990 582300
rect 131930 582240 131940 582280
rect 131980 582240 131990 582280
rect 131930 582170 131990 582240
rect 132050 582280 132110 582300
rect 132050 582240 132060 582280
rect 132100 582240 132110 582280
rect 132050 582170 132110 582240
rect 132150 582280 132280 582300
rect 132150 582240 132170 582280
rect 132260 582240 132280 582280
rect 132150 582220 132280 582240
rect 132320 582280 132380 582300
rect 132320 582240 132330 582280
rect 132370 582240 132380 582280
rect 132320 582170 132380 582240
rect 132440 582280 132500 582300
rect 132440 582240 132450 582280
rect 132490 582240 132500 582280
rect 132440 582170 132500 582240
rect 132540 582280 132670 582300
rect 132540 582240 132560 582280
rect 132650 582240 132670 582280
rect 132540 582220 132670 582240
rect 132710 582280 132770 582300
rect 132710 582240 132720 582280
rect 132760 582240 132770 582280
rect 132710 582170 132770 582240
rect 125420 582110 128370 582170
rect 128870 582110 132770 582170
rect 132860 581950 132890 582520
rect 133020 581950 133050 582520
rect 132860 581930 133050 581950
rect 119330 575566 119430 575608
rect 119312 575560 119430 575566
rect 119312 575480 119318 575560
rect 119410 575480 119430 575560
rect 119312 575442 119430 575480
rect 119130 575178 119230 575186
rect 119130 575094 119138 575178
rect 119220 575100 119230 575178
rect 119220 575094 119270 575100
rect 119130 575080 119270 575094
rect 119170 574870 119270 575080
rect 119170 574810 119190 574870
rect 119250 574810 119270 574870
rect 119170 574790 119270 574810
rect 119330 574390 119430 575442
rect 119490 575090 120114 575100
rect 119490 575084 120130 575090
rect 119490 575004 120036 575084
rect 120128 575004 120130 575084
rect 119490 575000 120130 575004
rect 119490 574980 119590 575000
rect 119490 574920 119510 574980
rect 119570 574920 119590 574980
rect 120030 574966 120130 575000
rect 119490 574900 119590 574920
rect 119920 574480 120020 574500
rect 120290 574480 120390 574490
rect 119920 574420 119940 574480
rect 120000 574470 120390 574480
rect 120000 574420 120310 574470
rect 119920 574400 120020 574420
rect 120290 574410 120310 574420
rect 120370 574410 120390 574470
rect 120290 574390 120390 574410
rect 119330 574340 119350 574390
rect 119390 574340 119430 574390
rect 119330 573960 119430 574340
rect 119680 574320 119780 574330
rect 119680 574240 119690 574320
rect 119770 574240 119780 574320
rect 119680 574230 119780 574240
rect 119920 574310 124382 574330
rect 119920 574250 119940 574310
rect 120000 574250 124382 574310
rect 119920 574230 124382 574250
rect 119330 573900 119350 573960
rect 119410 573900 119430 573960
rect 119330 573890 119430 573900
rect 124282 573524 124382 574230
rect 125340 574090 125760 574150
rect 125500 574060 125560 574090
rect 125390 574040 125450 574060
rect 125390 574000 125400 574040
rect 125440 574000 125450 574040
rect 125390 573870 125450 574000
rect 125490 574040 125570 574060
rect 125490 574000 125510 574040
rect 125550 574000 125570 574040
rect 125490 573980 125570 574000
rect 125610 574040 125670 574060
rect 125610 574000 125620 574040
rect 125660 574000 125670 574040
rect 125610 573870 125670 574000
rect 124282 573460 132758 573524
rect 124282 573424 125680 573460
rect 125670 573420 125680 573424
rect 125720 573424 126070 573460
rect 125720 573420 125730 573424
rect 125670 573400 125730 573420
rect 126060 573420 126070 573424
rect 126110 573424 126460 573460
rect 126110 573420 126120 573424
rect 126060 573400 126120 573420
rect 126450 573420 126460 573424
rect 126500 573424 126850 573460
rect 126500 573420 126510 573424
rect 126450 573400 126510 573420
rect 126840 573420 126850 573424
rect 126890 573424 127240 573460
rect 126890 573420 126900 573424
rect 126840 573400 126900 573420
rect 127230 573420 127240 573424
rect 127280 573424 127630 573460
rect 127280 573420 127290 573424
rect 127230 573400 127290 573420
rect 127620 573420 127630 573424
rect 127670 573424 128020 573460
rect 127670 573420 127680 573424
rect 127620 573400 127680 573420
rect 128010 573420 128020 573424
rect 128060 573424 128410 573460
rect 128060 573420 128070 573424
rect 128010 573400 128070 573420
rect 128400 573420 128410 573424
rect 128450 573424 128800 573460
rect 128450 573420 128460 573424
rect 128400 573400 128460 573420
rect 128790 573420 128800 573424
rect 128840 573424 129190 573460
rect 128840 573420 128850 573424
rect 128790 573400 128850 573420
rect 129180 573420 129190 573424
rect 129230 573424 129580 573460
rect 129230 573420 129240 573424
rect 129180 573400 129240 573420
rect 129570 573420 129580 573424
rect 129620 573424 129970 573460
rect 129620 573420 129630 573424
rect 129570 573400 129630 573420
rect 129960 573420 129970 573424
rect 130010 573424 130360 573460
rect 130010 573420 130020 573424
rect 129960 573400 130020 573420
rect 130350 573420 130360 573424
rect 130400 573424 130750 573460
rect 130400 573420 130410 573424
rect 130350 573400 130410 573420
rect 130740 573420 130750 573424
rect 130790 573424 131140 573460
rect 130790 573420 130800 573424
rect 130740 573400 130800 573420
rect 131130 573420 131140 573424
rect 131180 573424 131530 573460
rect 131180 573420 131190 573424
rect 131130 573400 131190 573420
rect 131520 573420 131530 573424
rect 131570 573424 131920 573460
rect 131570 573420 131580 573424
rect 131520 573400 131580 573420
rect 131910 573420 131920 573424
rect 131960 573424 132310 573460
rect 131960 573420 131970 573424
rect 131910 573400 131970 573420
rect 132300 573420 132310 573424
rect 132350 573424 132700 573460
rect 132350 573420 132360 573424
rect 132300 573400 132360 573420
rect 132690 573420 132700 573424
rect 132740 573424 132758 573460
rect 132900 573500 133090 573520
rect 132740 573420 132750 573424
rect 132690 573400 132750 573420
rect 125400 573310 128410 573370
rect 128910 573310 132810 573370
rect 125570 573280 125680 573310
rect 125960 573280 126070 573310
rect 126350 573280 126460 573310
rect 126740 573280 126850 573310
rect 127130 573280 127240 573310
rect 127520 573280 127630 573310
rect 127910 573280 128020 573310
rect 128300 573280 128410 573310
rect 128690 573280 128800 573310
rect 129080 573280 129190 573310
rect 129470 573280 129580 573310
rect 129860 573280 129970 573310
rect 130250 573280 130360 573310
rect 130640 573280 130750 573310
rect 131030 573280 131140 573310
rect 131420 573280 131530 573310
rect 131810 573280 131920 573310
rect 132200 573280 132310 573310
rect 132590 573280 132700 573310
rect 125460 573260 125520 573280
rect 125460 573120 125470 573260
rect 125510 573120 125520 573260
rect 125460 573050 125520 573120
rect 125560 573260 125690 573280
rect 125560 573120 125580 573260
rect 125670 573120 125690 573260
rect 125560 573100 125690 573120
rect 125730 573260 125790 573280
rect 125730 573120 125740 573260
rect 125780 573120 125790 573260
rect 125730 573050 125790 573120
rect 125850 573260 125910 573280
rect 125850 573120 125860 573260
rect 125900 573120 125910 573260
rect 125850 573050 125910 573120
rect 125950 573260 126080 573280
rect 125950 573120 125970 573260
rect 126060 573120 126080 573260
rect 125950 573100 126080 573120
rect 126120 573260 126180 573280
rect 126120 573120 126130 573260
rect 126170 573120 126180 573260
rect 126120 573050 126180 573120
rect 126240 573260 126300 573280
rect 126240 573120 126250 573260
rect 126290 573120 126300 573260
rect 126240 573050 126300 573120
rect 126340 573260 126470 573280
rect 126340 573120 126360 573260
rect 126450 573120 126470 573260
rect 126340 573100 126470 573120
rect 126510 573260 126570 573280
rect 126510 573120 126520 573260
rect 126560 573120 126570 573260
rect 126510 573050 126570 573120
rect 126630 573260 126690 573280
rect 126630 573120 126640 573260
rect 126680 573120 126690 573260
rect 126630 573050 126690 573120
rect 126730 573260 126860 573280
rect 126730 573120 126750 573260
rect 126840 573120 126860 573260
rect 126730 573100 126860 573120
rect 126900 573260 126960 573280
rect 126900 573120 126910 573260
rect 126950 573120 126960 573260
rect 126900 573050 126960 573120
rect 127020 573260 127080 573280
rect 127020 573120 127030 573260
rect 127070 573120 127080 573260
rect 127020 573050 127080 573120
rect 127120 573260 127250 573280
rect 127120 573120 127140 573260
rect 127230 573120 127250 573260
rect 127120 573100 127250 573120
rect 127290 573260 127350 573280
rect 127290 573120 127300 573260
rect 127340 573120 127350 573260
rect 127290 573050 127350 573120
rect 127410 573260 127470 573280
rect 127410 573120 127420 573260
rect 127460 573120 127470 573260
rect 127410 573050 127470 573120
rect 127510 573260 127640 573280
rect 127510 573120 127530 573260
rect 127620 573120 127640 573260
rect 127510 573100 127640 573120
rect 127680 573260 127740 573280
rect 127680 573120 127690 573260
rect 127730 573120 127740 573260
rect 127680 573050 127740 573120
rect 127800 573260 127860 573280
rect 127800 573120 127810 573260
rect 127850 573120 127860 573260
rect 127800 573050 127860 573120
rect 127900 573260 128030 573280
rect 127900 573120 127920 573260
rect 128010 573120 128030 573260
rect 127900 573100 128030 573120
rect 128070 573260 128130 573280
rect 128070 573120 128080 573260
rect 128120 573120 128130 573260
rect 128070 573050 128130 573120
rect 128190 573260 128250 573280
rect 128190 573120 128200 573260
rect 128240 573120 128250 573260
rect 128190 573050 128250 573120
rect 128290 573260 128420 573280
rect 128290 573120 128310 573260
rect 128400 573120 128420 573260
rect 128290 573100 128420 573120
rect 128460 573260 128520 573280
rect 128460 573120 128470 573260
rect 128510 573120 128520 573260
rect 128460 573050 128520 573120
rect 128580 573260 128640 573280
rect 128580 573120 128590 573260
rect 128630 573120 128640 573260
rect 128580 573050 128640 573120
rect 128680 573260 128810 573280
rect 128680 573120 128700 573260
rect 128790 573120 128810 573260
rect 128680 573100 128810 573120
rect 128850 573260 128910 573280
rect 128850 573120 128860 573260
rect 128900 573120 128910 573260
rect 128850 573050 128910 573120
rect 128970 573260 129030 573280
rect 128970 573120 128980 573260
rect 129020 573120 129030 573260
rect 128970 573050 129030 573120
rect 129070 573260 129200 573280
rect 129070 573120 129090 573260
rect 129180 573120 129200 573260
rect 129070 573100 129200 573120
rect 129240 573260 129300 573280
rect 129240 573120 129250 573260
rect 129290 573120 129300 573260
rect 129240 573050 129300 573120
rect 129360 573260 129420 573280
rect 129360 573120 129370 573260
rect 129410 573120 129420 573260
rect 129360 573050 129420 573120
rect 129460 573260 129590 573280
rect 129460 573120 129480 573260
rect 129570 573120 129590 573260
rect 129460 573100 129590 573120
rect 129630 573260 129690 573280
rect 129630 573120 129640 573260
rect 129680 573120 129690 573260
rect 129630 573050 129690 573120
rect 129750 573260 129810 573280
rect 129750 573120 129760 573260
rect 129800 573120 129810 573260
rect 129750 573050 129810 573120
rect 129850 573260 129980 573280
rect 129850 573120 129870 573260
rect 129960 573120 129980 573260
rect 129850 573100 129980 573120
rect 130020 573260 130080 573280
rect 130020 573120 130030 573260
rect 130070 573120 130080 573260
rect 130020 573050 130080 573120
rect 130140 573260 130200 573280
rect 130140 573120 130150 573260
rect 130190 573120 130200 573260
rect 130140 573050 130200 573120
rect 130240 573260 130370 573280
rect 130240 573120 130260 573260
rect 130350 573120 130370 573260
rect 130240 573100 130370 573120
rect 130410 573260 130470 573280
rect 130410 573120 130420 573260
rect 130460 573120 130470 573260
rect 130410 573050 130470 573120
rect 130530 573260 130590 573280
rect 130530 573120 130540 573260
rect 130580 573120 130590 573260
rect 130530 573050 130590 573120
rect 130630 573260 130760 573280
rect 130630 573120 130650 573260
rect 130740 573120 130760 573260
rect 130630 573100 130760 573120
rect 130800 573260 130860 573280
rect 130800 573120 130810 573260
rect 130850 573120 130860 573260
rect 130800 573050 130860 573120
rect 130920 573260 130980 573280
rect 130920 573120 130930 573260
rect 130970 573120 130980 573260
rect 130920 573050 130980 573120
rect 131020 573260 131150 573280
rect 131020 573120 131040 573260
rect 131130 573120 131150 573260
rect 131020 573100 131150 573120
rect 131190 573260 131250 573280
rect 131190 573120 131200 573260
rect 131240 573120 131250 573260
rect 131190 573050 131250 573120
rect 131310 573260 131370 573280
rect 131310 573120 131320 573260
rect 131360 573120 131370 573260
rect 131310 573050 131370 573120
rect 131410 573260 131540 573280
rect 131410 573120 131430 573260
rect 131520 573120 131540 573260
rect 131410 573100 131540 573120
rect 131580 573260 131640 573280
rect 131580 573120 131590 573260
rect 131630 573120 131640 573260
rect 131580 573050 131640 573120
rect 131700 573260 131760 573280
rect 131700 573120 131710 573260
rect 131750 573120 131760 573260
rect 131700 573050 131760 573120
rect 131800 573260 131930 573280
rect 131800 573120 131820 573260
rect 131910 573120 131930 573260
rect 131800 573100 131930 573120
rect 131970 573260 132030 573280
rect 131970 573120 131980 573260
rect 132020 573120 132030 573260
rect 131970 573050 132030 573120
rect 132090 573260 132150 573280
rect 132090 573120 132100 573260
rect 132140 573120 132150 573260
rect 132090 573050 132150 573120
rect 132190 573260 132320 573280
rect 132190 573120 132210 573260
rect 132300 573120 132320 573260
rect 132190 573100 132320 573120
rect 132360 573260 132420 573280
rect 132360 573120 132370 573260
rect 132410 573120 132420 573260
rect 132360 573050 132420 573120
rect 132480 573260 132540 573280
rect 132480 573120 132490 573260
rect 132530 573120 132540 573260
rect 132480 573050 132540 573120
rect 132580 573260 132710 573280
rect 132580 573120 132600 573260
rect 132690 573120 132710 573260
rect 132580 573100 132710 573120
rect 132750 573260 132810 573280
rect 132750 573120 132760 573260
rect 132800 573120 132810 573260
rect 132750 573050 132810 573120
rect 125460 572990 128410 573050
rect 128910 572990 132810 573050
rect 132900 572830 132930 573500
rect 133060 572830 133090 573500
rect 132900 572810 133090 572830
rect 119368 568042 119468 568048
rect 119368 568024 119374 568042
rect 119280 567962 119374 568024
rect 119466 568024 119468 568042
rect 119466 567962 119484 568024
rect 119280 567924 119484 567962
rect 119126 567510 119226 567518
rect 119126 567430 119134 567510
rect 119120 567426 119134 567430
rect 119216 567426 119226 567510
rect 119120 567412 119226 567426
rect 119120 567200 119220 567412
rect 119120 567140 119140 567200
rect 119200 567140 119220 567200
rect 119120 567120 119220 567140
rect 119280 566720 119380 567924
rect 119440 567388 120046 567430
rect 119440 567382 120088 567388
rect 119440 567330 119994 567382
rect 119440 567310 119540 567330
rect 119440 567250 119460 567310
rect 119520 567250 119540 567310
rect 119988 567302 119994 567330
rect 120086 567302 120088 567382
rect 119988 567264 120088 567302
rect 119440 567230 119540 567250
rect 119870 566810 119970 566830
rect 120240 566810 120340 566820
rect 119870 566750 119890 566810
rect 119950 566800 120340 566810
rect 119950 566750 120260 566800
rect 119870 566730 119970 566750
rect 120240 566740 120260 566750
rect 120320 566740 120340 566800
rect 120240 566720 120340 566740
rect 119280 566670 119300 566720
rect 119340 566670 119380 566720
rect 119280 566290 119380 566670
rect 119630 566650 119730 566660
rect 119630 566570 119640 566650
rect 119720 566570 119730 566650
rect 119630 566560 119730 566570
rect 119870 566640 124332 566660
rect 119870 566580 119890 566640
rect 119950 566580 124332 566640
rect 119870 566560 124332 566580
rect 119280 566230 119300 566290
rect 119360 566230 119380 566290
rect 119280 566220 119380 566230
rect 124232 565854 124332 566560
rect 125290 566420 125710 566480
rect 125450 566390 125510 566420
rect 125340 566370 125400 566390
rect 125340 566330 125350 566370
rect 125390 566330 125400 566370
rect 125340 566200 125400 566330
rect 125440 566370 125520 566390
rect 125440 566330 125460 566370
rect 125500 566330 125520 566370
rect 125440 566310 125520 566330
rect 125560 566370 125620 566390
rect 125560 566330 125570 566370
rect 125610 566330 125620 566370
rect 125560 566200 125620 566330
rect 124232 565790 132708 565854
rect 124232 565754 125630 565790
rect 125620 565750 125630 565754
rect 125670 565754 126020 565790
rect 125670 565750 125680 565754
rect 125620 565730 125680 565750
rect 126010 565750 126020 565754
rect 126060 565754 126410 565790
rect 126060 565750 126070 565754
rect 126010 565730 126070 565750
rect 126400 565750 126410 565754
rect 126450 565754 126800 565790
rect 126450 565750 126460 565754
rect 126400 565730 126460 565750
rect 126790 565750 126800 565754
rect 126840 565754 127190 565790
rect 126840 565750 126850 565754
rect 126790 565730 126850 565750
rect 127180 565750 127190 565754
rect 127230 565754 127580 565790
rect 127230 565750 127240 565754
rect 127180 565730 127240 565750
rect 127570 565750 127580 565754
rect 127620 565754 127970 565790
rect 127620 565750 127630 565754
rect 127570 565730 127630 565750
rect 127960 565750 127970 565754
rect 128010 565754 128360 565790
rect 128010 565750 128020 565754
rect 127960 565730 128020 565750
rect 128350 565750 128360 565754
rect 128400 565754 128750 565790
rect 128400 565750 128410 565754
rect 128350 565730 128410 565750
rect 128740 565750 128750 565754
rect 128790 565754 129140 565790
rect 128790 565750 128800 565754
rect 128740 565730 128800 565750
rect 129130 565750 129140 565754
rect 129180 565754 129530 565790
rect 129180 565750 129190 565754
rect 129130 565730 129190 565750
rect 129520 565750 129530 565754
rect 129570 565754 129920 565790
rect 129570 565750 129580 565754
rect 129520 565730 129580 565750
rect 129910 565750 129920 565754
rect 129960 565754 130310 565790
rect 129960 565750 129970 565754
rect 129910 565730 129970 565750
rect 130300 565750 130310 565754
rect 130350 565754 130700 565790
rect 130350 565750 130360 565754
rect 130300 565730 130360 565750
rect 130690 565750 130700 565754
rect 130740 565754 131090 565790
rect 130740 565750 130750 565754
rect 130690 565730 130750 565750
rect 131080 565750 131090 565754
rect 131130 565754 131480 565790
rect 131130 565750 131140 565754
rect 131080 565730 131140 565750
rect 131470 565750 131480 565754
rect 131520 565754 131870 565790
rect 131520 565750 131530 565754
rect 131470 565730 131530 565750
rect 131860 565750 131870 565754
rect 131910 565754 132260 565790
rect 131910 565750 131920 565754
rect 131860 565730 131920 565750
rect 132250 565750 132260 565754
rect 132300 565754 132650 565790
rect 132300 565750 132310 565754
rect 132250 565730 132310 565750
rect 132640 565750 132650 565754
rect 132690 565754 132708 565790
rect 132850 565830 133040 565850
rect 132690 565750 132700 565754
rect 132640 565730 132700 565750
rect 125350 565640 128360 565700
rect 128860 565640 132760 565700
rect 125520 565610 125630 565640
rect 125910 565610 126020 565640
rect 126300 565610 126410 565640
rect 126690 565610 126800 565640
rect 127080 565610 127190 565640
rect 127470 565610 127580 565640
rect 127860 565610 127970 565640
rect 128250 565610 128360 565640
rect 128640 565610 128750 565640
rect 129030 565610 129140 565640
rect 129420 565610 129530 565640
rect 129810 565610 129920 565640
rect 130200 565610 130310 565640
rect 130590 565610 130700 565640
rect 130980 565610 131090 565640
rect 131370 565610 131480 565640
rect 131760 565610 131870 565640
rect 132150 565610 132260 565640
rect 132540 565610 132650 565640
rect 125410 565590 125470 565610
rect 125410 565350 125420 565590
rect 125460 565350 125470 565590
rect 125410 565280 125470 565350
rect 125510 565590 125640 565610
rect 125510 565350 125530 565590
rect 125620 565350 125640 565590
rect 125510 565330 125640 565350
rect 125680 565590 125740 565610
rect 125680 565350 125690 565590
rect 125730 565350 125740 565590
rect 125680 565280 125740 565350
rect 125800 565590 125860 565610
rect 125800 565350 125810 565590
rect 125850 565350 125860 565590
rect 125800 565280 125860 565350
rect 125900 565590 126030 565610
rect 125900 565350 125920 565590
rect 126010 565350 126030 565590
rect 125900 565330 126030 565350
rect 126070 565590 126130 565610
rect 126070 565350 126080 565590
rect 126120 565350 126130 565590
rect 126070 565280 126130 565350
rect 126190 565590 126250 565610
rect 126190 565350 126200 565590
rect 126240 565350 126250 565590
rect 126190 565280 126250 565350
rect 126290 565590 126420 565610
rect 126290 565350 126310 565590
rect 126400 565350 126420 565590
rect 126290 565330 126420 565350
rect 126460 565590 126520 565610
rect 126460 565350 126470 565590
rect 126510 565350 126520 565590
rect 126460 565280 126520 565350
rect 126580 565590 126640 565610
rect 126580 565350 126590 565590
rect 126630 565350 126640 565590
rect 126580 565280 126640 565350
rect 126680 565590 126810 565610
rect 126680 565350 126700 565590
rect 126790 565350 126810 565590
rect 126680 565330 126810 565350
rect 126850 565590 126910 565610
rect 126850 565350 126860 565590
rect 126900 565350 126910 565590
rect 126850 565280 126910 565350
rect 126970 565590 127030 565610
rect 126970 565350 126980 565590
rect 127020 565350 127030 565590
rect 126970 565280 127030 565350
rect 127070 565590 127200 565610
rect 127070 565350 127090 565590
rect 127180 565350 127200 565590
rect 127070 565330 127200 565350
rect 127240 565590 127300 565610
rect 127240 565350 127250 565590
rect 127290 565350 127300 565590
rect 127240 565280 127300 565350
rect 127360 565590 127420 565610
rect 127360 565350 127370 565590
rect 127410 565350 127420 565590
rect 127360 565280 127420 565350
rect 127460 565590 127590 565610
rect 127460 565350 127480 565590
rect 127570 565350 127590 565590
rect 127460 565330 127590 565350
rect 127630 565590 127690 565610
rect 127630 565350 127640 565590
rect 127680 565350 127690 565590
rect 127630 565280 127690 565350
rect 127750 565590 127810 565610
rect 127750 565350 127760 565590
rect 127800 565350 127810 565590
rect 127750 565280 127810 565350
rect 127850 565590 127980 565610
rect 127850 565350 127870 565590
rect 127960 565350 127980 565590
rect 127850 565330 127980 565350
rect 128020 565590 128080 565610
rect 128020 565350 128030 565590
rect 128070 565350 128080 565590
rect 128020 565280 128080 565350
rect 128140 565590 128200 565610
rect 128140 565350 128150 565590
rect 128190 565350 128200 565590
rect 128140 565280 128200 565350
rect 128240 565590 128370 565610
rect 128240 565350 128260 565590
rect 128350 565350 128370 565590
rect 128240 565330 128370 565350
rect 128410 565590 128470 565610
rect 128410 565350 128420 565590
rect 128460 565350 128470 565590
rect 128410 565280 128470 565350
rect 128530 565590 128590 565610
rect 128530 565350 128540 565590
rect 128580 565350 128590 565590
rect 128530 565280 128590 565350
rect 128630 565590 128760 565610
rect 128630 565350 128650 565590
rect 128740 565350 128760 565590
rect 128630 565330 128760 565350
rect 128800 565590 128860 565610
rect 128800 565350 128810 565590
rect 128850 565350 128860 565590
rect 128800 565280 128860 565350
rect 128920 565590 128980 565610
rect 128920 565350 128930 565590
rect 128970 565350 128980 565590
rect 128920 565280 128980 565350
rect 129020 565590 129150 565610
rect 129020 565350 129040 565590
rect 129130 565350 129150 565590
rect 129020 565330 129150 565350
rect 129190 565590 129250 565610
rect 129190 565350 129200 565590
rect 129240 565350 129250 565590
rect 129190 565280 129250 565350
rect 129310 565590 129370 565610
rect 129310 565350 129320 565590
rect 129360 565350 129370 565590
rect 129310 565280 129370 565350
rect 129410 565590 129540 565610
rect 129410 565350 129430 565590
rect 129520 565350 129540 565590
rect 129410 565330 129540 565350
rect 129580 565590 129640 565610
rect 129580 565350 129590 565590
rect 129630 565350 129640 565590
rect 129580 565280 129640 565350
rect 129700 565590 129760 565610
rect 129700 565350 129710 565590
rect 129750 565350 129760 565590
rect 129700 565280 129760 565350
rect 129800 565590 129930 565610
rect 129800 565350 129820 565590
rect 129910 565350 129930 565590
rect 129800 565330 129930 565350
rect 129970 565590 130030 565610
rect 129970 565350 129980 565590
rect 130020 565350 130030 565590
rect 129970 565280 130030 565350
rect 130090 565590 130150 565610
rect 130090 565350 130100 565590
rect 130140 565350 130150 565590
rect 130090 565280 130150 565350
rect 130190 565590 130320 565610
rect 130190 565350 130210 565590
rect 130300 565350 130320 565590
rect 130190 565330 130320 565350
rect 130360 565590 130420 565610
rect 130360 565350 130370 565590
rect 130410 565350 130420 565590
rect 130360 565280 130420 565350
rect 130480 565590 130540 565610
rect 130480 565350 130490 565590
rect 130530 565350 130540 565590
rect 130480 565280 130540 565350
rect 130580 565590 130710 565610
rect 130580 565350 130600 565590
rect 130690 565350 130710 565590
rect 130580 565330 130710 565350
rect 130750 565590 130810 565610
rect 130750 565350 130760 565590
rect 130800 565350 130810 565590
rect 130750 565280 130810 565350
rect 130870 565590 130930 565610
rect 130870 565350 130880 565590
rect 130920 565350 130930 565590
rect 130870 565280 130930 565350
rect 130970 565590 131100 565610
rect 130970 565350 130990 565590
rect 131080 565350 131100 565590
rect 130970 565330 131100 565350
rect 131140 565590 131200 565610
rect 131140 565350 131150 565590
rect 131190 565350 131200 565590
rect 131140 565280 131200 565350
rect 131260 565590 131320 565610
rect 131260 565350 131270 565590
rect 131310 565350 131320 565590
rect 131260 565280 131320 565350
rect 131360 565590 131490 565610
rect 131360 565350 131380 565590
rect 131470 565350 131490 565590
rect 131360 565330 131490 565350
rect 131530 565590 131590 565610
rect 131530 565350 131540 565590
rect 131580 565350 131590 565590
rect 131530 565280 131590 565350
rect 131650 565590 131710 565610
rect 131650 565350 131660 565590
rect 131700 565350 131710 565590
rect 131650 565280 131710 565350
rect 131750 565590 131880 565610
rect 131750 565350 131770 565590
rect 131860 565350 131880 565590
rect 131750 565330 131880 565350
rect 131920 565590 131980 565610
rect 131920 565350 131930 565590
rect 131970 565350 131980 565590
rect 131920 565280 131980 565350
rect 132040 565590 132100 565610
rect 132040 565350 132050 565590
rect 132090 565350 132100 565590
rect 132040 565280 132100 565350
rect 132140 565590 132270 565610
rect 132140 565350 132160 565590
rect 132250 565350 132270 565590
rect 132140 565330 132270 565350
rect 132310 565590 132370 565610
rect 132310 565350 132320 565590
rect 132360 565350 132370 565590
rect 132310 565280 132370 565350
rect 132430 565590 132490 565610
rect 132430 565350 132440 565590
rect 132480 565350 132490 565590
rect 132430 565280 132490 565350
rect 132530 565590 132660 565610
rect 132530 565350 132550 565590
rect 132640 565350 132660 565590
rect 132530 565330 132660 565350
rect 132700 565590 132760 565610
rect 132700 565350 132710 565590
rect 132750 565350 132760 565590
rect 132700 565280 132760 565350
rect 125410 565220 128360 565280
rect 128860 565220 132760 565280
rect 132850 565060 132880 565830
rect 133010 565060 133040 565830
rect 132850 565040 133040 565060
rect 311944 561524 312040 563752
rect 119308 561424 119408 561430
rect 119308 561388 119314 561424
rect 119280 561344 119314 561388
rect 119406 561344 119408 561424
rect 119280 561306 119408 561344
rect 311944 561428 312200 561524
rect 119116 560948 119216 560956
rect 119116 560864 119124 560948
rect 119206 560890 119216 560948
rect 119206 560864 119220 560890
rect 119116 560850 119220 560864
rect 119120 560660 119220 560850
rect 119120 560600 119140 560660
rect 119200 560600 119220 560660
rect 119120 560580 119220 560600
rect 119280 560180 119380 561306
rect 120028 560958 120128 560960
rect 119440 560954 120128 560958
rect 119440 560874 120034 560954
rect 120126 560874 120128 560954
rect 119440 560858 120128 560874
rect 119440 560770 119540 560858
rect 120028 560836 120128 560858
rect 119440 560710 119460 560770
rect 119520 560710 119540 560770
rect 119440 560690 119540 560710
rect 311944 560570 312038 561428
rect 370436 560977 371064 560980
rect 371755 560977 371851 563752
rect 375661 561624 375757 563752
rect 435472 561925 435568 563752
rect 435472 561817 435568 561829
rect 375661 561539 377172 561624
rect 375662 561528 377172 561539
rect 370436 560884 371851 560977
rect 311942 560436 312038 560570
rect 370968 560881 371851 560884
rect 311942 560340 312200 560436
rect 119870 560270 119970 560290
rect 120240 560270 120340 560280
rect 119870 560210 119890 560270
rect 119950 560260 120340 560270
rect 119950 560210 120260 560260
rect 119870 560190 119970 560210
rect 120240 560200 120260 560210
rect 120320 560200 120340 560260
rect 120240 560180 120340 560200
rect 119280 560130 119300 560180
rect 119340 560130 119380 560180
rect 119280 559750 119380 560130
rect 119630 560110 119730 560120
rect 119630 560030 119640 560110
rect 119720 560030 119730 560110
rect 119630 560020 119730 560030
rect 119870 560100 124332 560120
rect 119870 560040 119890 560100
rect 119950 560040 124332 560100
rect 119870 560020 124332 560040
rect 119280 559690 119300 559750
rect 119360 559690 119380 559750
rect 119280 559680 119380 559690
rect 124232 559314 124332 560020
rect 125290 559880 125710 559940
rect 125450 559850 125510 559880
rect 125340 559830 125400 559850
rect 125340 559790 125350 559830
rect 125390 559790 125400 559830
rect 125340 559660 125400 559790
rect 125440 559830 125520 559850
rect 125440 559790 125460 559830
rect 125500 559790 125520 559830
rect 125440 559770 125520 559790
rect 125560 559830 125620 559850
rect 125560 559790 125570 559830
rect 125610 559790 125620 559830
rect 125560 559660 125620 559790
rect 311942 559348 312038 560340
rect 370968 559892 371064 560881
rect 370436 559796 371064 559892
rect 124232 559250 132708 559314
rect 124232 559214 125630 559250
rect 125620 559210 125630 559214
rect 125670 559214 126020 559250
rect 125670 559210 125680 559214
rect 125620 559190 125680 559210
rect 126010 559210 126020 559214
rect 126060 559214 126410 559250
rect 126060 559210 126070 559214
rect 126010 559190 126070 559210
rect 126400 559210 126410 559214
rect 126450 559214 126800 559250
rect 126450 559210 126460 559214
rect 126400 559190 126460 559210
rect 126790 559210 126800 559214
rect 126840 559214 127190 559250
rect 126840 559210 126850 559214
rect 126790 559190 126850 559210
rect 127180 559210 127190 559214
rect 127230 559214 127580 559250
rect 127230 559210 127240 559214
rect 127180 559190 127240 559210
rect 127570 559210 127580 559214
rect 127620 559214 127970 559250
rect 127620 559210 127630 559214
rect 127570 559190 127630 559210
rect 127960 559210 127970 559214
rect 128010 559214 128360 559250
rect 128010 559210 128020 559214
rect 127960 559190 128020 559210
rect 128350 559210 128360 559214
rect 128400 559214 128750 559250
rect 128400 559210 128410 559214
rect 128350 559190 128410 559210
rect 128740 559210 128750 559214
rect 128790 559214 129140 559250
rect 128790 559210 128800 559214
rect 128740 559190 128800 559210
rect 129130 559210 129140 559214
rect 129180 559214 129530 559250
rect 129180 559210 129190 559214
rect 129130 559190 129190 559210
rect 129520 559210 129530 559214
rect 129570 559214 129920 559250
rect 129570 559210 129580 559214
rect 129520 559190 129580 559210
rect 129910 559210 129920 559214
rect 129960 559214 130310 559250
rect 129960 559210 129970 559214
rect 129910 559190 129970 559210
rect 130300 559210 130310 559214
rect 130350 559214 130700 559250
rect 130350 559210 130360 559214
rect 130300 559190 130360 559210
rect 130690 559210 130700 559214
rect 130740 559214 131090 559250
rect 130740 559210 130750 559214
rect 130690 559190 130750 559210
rect 131080 559210 131090 559214
rect 131130 559214 131480 559250
rect 131130 559210 131140 559214
rect 131080 559190 131140 559210
rect 131470 559210 131480 559214
rect 131520 559214 131870 559250
rect 131520 559210 131530 559214
rect 131470 559190 131530 559210
rect 131860 559210 131870 559214
rect 131910 559214 132260 559250
rect 131910 559210 131920 559214
rect 131860 559190 131920 559210
rect 132250 559210 132260 559214
rect 132300 559214 132650 559250
rect 132300 559210 132310 559214
rect 132250 559190 132310 559210
rect 132640 559210 132650 559214
rect 132690 559214 132708 559250
rect 132850 559290 133040 559310
rect 132690 559210 132700 559214
rect 132640 559190 132700 559210
rect 125350 559100 128360 559160
rect 128860 559100 132760 559160
rect 125520 559070 125630 559100
rect 125910 559070 126020 559100
rect 126300 559070 126410 559100
rect 126690 559070 126800 559100
rect 127080 559070 127190 559100
rect 127470 559070 127580 559100
rect 127860 559070 127970 559100
rect 128250 559070 128360 559100
rect 128640 559070 128750 559100
rect 129030 559070 129140 559100
rect 129420 559070 129530 559100
rect 129810 559070 129920 559100
rect 130200 559070 130310 559100
rect 130590 559070 130700 559100
rect 130980 559070 131090 559100
rect 131370 559070 131480 559100
rect 131760 559070 131870 559100
rect 132150 559070 132260 559100
rect 132540 559070 132650 559100
rect 125410 559050 125470 559070
rect 125410 558710 125420 559050
rect 125460 558710 125470 559050
rect 125410 558640 125470 558710
rect 125510 559050 125640 559070
rect 125510 558710 125530 559050
rect 125620 558710 125640 559050
rect 125510 558690 125640 558710
rect 125680 559050 125740 559070
rect 125680 558710 125690 559050
rect 125730 558710 125740 559050
rect 125680 558640 125740 558710
rect 125800 559050 125860 559070
rect 125800 558710 125810 559050
rect 125850 558710 125860 559050
rect 125800 558640 125860 558710
rect 125900 559050 126030 559070
rect 125900 558710 125920 559050
rect 126010 558710 126030 559050
rect 125900 558690 126030 558710
rect 126070 559050 126130 559070
rect 126070 558710 126080 559050
rect 126120 558710 126130 559050
rect 126070 558640 126130 558710
rect 126190 559050 126250 559070
rect 126190 558710 126200 559050
rect 126240 558710 126250 559050
rect 126190 558640 126250 558710
rect 126290 559050 126420 559070
rect 126290 558710 126310 559050
rect 126400 558710 126420 559050
rect 126290 558690 126420 558710
rect 126460 559050 126520 559070
rect 126460 558710 126470 559050
rect 126510 558710 126520 559050
rect 126460 558640 126520 558710
rect 126580 559050 126640 559070
rect 126580 558710 126590 559050
rect 126630 558710 126640 559050
rect 126580 558640 126640 558710
rect 126680 559050 126810 559070
rect 126680 558710 126700 559050
rect 126790 558710 126810 559050
rect 126680 558690 126810 558710
rect 126850 559050 126910 559070
rect 126850 558710 126860 559050
rect 126900 558710 126910 559050
rect 126850 558640 126910 558710
rect 126970 559050 127030 559070
rect 126970 558710 126980 559050
rect 127020 558710 127030 559050
rect 126970 558640 127030 558710
rect 127070 559050 127200 559070
rect 127070 558710 127090 559050
rect 127180 558710 127200 559050
rect 127070 558690 127200 558710
rect 127240 559050 127300 559070
rect 127240 558710 127250 559050
rect 127290 558710 127300 559050
rect 127240 558640 127300 558710
rect 127360 559050 127420 559070
rect 127360 558710 127370 559050
rect 127410 558710 127420 559050
rect 127360 558640 127420 558710
rect 127460 559050 127590 559070
rect 127460 558710 127480 559050
rect 127570 558710 127590 559050
rect 127460 558690 127590 558710
rect 127630 559050 127690 559070
rect 127630 558710 127640 559050
rect 127680 558710 127690 559050
rect 127630 558640 127690 558710
rect 127750 559050 127810 559070
rect 127750 558710 127760 559050
rect 127800 558710 127810 559050
rect 127750 558640 127810 558710
rect 127850 559050 127980 559070
rect 127850 558710 127870 559050
rect 127960 558710 127980 559050
rect 127850 558690 127980 558710
rect 128020 559050 128080 559070
rect 128020 558710 128030 559050
rect 128070 558710 128080 559050
rect 128020 558640 128080 558710
rect 128140 559050 128200 559070
rect 128140 558710 128150 559050
rect 128190 558710 128200 559050
rect 128140 558640 128200 558710
rect 128240 559050 128370 559070
rect 128240 558710 128260 559050
rect 128350 558710 128370 559050
rect 128240 558690 128370 558710
rect 128410 559050 128470 559070
rect 128410 558710 128420 559050
rect 128460 558710 128470 559050
rect 128410 558640 128470 558710
rect 128530 559050 128590 559070
rect 128530 558710 128540 559050
rect 128580 558710 128590 559050
rect 128530 558640 128590 558710
rect 128630 559050 128760 559070
rect 128630 558710 128650 559050
rect 128740 558710 128760 559050
rect 128630 558690 128760 558710
rect 128800 559050 128860 559070
rect 128800 558710 128810 559050
rect 128850 558710 128860 559050
rect 128800 558640 128860 558710
rect 128920 559050 128980 559070
rect 128920 558710 128930 559050
rect 128970 558710 128980 559050
rect 128920 558640 128980 558710
rect 129020 559050 129150 559070
rect 129020 558710 129040 559050
rect 129130 558710 129150 559050
rect 129020 558690 129150 558710
rect 129190 559050 129250 559070
rect 129190 558710 129200 559050
rect 129240 558710 129250 559050
rect 129190 558640 129250 558710
rect 129310 559050 129370 559070
rect 129310 558710 129320 559050
rect 129360 558710 129370 559050
rect 129310 558640 129370 558710
rect 129410 559050 129540 559070
rect 129410 558710 129430 559050
rect 129520 558710 129540 559050
rect 129410 558690 129540 558710
rect 129580 559050 129640 559070
rect 129580 558710 129590 559050
rect 129630 558710 129640 559050
rect 129580 558640 129640 558710
rect 129700 559050 129760 559070
rect 129700 558710 129710 559050
rect 129750 558710 129760 559050
rect 129700 558640 129760 558710
rect 129800 559050 129930 559070
rect 129800 558710 129820 559050
rect 129910 558710 129930 559050
rect 129800 558690 129930 558710
rect 129970 559050 130030 559070
rect 129970 558710 129980 559050
rect 130020 558710 130030 559050
rect 129970 558640 130030 558710
rect 130090 559050 130150 559070
rect 130090 558710 130100 559050
rect 130140 558710 130150 559050
rect 130090 558640 130150 558710
rect 130190 559050 130320 559070
rect 130190 558710 130210 559050
rect 130300 558710 130320 559050
rect 130190 558690 130320 558710
rect 130360 559050 130420 559070
rect 130360 558710 130370 559050
rect 130410 558710 130420 559050
rect 130360 558640 130420 558710
rect 130480 559050 130540 559070
rect 130480 558710 130490 559050
rect 130530 558710 130540 559050
rect 130480 558640 130540 558710
rect 130580 559050 130710 559070
rect 130580 558710 130600 559050
rect 130690 558710 130710 559050
rect 130580 558690 130710 558710
rect 130750 559050 130810 559070
rect 130750 558710 130760 559050
rect 130800 558710 130810 559050
rect 130750 558640 130810 558710
rect 130870 559050 130930 559070
rect 130870 558710 130880 559050
rect 130920 558710 130930 559050
rect 130870 558640 130930 558710
rect 130970 559050 131100 559070
rect 130970 558710 130990 559050
rect 131080 558710 131100 559050
rect 130970 558690 131100 558710
rect 131140 559050 131200 559070
rect 131140 558710 131150 559050
rect 131190 558710 131200 559050
rect 131140 558640 131200 558710
rect 131260 559050 131320 559070
rect 131260 558710 131270 559050
rect 131310 558710 131320 559050
rect 131260 558640 131320 558710
rect 131360 559050 131490 559070
rect 131360 558710 131380 559050
rect 131470 558710 131490 559050
rect 131360 558690 131490 558710
rect 131530 559050 131590 559070
rect 131530 558710 131540 559050
rect 131580 558710 131590 559050
rect 131530 558640 131590 558710
rect 131650 559050 131710 559070
rect 131650 558710 131660 559050
rect 131700 558710 131710 559050
rect 131650 558640 131710 558710
rect 131750 559050 131880 559070
rect 131750 558710 131770 559050
rect 131860 558710 131880 559050
rect 131750 558690 131880 558710
rect 131920 559050 131980 559070
rect 131920 558710 131930 559050
rect 131970 558710 131980 559050
rect 131920 558640 131980 558710
rect 132040 559050 132100 559070
rect 132040 558710 132050 559050
rect 132090 558710 132100 559050
rect 132040 558640 132100 558710
rect 132140 559050 132270 559070
rect 132140 558710 132160 559050
rect 132250 558710 132270 559050
rect 132140 558690 132270 558710
rect 132310 559050 132370 559070
rect 132310 558710 132320 559050
rect 132360 558710 132370 559050
rect 132310 558640 132370 558710
rect 132430 559050 132490 559070
rect 132430 558710 132440 559050
rect 132480 558710 132490 559050
rect 132430 558640 132490 558710
rect 132530 559050 132660 559070
rect 132530 558710 132550 559050
rect 132640 558710 132660 559050
rect 132530 558690 132660 558710
rect 132700 559050 132760 559070
rect 132700 558710 132710 559050
rect 132750 558710 132760 559050
rect 132700 558640 132760 558710
rect 125410 558580 128360 558640
rect 128860 558580 132760 558640
rect 132850 558420 132880 559290
rect 133010 558420 133040 559290
rect 132850 558400 133040 558420
rect 311942 559252 312200 559348
rect 311942 558260 312038 559252
rect 370968 558804 371064 559796
rect 370436 558708 371064 558804
rect 311942 558164 312200 558260
rect 311942 557172 312038 558164
rect 370968 557716 371064 558708
rect 370436 557620 371064 557716
rect 311942 557076 312200 557172
rect 311942 556084 312038 557076
rect 370968 556628 371064 557620
rect 370436 556532 371064 556628
rect 311942 555988 312200 556084
rect 311942 554996 312038 555988
rect 370968 555540 371064 556532
rect 370436 555444 371064 555540
rect 311942 554900 312200 554996
rect 119344 554640 119444 554646
rect 119344 554560 119350 554640
rect 119442 554594 119444 554640
rect 119442 554560 119450 554594
rect 119344 554522 119450 554560
rect 119124 554062 119224 554070
rect 119124 553978 119132 554062
rect 119214 554060 119224 554062
rect 119214 553978 119290 554060
rect 119124 553964 119290 553978
rect 119190 553830 119290 553964
rect 119190 553770 119210 553830
rect 119270 553770 119290 553830
rect 119190 553750 119290 553770
rect 119350 553350 119450 554522
rect 119510 554038 120156 554060
rect 119510 554032 120172 554038
rect 119510 553960 120078 554032
rect 119510 553940 119610 553960
rect 119510 553880 119530 553940
rect 119590 553880 119610 553940
rect 120072 553952 120078 553960
rect 120170 553952 120172 554032
rect 124940 554020 125360 554080
rect 125100 553990 125160 554020
rect 120072 553914 120172 553952
rect 124990 553970 125050 553990
rect 124990 553930 125000 553970
rect 125040 553930 125050 553970
rect 119510 553860 119610 553880
rect 124990 553800 125050 553930
rect 125090 553970 125170 553990
rect 125090 553930 125110 553970
rect 125150 553930 125170 553970
rect 125090 553910 125170 553930
rect 125210 553970 125270 553990
rect 125210 553930 125220 553970
rect 125260 553930 125270 553970
rect 125210 553800 125270 553930
rect 311942 553908 312038 554900
rect 370968 554452 371064 555444
rect 370436 554356 371064 554452
rect 311942 553812 312200 553908
rect 119940 553440 120040 553460
rect 120310 553440 120410 553450
rect 119940 553380 119960 553440
rect 120020 553430 120410 553440
rect 120020 553380 120330 553430
rect 119940 553360 120040 553380
rect 120310 553370 120330 553380
rect 120390 553370 120410 553430
rect 120310 553350 120410 553370
rect 119350 553300 119370 553350
rect 119410 553300 119450 553350
rect 119350 552920 119450 553300
rect 119700 553280 119800 553290
rect 119700 553200 119710 553280
rect 119790 553200 119800 553280
rect 119700 553190 119800 553200
rect 119940 553270 124402 553290
rect 119940 553210 119960 553270
rect 120020 553210 124402 553270
rect 119940 553190 124402 553210
rect 119350 552860 119370 552920
rect 119430 552860 119450 552920
rect 119350 552850 119450 552860
rect 124302 552484 124402 553190
rect 311942 552820 312038 553812
rect 370968 553364 371064 554356
rect 370436 553268 371064 553364
rect 311942 552724 312200 552820
rect 124302 552420 133728 552484
rect 124302 552384 125750 552420
rect 125740 552380 125750 552384
rect 125790 552384 126190 552420
rect 125790 552380 125800 552384
rect 125740 552360 125800 552380
rect 126180 552380 126190 552384
rect 126230 552384 126630 552420
rect 126230 552380 126240 552384
rect 126180 552360 126240 552380
rect 126620 552380 126630 552384
rect 126670 552384 127070 552420
rect 126670 552380 126680 552384
rect 126620 552360 126680 552380
rect 127060 552380 127070 552384
rect 127110 552384 127510 552420
rect 127110 552380 127120 552384
rect 127060 552360 127120 552380
rect 127500 552380 127510 552384
rect 127550 552384 127950 552420
rect 127550 552380 127560 552384
rect 127500 552360 127560 552380
rect 127940 552380 127950 552384
rect 127990 552384 128390 552420
rect 127990 552380 128000 552384
rect 127940 552360 128000 552380
rect 128380 552380 128390 552384
rect 128430 552384 128830 552420
rect 128430 552380 128440 552384
rect 128380 552360 128440 552380
rect 128820 552380 128830 552384
rect 128870 552384 129270 552420
rect 128870 552380 128880 552384
rect 128820 552360 128880 552380
rect 129260 552380 129270 552384
rect 129310 552384 129710 552420
rect 129310 552380 129320 552384
rect 129260 552360 129320 552380
rect 129700 552380 129710 552384
rect 129750 552384 130150 552420
rect 129750 552380 129760 552384
rect 129700 552360 129760 552380
rect 130140 552380 130150 552384
rect 130190 552384 130590 552420
rect 130190 552380 130200 552384
rect 130140 552360 130200 552380
rect 130580 552380 130590 552384
rect 130630 552384 131030 552420
rect 130630 552380 130640 552384
rect 130580 552360 130640 552380
rect 131020 552380 131030 552384
rect 131070 552384 131470 552420
rect 131070 552380 131080 552384
rect 131020 552360 131080 552380
rect 131460 552380 131470 552384
rect 131510 552384 131910 552420
rect 131510 552380 131520 552384
rect 131460 552360 131520 552380
rect 131900 552380 131910 552384
rect 131950 552384 132350 552420
rect 131950 552380 131960 552384
rect 131900 552360 131960 552380
rect 132340 552380 132350 552384
rect 132390 552384 132790 552420
rect 132390 552380 132400 552384
rect 132340 552360 132400 552380
rect 132780 552380 132790 552384
rect 132830 552384 133230 552420
rect 132830 552380 132840 552384
rect 132780 552360 132840 552380
rect 133220 552380 133230 552384
rect 133270 552384 133670 552420
rect 133270 552380 133280 552384
rect 133220 552360 133280 552380
rect 133660 552380 133670 552384
rect 133710 552384 133728 552420
rect 133870 552460 134060 552480
rect 133710 552380 133720 552384
rect 133660 552360 133720 552380
rect 125420 552270 128830 552330
rect 129380 552270 133780 552330
rect 125590 552240 125750 552270
rect 126030 552240 126190 552270
rect 126470 552240 126630 552270
rect 126910 552240 127070 552270
rect 127350 552240 127510 552270
rect 127790 552240 127950 552270
rect 128230 552240 128390 552270
rect 128670 552240 128830 552270
rect 129110 552240 129270 552270
rect 129550 552240 129710 552270
rect 129990 552240 130150 552270
rect 130430 552240 130590 552270
rect 130870 552240 131030 552270
rect 131310 552240 131470 552270
rect 131750 552240 131910 552270
rect 132190 552240 132350 552270
rect 132630 552240 132790 552270
rect 133070 552240 133230 552270
rect 133510 552240 133670 552270
rect 125480 552220 125540 552240
rect 125480 552180 125490 552220
rect 125530 552180 125540 552220
rect 125480 552110 125540 552180
rect 125580 552220 125760 552240
rect 125580 552180 125600 552220
rect 125740 552180 125760 552220
rect 125580 552160 125760 552180
rect 125800 552220 125860 552240
rect 125800 552180 125810 552220
rect 125850 552180 125860 552220
rect 125800 552110 125860 552180
rect 125920 552220 125980 552240
rect 125920 552180 125930 552220
rect 125970 552180 125980 552220
rect 125920 552110 125980 552180
rect 126020 552220 126200 552240
rect 126020 552180 126040 552220
rect 126180 552180 126200 552220
rect 126020 552160 126200 552180
rect 126240 552220 126300 552240
rect 126240 552180 126250 552220
rect 126290 552180 126300 552220
rect 126240 552110 126300 552180
rect 126360 552220 126420 552240
rect 126360 552180 126370 552220
rect 126410 552180 126420 552220
rect 126360 552110 126420 552180
rect 126460 552220 126640 552240
rect 126460 552180 126480 552220
rect 126620 552180 126640 552220
rect 126460 552160 126640 552180
rect 126680 552220 126740 552240
rect 126680 552180 126690 552220
rect 126730 552180 126740 552220
rect 126680 552110 126740 552180
rect 126800 552220 126860 552240
rect 126800 552180 126810 552220
rect 126850 552180 126860 552220
rect 126800 552110 126860 552180
rect 126900 552220 127080 552240
rect 126900 552180 126920 552220
rect 127060 552180 127080 552220
rect 126900 552160 127080 552180
rect 127120 552220 127180 552240
rect 127120 552180 127130 552220
rect 127170 552180 127180 552220
rect 127120 552110 127180 552180
rect 127240 552220 127300 552240
rect 127240 552180 127250 552220
rect 127290 552180 127300 552220
rect 127240 552110 127300 552180
rect 127340 552220 127520 552240
rect 127340 552180 127360 552220
rect 127500 552180 127520 552220
rect 127340 552160 127520 552180
rect 127560 552220 127620 552240
rect 127560 552180 127570 552220
rect 127610 552180 127620 552220
rect 127560 552110 127620 552180
rect 127680 552220 127740 552240
rect 127680 552180 127690 552220
rect 127730 552180 127740 552220
rect 127680 552110 127740 552180
rect 127780 552220 127960 552240
rect 127780 552180 127800 552220
rect 127940 552180 127960 552220
rect 127780 552160 127960 552180
rect 128000 552220 128060 552240
rect 128000 552180 128010 552220
rect 128050 552180 128060 552220
rect 128000 552110 128060 552180
rect 128120 552220 128180 552240
rect 128120 552180 128130 552220
rect 128170 552180 128180 552220
rect 128120 552110 128180 552180
rect 128220 552220 128400 552240
rect 128220 552180 128240 552220
rect 128380 552180 128400 552220
rect 128220 552160 128400 552180
rect 128440 552220 128500 552240
rect 128440 552180 128450 552220
rect 128490 552180 128500 552220
rect 128440 552110 128500 552180
rect 128560 552220 128620 552240
rect 128560 552180 128570 552220
rect 128610 552180 128620 552220
rect 128560 552110 128620 552180
rect 128660 552220 128840 552240
rect 128660 552180 128680 552220
rect 128820 552180 128840 552220
rect 128660 552160 128840 552180
rect 128880 552220 128940 552240
rect 128880 552180 128890 552220
rect 128930 552180 128940 552220
rect 128880 552110 128940 552180
rect 129000 552220 129060 552240
rect 129000 552180 129010 552220
rect 129050 552180 129060 552220
rect 129000 552110 129060 552180
rect 129100 552220 129280 552240
rect 129100 552180 129120 552220
rect 129260 552180 129280 552220
rect 129100 552160 129280 552180
rect 129320 552220 129380 552240
rect 129320 552180 129330 552220
rect 129370 552180 129380 552220
rect 129320 552110 129380 552180
rect 129440 552220 129500 552240
rect 129440 552180 129450 552220
rect 129490 552180 129500 552220
rect 129440 552110 129500 552180
rect 129540 552220 129720 552240
rect 129540 552180 129560 552220
rect 129700 552180 129720 552220
rect 129540 552160 129720 552180
rect 129760 552220 129820 552240
rect 129760 552180 129770 552220
rect 129810 552180 129820 552220
rect 129760 552110 129820 552180
rect 129880 552220 129940 552240
rect 129880 552180 129890 552220
rect 129930 552180 129940 552220
rect 129880 552110 129940 552180
rect 129980 552220 130160 552240
rect 129980 552180 130000 552220
rect 130140 552180 130160 552220
rect 129980 552160 130160 552180
rect 130200 552220 130260 552240
rect 130200 552180 130210 552220
rect 130250 552180 130260 552220
rect 130200 552110 130260 552180
rect 130320 552220 130380 552240
rect 130320 552180 130330 552220
rect 130370 552180 130380 552220
rect 130320 552110 130380 552180
rect 130420 552220 130600 552240
rect 130420 552180 130440 552220
rect 130580 552180 130600 552220
rect 130420 552160 130600 552180
rect 130640 552220 130700 552240
rect 130640 552180 130650 552220
rect 130690 552180 130700 552220
rect 130640 552110 130700 552180
rect 130760 552220 130820 552240
rect 130760 552180 130770 552220
rect 130810 552180 130820 552220
rect 130760 552110 130820 552180
rect 130860 552220 131040 552240
rect 130860 552180 130880 552220
rect 131020 552180 131040 552220
rect 130860 552160 131040 552180
rect 131080 552220 131140 552240
rect 131080 552180 131090 552220
rect 131130 552180 131140 552220
rect 131080 552110 131140 552180
rect 131200 552220 131260 552240
rect 131200 552180 131210 552220
rect 131250 552180 131260 552220
rect 131200 552110 131260 552180
rect 131300 552220 131480 552240
rect 131300 552180 131320 552220
rect 131460 552180 131480 552220
rect 131300 552160 131480 552180
rect 131520 552220 131580 552240
rect 131520 552180 131530 552220
rect 131570 552180 131580 552220
rect 131520 552110 131580 552180
rect 131640 552220 131700 552240
rect 131640 552180 131650 552220
rect 131690 552180 131700 552220
rect 131640 552110 131700 552180
rect 131740 552220 131920 552240
rect 131740 552180 131760 552220
rect 131900 552180 131920 552220
rect 131740 552160 131920 552180
rect 131960 552220 132020 552240
rect 131960 552180 131970 552220
rect 132010 552180 132020 552220
rect 131960 552110 132020 552180
rect 132080 552220 132140 552240
rect 132080 552180 132090 552220
rect 132130 552180 132140 552220
rect 132080 552110 132140 552180
rect 132180 552220 132360 552240
rect 132180 552180 132200 552220
rect 132340 552180 132360 552220
rect 132180 552160 132360 552180
rect 132400 552220 132460 552240
rect 132400 552180 132410 552220
rect 132450 552180 132460 552220
rect 132400 552110 132460 552180
rect 132520 552220 132580 552240
rect 132520 552180 132530 552220
rect 132570 552180 132580 552220
rect 132520 552110 132580 552180
rect 132620 552220 132800 552240
rect 132620 552180 132640 552220
rect 132780 552180 132800 552220
rect 132620 552160 132800 552180
rect 132840 552220 132900 552240
rect 132840 552180 132850 552220
rect 132890 552180 132900 552220
rect 132840 552110 132900 552180
rect 132960 552220 133020 552240
rect 132960 552180 132970 552220
rect 133010 552180 133020 552220
rect 132960 552110 133020 552180
rect 133060 552220 133240 552240
rect 133060 552180 133080 552220
rect 133220 552180 133240 552220
rect 133060 552160 133240 552180
rect 133280 552220 133340 552240
rect 133280 552180 133290 552220
rect 133330 552180 133340 552220
rect 133280 552110 133340 552180
rect 133400 552220 133460 552240
rect 133400 552180 133410 552220
rect 133450 552180 133460 552220
rect 133400 552110 133460 552180
rect 133500 552220 133680 552240
rect 133500 552180 133520 552220
rect 133660 552180 133680 552220
rect 133500 552160 133680 552180
rect 133720 552220 133780 552240
rect 133720 552180 133730 552220
rect 133770 552180 133780 552220
rect 133720 552110 133780 552180
rect 125480 552050 128830 552110
rect 129380 552050 133780 552110
rect 133870 551890 133900 552460
rect 134030 551890 134060 552460
rect 133870 551870 134060 551890
rect 311942 551732 312038 552724
rect 370968 552276 371064 553268
rect 370436 552180 371064 552276
rect 311942 551636 312200 551732
rect 311942 550644 312038 551636
rect 370968 551188 371064 552180
rect 370436 551092 371064 551188
rect 311942 550548 312200 550644
rect 311942 549556 312038 550548
rect 370968 550100 371064 551092
rect 370436 550004 371064 550100
rect 311942 549460 312200 549556
rect 311942 548468 312038 549460
rect 370968 549012 371064 550004
rect 370436 548916 371064 549012
rect 311942 548372 312200 548468
rect 311942 547380 312038 548372
rect 370968 547924 371064 548916
rect 370436 547828 371064 547924
rect 311942 547284 312200 547380
rect 119350 547028 119450 547058
rect 119330 547022 119450 547028
rect 119330 546942 119336 547022
rect 119428 546942 119450 547022
rect 119330 546904 119450 546942
rect 119120 546492 119220 546500
rect 119120 546408 119128 546492
rect 119210 546490 119220 546492
rect 119210 546408 119290 546490
rect 119120 546394 119290 546408
rect 119190 546260 119290 546394
rect 119190 546200 119210 546260
rect 119270 546200 119290 546260
rect 119190 546180 119290 546200
rect 119350 545780 119450 546904
rect 119510 546448 120268 546490
rect 124940 546450 125360 546510
rect 119510 546390 120170 546448
rect 119510 546370 119610 546390
rect 119510 546310 119530 546370
rect 119590 546310 119610 546370
rect 120164 546368 120170 546390
rect 120262 546390 120268 546448
rect 125100 546420 125160 546450
rect 124990 546400 125050 546420
rect 120262 546368 120264 546390
rect 120164 546330 120264 546368
rect 124990 546360 125000 546400
rect 125040 546360 125050 546400
rect 119510 546290 119610 546310
rect 124990 546230 125050 546360
rect 125090 546400 125170 546420
rect 125090 546360 125110 546400
rect 125150 546360 125170 546400
rect 125090 546340 125170 546360
rect 125210 546400 125270 546420
rect 125210 546360 125220 546400
rect 125260 546360 125270 546400
rect 125210 546230 125270 546360
rect 311942 546292 312038 547284
rect 370968 546836 371064 547828
rect 370436 546740 371064 546836
rect 311942 546196 312200 546292
rect 119940 545870 120040 545890
rect 120310 545870 120410 545880
rect 119940 545810 119960 545870
rect 120020 545860 120410 545870
rect 120020 545810 120330 545860
rect 119940 545790 120040 545810
rect 120310 545800 120330 545810
rect 120390 545800 120410 545860
rect 120310 545780 120410 545800
rect 119350 545730 119370 545780
rect 119410 545730 119450 545780
rect 119350 545350 119450 545730
rect 119700 545710 119800 545720
rect 119700 545630 119710 545710
rect 119790 545630 119800 545710
rect 119700 545620 119800 545630
rect 119940 545700 124402 545720
rect 119940 545640 119960 545700
rect 120020 545640 124402 545700
rect 119940 545620 124402 545640
rect 119350 545290 119370 545350
rect 119430 545290 119450 545350
rect 119350 545280 119450 545290
rect 124302 544914 124402 545620
rect 311942 545204 312038 546196
rect 370968 545748 371064 546740
rect 370436 545652 371064 545748
rect 311942 545108 312200 545204
rect 124302 544850 133728 544914
rect 124302 544814 125750 544850
rect 125740 544810 125750 544814
rect 125790 544814 126190 544850
rect 125790 544810 125800 544814
rect 125740 544790 125800 544810
rect 126180 544810 126190 544814
rect 126230 544814 126630 544850
rect 126230 544810 126240 544814
rect 126180 544790 126240 544810
rect 126620 544810 126630 544814
rect 126670 544814 127070 544850
rect 126670 544810 126680 544814
rect 126620 544790 126680 544810
rect 127060 544810 127070 544814
rect 127110 544814 127510 544850
rect 127110 544810 127120 544814
rect 127060 544790 127120 544810
rect 127500 544810 127510 544814
rect 127550 544814 127950 544850
rect 127550 544810 127560 544814
rect 127500 544790 127560 544810
rect 127940 544810 127950 544814
rect 127990 544814 128390 544850
rect 127990 544810 128000 544814
rect 127940 544790 128000 544810
rect 128380 544810 128390 544814
rect 128430 544814 128830 544850
rect 128430 544810 128440 544814
rect 128380 544790 128440 544810
rect 128820 544810 128830 544814
rect 128870 544814 129270 544850
rect 128870 544810 128880 544814
rect 128820 544790 128880 544810
rect 129260 544810 129270 544814
rect 129310 544814 129710 544850
rect 129310 544810 129320 544814
rect 129260 544790 129320 544810
rect 129700 544810 129710 544814
rect 129750 544814 130150 544850
rect 129750 544810 129760 544814
rect 129700 544790 129760 544810
rect 130140 544810 130150 544814
rect 130190 544814 130590 544850
rect 130190 544810 130200 544814
rect 130140 544790 130200 544810
rect 130580 544810 130590 544814
rect 130630 544814 131030 544850
rect 130630 544810 130640 544814
rect 130580 544790 130640 544810
rect 131020 544810 131030 544814
rect 131070 544814 131470 544850
rect 131070 544810 131080 544814
rect 131020 544790 131080 544810
rect 131460 544810 131470 544814
rect 131510 544814 131910 544850
rect 131510 544810 131520 544814
rect 131460 544790 131520 544810
rect 131900 544810 131910 544814
rect 131950 544814 132350 544850
rect 131950 544810 131960 544814
rect 131900 544790 131960 544810
rect 132340 544810 132350 544814
rect 132390 544814 132790 544850
rect 132390 544810 132400 544814
rect 132340 544790 132400 544810
rect 132780 544810 132790 544814
rect 132830 544814 133230 544850
rect 132830 544810 132840 544814
rect 132780 544790 132840 544810
rect 133220 544810 133230 544814
rect 133270 544814 133670 544850
rect 133270 544810 133280 544814
rect 133220 544790 133280 544810
rect 133660 544810 133670 544814
rect 133710 544814 133728 544850
rect 133870 544890 134060 544910
rect 133710 544810 133720 544814
rect 133660 544790 133720 544810
rect 125420 544700 128830 544760
rect 129380 544700 133780 544760
rect 125590 544670 125750 544700
rect 126030 544670 126190 544700
rect 126470 544670 126630 544700
rect 126910 544670 127070 544700
rect 127350 544670 127510 544700
rect 127790 544670 127950 544700
rect 128230 544670 128390 544700
rect 128670 544670 128830 544700
rect 129110 544670 129270 544700
rect 129550 544670 129710 544700
rect 129990 544670 130150 544700
rect 130430 544670 130590 544700
rect 130870 544670 131030 544700
rect 131310 544670 131470 544700
rect 131750 544670 131910 544700
rect 132190 544670 132350 544700
rect 132630 544670 132790 544700
rect 133070 544670 133230 544700
rect 133510 544670 133670 544700
rect 125480 544650 125540 544670
rect 125480 544410 125490 544650
rect 125530 544410 125540 544650
rect 125480 544340 125540 544410
rect 125580 544650 125760 544670
rect 125580 544410 125600 544650
rect 125740 544410 125760 544650
rect 125580 544390 125760 544410
rect 125800 544650 125860 544670
rect 125800 544410 125810 544650
rect 125850 544410 125860 544650
rect 125800 544340 125860 544410
rect 125920 544650 125980 544670
rect 125920 544410 125930 544650
rect 125970 544410 125980 544650
rect 125920 544340 125980 544410
rect 126020 544650 126200 544670
rect 126020 544410 126040 544650
rect 126180 544410 126200 544650
rect 126020 544390 126200 544410
rect 126240 544650 126300 544670
rect 126240 544410 126250 544650
rect 126290 544410 126300 544650
rect 126240 544340 126300 544410
rect 126360 544650 126420 544670
rect 126360 544410 126370 544650
rect 126410 544410 126420 544650
rect 126360 544340 126420 544410
rect 126460 544650 126640 544670
rect 126460 544410 126480 544650
rect 126620 544410 126640 544650
rect 126460 544390 126640 544410
rect 126680 544650 126740 544670
rect 126680 544410 126690 544650
rect 126730 544410 126740 544650
rect 126680 544340 126740 544410
rect 126800 544650 126860 544670
rect 126800 544410 126810 544650
rect 126850 544410 126860 544650
rect 126800 544340 126860 544410
rect 126900 544650 127080 544670
rect 126900 544410 126920 544650
rect 127060 544410 127080 544650
rect 126900 544390 127080 544410
rect 127120 544650 127180 544670
rect 127120 544410 127130 544650
rect 127170 544410 127180 544650
rect 127120 544340 127180 544410
rect 127240 544650 127300 544670
rect 127240 544410 127250 544650
rect 127290 544410 127300 544650
rect 127240 544340 127300 544410
rect 127340 544650 127520 544670
rect 127340 544410 127360 544650
rect 127500 544410 127520 544650
rect 127340 544390 127520 544410
rect 127560 544650 127620 544670
rect 127560 544410 127570 544650
rect 127610 544410 127620 544650
rect 127560 544340 127620 544410
rect 127680 544650 127740 544670
rect 127680 544410 127690 544650
rect 127730 544410 127740 544650
rect 127680 544340 127740 544410
rect 127780 544650 127960 544670
rect 127780 544410 127800 544650
rect 127940 544410 127960 544650
rect 127780 544390 127960 544410
rect 128000 544650 128060 544670
rect 128000 544410 128010 544650
rect 128050 544410 128060 544650
rect 128000 544340 128060 544410
rect 128120 544650 128180 544670
rect 128120 544410 128130 544650
rect 128170 544410 128180 544650
rect 128120 544340 128180 544410
rect 128220 544650 128400 544670
rect 128220 544410 128240 544650
rect 128380 544410 128400 544650
rect 128220 544390 128400 544410
rect 128440 544650 128500 544670
rect 128440 544410 128450 544650
rect 128490 544410 128500 544650
rect 128440 544340 128500 544410
rect 128560 544650 128620 544670
rect 128560 544410 128570 544650
rect 128610 544410 128620 544650
rect 128560 544340 128620 544410
rect 128660 544650 128840 544670
rect 128660 544410 128680 544650
rect 128820 544410 128840 544650
rect 128660 544390 128840 544410
rect 128880 544650 128940 544670
rect 128880 544410 128890 544650
rect 128930 544410 128940 544650
rect 128880 544340 128940 544410
rect 129000 544650 129060 544670
rect 129000 544410 129010 544650
rect 129050 544410 129060 544650
rect 129000 544340 129060 544410
rect 129100 544650 129280 544670
rect 129100 544410 129120 544650
rect 129260 544410 129280 544650
rect 129100 544390 129280 544410
rect 129320 544650 129380 544670
rect 129320 544410 129330 544650
rect 129370 544410 129380 544650
rect 129320 544340 129380 544410
rect 129440 544650 129500 544670
rect 129440 544410 129450 544650
rect 129490 544410 129500 544650
rect 129440 544340 129500 544410
rect 129540 544650 129720 544670
rect 129540 544410 129560 544650
rect 129700 544410 129720 544650
rect 129540 544390 129720 544410
rect 129760 544650 129820 544670
rect 129760 544410 129770 544650
rect 129810 544410 129820 544650
rect 129760 544340 129820 544410
rect 129880 544650 129940 544670
rect 129880 544410 129890 544650
rect 129930 544410 129940 544650
rect 129880 544340 129940 544410
rect 129980 544650 130160 544670
rect 129980 544410 130000 544650
rect 130140 544410 130160 544650
rect 129980 544390 130160 544410
rect 130200 544650 130260 544670
rect 130200 544410 130210 544650
rect 130250 544410 130260 544650
rect 130200 544340 130260 544410
rect 130320 544650 130380 544670
rect 130320 544410 130330 544650
rect 130370 544410 130380 544650
rect 130320 544340 130380 544410
rect 130420 544650 130600 544670
rect 130420 544410 130440 544650
rect 130580 544410 130600 544650
rect 130420 544390 130600 544410
rect 130640 544650 130700 544670
rect 130640 544410 130650 544650
rect 130690 544410 130700 544650
rect 130640 544340 130700 544410
rect 130760 544650 130820 544670
rect 130760 544410 130770 544650
rect 130810 544410 130820 544650
rect 130760 544340 130820 544410
rect 130860 544650 131040 544670
rect 130860 544410 130880 544650
rect 131020 544410 131040 544650
rect 130860 544390 131040 544410
rect 131080 544650 131140 544670
rect 131080 544410 131090 544650
rect 131130 544410 131140 544650
rect 131080 544340 131140 544410
rect 131200 544650 131260 544670
rect 131200 544410 131210 544650
rect 131250 544410 131260 544650
rect 131200 544340 131260 544410
rect 131300 544650 131480 544670
rect 131300 544410 131320 544650
rect 131460 544410 131480 544650
rect 131300 544390 131480 544410
rect 131520 544650 131580 544670
rect 131520 544410 131530 544650
rect 131570 544410 131580 544650
rect 131520 544340 131580 544410
rect 131640 544650 131700 544670
rect 131640 544410 131650 544650
rect 131690 544410 131700 544650
rect 131640 544340 131700 544410
rect 131740 544650 131920 544670
rect 131740 544410 131760 544650
rect 131900 544410 131920 544650
rect 131740 544390 131920 544410
rect 131960 544650 132020 544670
rect 131960 544410 131970 544650
rect 132010 544410 132020 544650
rect 131960 544340 132020 544410
rect 132080 544650 132140 544670
rect 132080 544410 132090 544650
rect 132130 544410 132140 544650
rect 132080 544340 132140 544410
rect 132180 544650 132360 544670
rect 132180 544410 132200 544650
rect 132340 544410 132360 544650
rect 132180 544390 132360 544410
rect 132400 544650 132460 544670
rect 132400 544410 132410 544650
rect 132450 544410 132460 544650
rect 132400 544340 132460 544410
rect 132520 544650 132580 544670
rect 132520 544410 132530 544650
rect 132570 544410 132580 544650
rect 132520 544340 132580 544410
rect 132620 544650 132800 544670
rect 132620 544410 132640 544650
rect 132780 544410 132800 544650
rect 132620 544390 132800 544410
rect 132840 544650 132900 544670
rect 132840 544410 132850 544650
rect 132890 544410 132900 544650
rect 132840 544340 132900 544410
rect 132960 544650 133020 544670
rect 132960 544410 132970 544650
rect 133010 544410 133020 544650
rect 132960 544340 133020 544410
rect 133060 544650 133240 544670
rect 133060 544410 133080 544650
rect 133220 544410 133240 544650
rect 133060 544390 133240 544410
rect 133280 544650 133340 544670
rect 133280 544410 133290 544650
rect 133330 544410 133340 544650
rect 133280 544340 133340 544410
rect 133400 544650 133460 544670
rect 133400 544410 133410 544650
rect 133450 544410 133460 544650
rect 133400 544340 133460 544410
rect 133500 544650 133680 544670
rect 133500 544410 133520 544650
rect 133660 544410 133680 544650
rect 133500 544390 133680 544410
rect 133720 544650 133780 544670
rect 133720 544410 133730 544650
rect 133770 544410 133780 544650
rect 133720 544340 133780 544410
rect 125480 544280 128830 544340
rect 129380 544280 133780 544340
rect 133870 544120 133900 544890
rect 134030 544120 134060 544890
rect 133870 544100 134060 544120
rect 311942 544116 312038 545108
rect 370968 544660 371064 545652
rect 370436 544564 371064 544660
rect 311942 544020 312200 544116
rect 311942 543028 312038 544020
rect 370968 543572 371064 544564
rect 370436 543476 371064 543572
rect 311942 542932 312200 543028
rect 311942 541940 312038 542932
rect 370968 542484 371064 543476
rect 370436 542388 371064 542484
rect 311942 541844 312200 541940
rect 311942 540852 312038 541844
rect 370968 541396 371064 542388
rect 370436 541300 371064 541396
rect 311942 540756 312200 540852
rect 311942 539764 312038 540756
rect 370968 540308 371064 541300
rect 370436 540212 371064 540308
rect 311942 539668 312200 539764
rect 119312 538982 119412 538988
rect 119312 538902 119318 538982
rect 119410 538940 119412 538982
rect 119410 538902 119420 538940
rect 119312 538864 119420 538902
rect 119124 538474 119224 538482
rect 119124 538390 119132 538474
rect 119214 538430 119224 538474
rect 119214 538390 119260 538430
rect 119124 538376 119260 538390
rect 119160 538200 119260 538376
rect 119160 538140 119180 538200
rect 119240 538140 119260 538200
rect 119160 538120 119260 538140
rect 119320 537720 119420 538864
rect 311942 538676 312038 539668
rect 370968 539220 371064 540212
rect 370436 539124 371064 539220
rect 311942 538580 312200 538676
rect 119480 538424 120140 538430
rect 119480 538344 120046 538424
rect 120138 538344 120140 538424
rect 124910 538390 125330 538450
rect 125070 538360 125130 538390
rect 119480 538330 120140 538344
rect 119480 538310 119580 538330
rect 119480 538250 119500 538310
rect 119560 538250 119580 538310
rect 120040 538306 120140 538330
rect 124960 538340 125020 538360
rect 119480 538230 119580 538250
rect 124960 538300 124970 538340
rect 125010 538300 125020 538340
rect 124960 538170 125020 538300
rect 125060 538340 125140 538360
rect 125060 538300 125080 538340
rect 125120 538300 125140 538340
rect 125060 538280 125140 538300
rect 125180 538340 125240 538360
rect 125180 538300 125190 538340
rect 125230 538300 125240 538340
rect 125180 538170 125240 538300
rect 119910 537810 120010 537830
rect 120280 537810 120380 537820
rect 119910 537750 119930 537810
rect 119990 537800 120380 537810
rect 119990 537750 120300 537800
rect 119910 537730 120010 537750
rect 120280 537740 120300 537750
rect 120360 537740 120380 537800
rect 120280 537720 120380 537740
rect 119320 537670 119340 537720
rect 119380 537670 119420 537720
rect 119320 537290 119420 537670
rect 119670 537650 119770 537660
rect 119670 537570 119680 537650
rect 119760 537570 119770 537650
rect 119670 537560 119770 537570
rect 119910 537640 124372 537660
rect 119910 537580 119930 537640
rect 119990 537580 124372 537640
rect 119910 537560 124372 537580
rect 119320 537230 119340 537290
rect 119400 537230 119420 537290
rect 119320 537220 119420 537230
rect 124272 536854 124372 537560
rect 311942 537588 312038 538580
rect 370968 538132 371064 539124
rect 370436 538036 371064 538132
rect 311942 537492 312200 537588
rect 124272 536790 133698 536854
rect 124272 536754 125720 536790
rect 125710 536750 125720 536754
rect 125760 536754 126160 536790
rect 125760 536750 125770 536754
rect 125710 536730 125770 536750
rect 126150 536750 126160 536754
rect 126200 536754 126600 536790
rect 126200 536750 126210 536754
rect 126150 536730 126210 536750
rect 126590 536750 126600 536754
rect 126640 536754 127040 536790
rect 126640 536750 126650 536754
rect 126590 536730 126650 536750
rect 127030 536750 127040 536754
rect 127080 536754 127480 536790
rect 127080 536750 127090 536754
rect 127030 536730 127090 536750
rect 127470 536750 127480 536754
rect 127520 536754 127920 536790
rect 127520 536750 127530 536754
rect 127470 536730 127530 536750
rect 127910 536750 127920 536754
rect 127960 536754 128360 536790
rect 127960 536750 127970 536754
rect 127910 536730 127970 536750
rect 128350 536750 128360 536754
rect 128400 536754 128800 536790
rect 128400 536750 128410 536754
rect 128350 536730 128410 536750
rect 128790 536750 128800 536754
rect 128840 536754 129240 536790
rect 128840 536750 128850 536754
rect 128790 536730 128850 536750
rect 129230 536750 129240 536754
rect 129280 536754 129680 536790
rect 129280 536750 129290 536754
rect 129230 536730 129290 536750
rect 129670 536750 129680 536754
rect 129720 536754 130120 536790
rect 129720 536750 129730 536754
rect 129670 536730 129730 536750
rect 130110 536750 130120 536754
rect 130160 536754 130560 536790
rect 130160 536750 130170 536754
rect 130110 536730 130170 536750
rect 130550 536750 130560 536754
rect 130600 536754 131000 536790
rect 130600 536750 130610 536754
rect 130550 536730 130610 536750
rect 130990 536750 131000 536754
rect 131040 536754 131440 536790
rect 131040 536750 131050 536754
rect 130990 536730 131050 536750
rect 131430 536750 131440 536754
rect 131480 536754 131880 536790
rect 131480 536750 131490 536754
rect 131430 536730 131490 536750
rect 131870 536750 131880 536754
rect 131920 536754 132320 536790
rect 131920 536750 131930 536754
rect 131870 536730 131930 536750
rect 132310 536750 132320 536754
rect 132360 536754 132760 536790
rect 132360 536750 132370 536754
rect 132310 536730 132370 536750
rect 132750 536750 132760 536754
rect 132800 536754 133200 536790
rect 132800 536750 132810 536754
rect 132750 536730 132810 536750
rect 133190 536750 133200 536754
rect 133240 536754 133640 536790
rect 133240 536750 133250 536754
rect 133190 536730 133250 536750
rect 133630 536750 133640 536754
rect 133680 536754 133698 536790
rect 133840 536830 134030 536850
rect 133680 536750 133690 536754
rect 133630 536730 133690 536750
rect 125390 536640 128800 536700
rect 129350 536640 133750 536700
rect 125560 536610 125720 536640
rect 126000 536610 126160 536640
rect 126440 536610 126600 536640
rect 126880 536610 127040 536640
rect 127320 536610 127480 536640
rect 127760 536610 127920 536640
rect 128200 536610 128360 536640
rect 128640 536610 128800 536640
rect 129080 536610 129240 536640
rect 129520 536610 129680 536640
rect 129960 536610 130120 536640
rect 130400 536610 130560 536640
rect 130840 536610 131000 536640
rect 131280 536610 131440 536640
rect 131720 536610 131880 536640
rect 132160 536610 132320 536640
rect 132600 536610 132760 536640
rect 133040 536610 133200 536640
rect 133480 536610 133640 536640
rect 125450 536590 125510 536610
rect 125450 536150 125460 536590
rect 125500 536150 125510 536590
rect 125450 536080 125510 536150
rect 125550 536590 125730 536610
rect 125550 536150 125570 536590
rect 125710 536150 125730 536590
rect 125550 536130 125730 536150
rect 125770 536590 125830 536610
rect 125770 536150 125780 536590
rect 125820 536150 125830 536590
rect 125770 536080 125830 536150
rect 125890 536590 125950 536610
rect 125890 536150 125900 536590
rect 125940 536150 125950 536590
rect 125890 536080 125950 536150
rect 125990 536590 126170 536610
rect 125990 536150 126010 536590
rect 126150 536150 126170 536590
rect 125990 536130 126170 536150
rect 126210 536590 126270 536610
rect 126210 536150 126220 536590
rect 126260 536150 126270 536590
rect 126210 536080 126270 536150
rect 126330 536590 126390 536610
rect 126330 536150 126340 536590
rect 126380 536150 126390 536590
rect 126330 536080 126390 536150
rect 126430 536590 126610 536610
rect 126430 536150 126450 536590
rect 126590 536150 126610 536590
rect 126430 536130 126610 536150
rect 126650 536590 126710 536610
rect 126650 536150 126660 536590
rect 126700 536150 126710 536590
rect 126650 536080 126710 536150
rect 126770 536590 126830 536610
rect 126770 536150 126780 536590
rect 126820 536150 126830 536590
rect 126770 536080 126830 536150
rect 126870 536590 127050 536610
rect 126870 536150 126890 536590
rect 127030 536150 127050 536590
rect 126870 536130 127050 536150
rect 127090 536590 127150 536610
rect 127090 536150 127100 536590
rect 127140 536150 127150 536590
rect 127090 536080 127150 536150
rect 127210 536590 127270 536610
rect 127210 536150 127220 536590
rect 127260 536150 127270 536590
rect 127210 536080 127270 536150
rect 127310 536590 127490 536610
rect 127310 536150 127330 536590
rect 127470 536150 127490 536590
rect 127310 536130 127490 536150
rect 127530 536590 127590 536610
rect 127530 536150 127540 536590
rect 127580 536150 127590 536590
rect 127530 536080 127590 536150
rect 127650 536590 127710 536610
rect 127650 536150 127660 536590
rect 127700 536150 127710 536590
rect 127650 536080 127710 536150
rect 127750 536590 127930 536610
rect 127750 536150 127770 536590
rect 127910 536150 127930 536590
rect 127750 536130 127930 536150
rect 127970 536590 128030 536610
rect 127970 536150 127980 536590
rect 128020 536150 128030 536590
rect 127970 536080 128030 536150
rect 128090 536590 128150 536610
rect 128090 536150 128100 536590
rect 128140 536150 128150 536590
rect 128090 536080 128150 536150
rect 128190 536590 128370 536610
rect 128190 536150 128210 536590
rect 128350 536150 128370 536590
rect 128190 536130 128370 536150
rect 128410 536590 128470 536610
rect 128410 536150 128420 536590
rect 128460 536150 128470 536590
rect 128410 536080 128470 536150
rect 128530 536590 128590 536610
rect 128530 536150 128540 536590
rect 128580 536150 128590 536590
rect 128530 536080 128590 536150
rect 128630 536590 128810 536610
rect 128630 536150 128650 536590
rect 128790 536150 128810 536590
rect 128630 536130 128810 536150
rect 128850 536590 128910 536610
rect 128850 536150 128860 536590
rect 128900 536150 128910 536590
rect 128850 536080 128910 536150
rect 128970 536590 129030 536610
rect 128970 536150 128980 536590
rect 129020 536150 129030 536590
rect 128970 536080 129030 536150
rect 129070 536590 129250 536610
rect 129070 536150 129090 536590
rect 129230 536150 129250 536590
rect 129070 536130 129250 536150
rect 129290 536590 129350 536610
rect 129290 536150 129300 536590
rect 129340 536150 129350 536590
rect 129290 536080 129350 536150
rect 129410 536590 129470 536610
rect 129410 536150 129420 536590
rect 129460 536150 129470 536590
rect 129410 536080 129470 536150
rect 129510 536590 129690 536610
rect 129510 536150 129530 536590
rect 129670 536150 129690 536590
rect 129510 536130 129690 536150
rect 129730 536590 129790 536610
rect 129730 536150 129740 536590
rect 129780 536150 129790 536590
rect 129730 536080 129790 536150
rect 129850 536590 129910 536610
rect 129850 536150 129860 536590
rect 129900 536150 129910 536590
rect 129850 536080 129910 536150
rect 129950 536590 130130 536610
rect 129950 536150 129970 536590
rect 130110 536150 130130 536590
rect 129950 536130 130130 536150
rect 130170 536590 130230 536610
rect 130170 536150 130180 536590
rect 130220 536150 130230 536590
rect 130170 536080 130230 536150
rect 130290 536590 130350 536610
rect 130290 536150 130300 536590
rect 130340 536150 130350 536590
rect 130290 536080 130350 536150
rect 130390 536590 130570 536610
rect 130390 536150 130410 536590
rect 130550 536150 130570 536590
rect 130390 536130 130570 536150
rect 130610 536590 130670 536610
rect 130610 536150 130620 536590
rect 130660 536150 130670 536590
rect 130610 536080 130670 536150
rect 130730 536590 130790 536610
rect 130730 536150 130740 536590
rect 130780 536150 130790 536590
rect 130730 536080 130790 536150
rect 130830 536590 131010 536610
rect 130830 536150 130850 536590
rect 130990 536150 131010 536590
rect 130830 536130 131010 536150
rect 131050 536590 131110 536610
rect 131050 536150 131060 536590
rect 131100 536150 131110 536590
rect 131050 536080 131110 536150
rect 131170 536590 131230 536610
rect 131170 536150 131180 536590
rect 131220 536150 131230 536590
rect 131170 536080 131230 536150
rect 131270 536590 131450 536610
rect 131270 536150 131290 536590
rect 131430 536150 131450 536590
rect 131270 536130 131450 536150
rect 131490 536590 131550 536610
rect 131490 536150 131500 536590
rect 131540 536150 131550 536590
rect 131490 536080 131550 536150
rect 131610 536590 131670 536610
rect 131610 536150 131620 536590
rect 131660 536150 131670 536590
rect 131610 536080 131670 536150
rect 131710 536590 131890 536610
rect 131710 536150 131730 536590
rect 131870 536150 131890 536590
rect 131710 536130 131890 536150
rect 131930 536590 131990 536610
rect 131930 536150 131940 536590
rect 131980 536150 131990 536590
rect 131930 536080 131990 536150
rect 132050 536590 132110 536610
rect 132050 536150 132060 536590
rect 132100 536150 132110 536590
rect 132050 536080 132110 536150
rect 132150 536590 132330 536610
rect 132150 536150 132170 536590
rect 132310 536150 132330 536590
rect 132150 536130 132330 536150
rect 132370 536590 132430 536610
rect 132370 536150 132380 536590
rect 132420 536150 132430 536590
rect 132370 536080 132430 536150
rect 132490 536590 132550 536610
rect 132490 536150 132500 536590
rect 132540 536150 132550 536590
rect 132490 536080 132550 536150
rect 132590 536590 132770 536610
rect 132590 536150 132610 536590
rect 132750 536150 132770 536590
rect 132590 536130 132770 536150
rect 132810 536590 132870 536610
rect 132810 536150 132820 536590
rect 132860 536150 132870 536590
rect 132810 536080 132870 536150
rect 132930 536590 132990 536610
rect 132930 536150 132940 536590
rect 132980 536150 132990 536590
rect 132930 536080 132990 536150
rect 133030 536590 133210 536610
rect 133030 536150 133050 536590
rect 133190 536150 133210 536590
rect 133030 536130 133210 536150
rect 133250 536590 133310 536610
rect 133250 536150 133260 536590
rect 133300 536150 133310 536590
rect 133250 536080 133310 536150
rect 133370 536590 133430 536610
rect 133370 536150 133380 536590
rect 133420 536150 133430 536590
rect 133370 536080 133430 536150
rect 133470 536590 133650 536610
rect 133470 536150 133490 536590
rect 133630 536150 133650 536590
rect 133470 536130 133650 536150
rect 133690 536590 133750 536610
rect 133690 536150 133700 536590
rect 133740 536150 133750 536590
rect 133690 536080 133750 536150
rect 125450 536020 128800 536080
rect 129350 536020 133750 536080
rect 133840 535860 133870 536830
rect 134000 535860 134030 536830
rect 133840 535840 134030 535860
rect 311942 536500 312038 537492
rect 370968 537044 371064 538036
rect 370436 536948 371064 537044
rect 311942 536404 312200 536500
rect 311942 535412 312038 536404
rect 370968 535956 371064 536948
rect 370436 535860 371064 535956
rect 311942 535316 312200 535412
rect 311942 534324 312038 535316
rect 370968 534868 371064 535860
rect 370436 534772 371064 534868
rect 311942 534228 312200 534324
rect 311942 533236 312038 534228
rect 370968 533780 371064 534772
rect 370436 533684 371064 533780
rect 311942 533140 312200 533236
rect 311942 532148 312038 533140
rect 370968 532692 371064 533684
rect 370436 532596 371064 532692
rect 311942 532052 312200 532148
rect 311942 531060 312038 532052
rect 370968 531604 371064 532596
rect 370436 531508 371064 531604
rect 311942 530977 312200 531060
rect 306149 530964 312200 530977
rect 370968 530977 371064 531508
rect 376448 560536 376544 561528
rect 437264 561524 437360 563752
rect 437264 561428 437520 561524
rect 435474 561392 435568 561420
rect 435216 561001 435568 561080
rect 435216 560984 435466 561001
rect 435460 560905 435466 560984
rect 435574 560905 435580 561001
rect 435474 560781 435568 560905
rect 376448 560440 377076 560536
rect 376448 559448 376544 560440
rect 435474 559992 435570 560781
rect 437264 560570 437358 561428
rect 495756 560977 496384 560980
rect 497075 560977 497171 563752
rect 500981 561624 501077 563752
rect 560792 561925 560888 563752
rect 560792 561817 560888 561829
rect 500981 561539 502492 561624
rect 500982 561528 502492 561539
rect 495756 560884 497171 560977
rect 435216 559896 435570 559992
rect 376448 559352 377076 559448
rect 376448 558360 376544 559352
rect 435474 558904 435570 559896
rect 435312 558808 435570 558904
rect 376448 558264 377076 558360
rect 376448 557272 376544 558264
rect 435474 557816 435570 558808
rect 435312 557720 435570 557816
rect 376448 557176 377076 557272
rect 376448 556184 376544 557176
rect 435474 556728 435570 557720
rect 435312 556632 435570 556728
rect 376448 556088 377076 556184
rect 376448 555096 376544 556088
rect 435474 555640 435570 556632
rect 435312 555544 435570 555640
rect 376448 555000 377076 555096
rect 376448 554008 376544 555000
rect 435474 554552 435570 555544
rect 435312 554456 435570 554552
rect 376448 553912 377076 554008
rect 376448 552920 376544 553912
rect 435474 553464 435570 554456
rect 435312 553368 435570 553464
rect 376448 552824 377076 552920
rect 376448 551832 376544 552824
rect 435474 552376 435570 553368
rect 435312 552280 435570 552376
rect 376448 551736 377076 551832
rect 376448 550744 376544 551736
rect 435474 551288 435570 552280
rect 435312 551192 435570 551288
rect 376448 550648 377076 550744
rect 376448 549656 376544 550648
rect 435474 550200 435570 551192
rect 435312 550104 435570 550200
rect 376448 549560 377076 549656
rect 376448 548568 376544 549560
rect 435474 549112 435570 550104
rect 435312 549016 435570 549112
rect 376448 548472 377076 548568
rect 376448 547480 376544 548472
rect 435474 548024 435570 549016
rect 435312 547928 435570 548024
rect 376448 547384 377076 547480
rect 376448 546392 376544 547384
rect 435474 546936 435570 547928
rect 435312 546840 435570 546936
rect 376448 546296 377076 546392
rect 376448 545304 376544 546296
rect 435474 545848 435570 546840
rect 435312 545752 435570 545848
rect 376448 545208 377076 545304
rect 376448 544216 376544 545208
rect 435474 544760 435570 545752
rect 435312 544664 435570 544760
rect 376448 544120 377076 544216
rect 376448 543128 376544 544120
rect 435474 543672 435570 544664
rect 435312 543576 435570 543672
rect 376448 543032 377076 543128
rect 376448 542040 376544 543032
rect 435474 542584 435570 543576
rect 435312 542488 435570 542584
rect 376448 541944 377076 542040
rect 376448 540952 376544 541944
rect 435474 541496 435570 542488
rect 435312 541400 435570 541496
rect 376448 540856 377076 540952
rect 376448 539864 376544 540856
rect 435474 540408 435570 541400
rect 435312 540312 435570 540408
rect 376448 539768 377076 539864
rect 376448 538776 376544 539768
rect 435474 539320 435570 540312
rect 435312 539224 435570 539320
rect 376448 538680 377076 538776
rect 376448 537688 376544 538680
rect 435474 538232 435570 539224
rect 435312 538136 435570 538232
rect 376448 537592 377076 537688
rect 376448 536600 376544 537592
rect 435474 537144 435570 538136
rect 435312 537048 435570 537144
rect 376448 536504 377076 536600
rect 376448 535512 376544 536504
rect 435474 536056 435570 537048
rect 435312 535960 435570 536056
rect 376448 535416 377076 535512
rect 376448 534424 376544 535416
rect 435474 534968 435570 535960
rect 435312 534872 435570 534968
rect 376448 534328 377076 534424
rect 376448 533336 376544 534328
rect 435474 533880 435570 534872
rect 435312 533784 435570 533880
rect 376448 533240 377076 533336
rect 376448 532248 376544 533240
rect 435474 532792 435570 533784
rect 435312 532696 435570 532792
rect 376448 532152 377076 532248
rect 376448 531160 376544 532152
rect 435474 531704 435570 532696
rect 435312 531608 435570 531704
rect 376448 531064 377076 531160
rect 376448 530977 376544 531064
rect 306149 530929 312038 530964
rect 306149 530001 307383 530929
rect 308407 530001 312038 530929
rect 370968 530929 376544 530977
rect 370968 530516 373176 530929
rect 370436 530420 373176 530516
rect 306149 529972 312038 530001
rect 370968 530001 373176 530420
rect 374200 530072 376544 530929
rect 435474 530616 435570 531608
rect 435312 530520 435570 530616
rect 374200 530001 377076 530072
rect 370968 529976 377076 530001
rect 306149 529953 312200 529972
rect 311942 529876 312200 529953
rect 370968 529953 376544 529976
rect 311942 528884 312038 529876
rect 370968 529428 371064 529953
rect 370436 529332 371064 529428
rect 311942 528788 312200 528884
rect 311942 527796 312038 528788
rect 370968 528340 371064 529332
rect 370436 528244 371064 528340
rect 311942 527700 312200 527796
rect 311942 526708 312038 527700
rect 370968 527252 371064 528244
rect 370436 527156 371064 527252
rect 311942 526612 312200 526708
rect 311942 525620 312038 526612
rect 370968 526164 371064 527156
rect 370436 526068 371064 526164
rect 311942 525524 312200 525620
rect 311942 524532 312038 525524
rect 370968 525076 371064 526068
rect 370436 524980 371064 525076
rect 311942 524436 312200 524532
rect 311942 523444 312038 524436
rect 370968 523988 371064 524980
rect 370436 523892 371064 523988
rect 311942 523348 312200 523444
rect 311942 522356 312038 523348
rect 370968 522900 371064 523892
rect 370436 522804 371064 522900
rect 311942 522260 312200 522356
rect 311942 521268 312038 522260
rect 370968 521812 371064 522804
rect 370436 521716 371064 521812
rect 311942 521172 312200 521268
rect 311942 520180 312038 521172
rect 370968 520724 371064 521716
rect 370436 520628 371064 520724
rect 311942 520084 312200 520180
rect 311942 519092 312038 520084
rect 370968 519636 371064 520628
rect 370436 519540 371064 519636
rect 311942 518996 312200 519092
rect 311942 518004 312038 518996
rect 370968 518548 371064 519540
rect 370436 518452 371064 518548
rect 311942 517908 312200 518004
rect 311942 516916 312038 517908
rect 370968 517460 371064 518452
rect 370436 517364 371064 517460
rect 311942 516820 312200 516916
rect 311942 515828 312038 516820
rect 370968 516372 371064 517364
rect 370436 516276 371064 516372
rect 311942 515732 312200 515828
rect 311942 514740 312038 515732
rect 370968 515284 371064 516276
rect 370436 515188 371064 515284
rect 311942 514644 312200 514740
rect 311942 513652 312038 514644
rect 370968 514196 371064 515188
rect 370436 514100 371064 514196
rect 311942 513556 312200 513652
rect 311942 512564 312038 513556
rect 370968 513108 371064 514100
rect 370436 513012 371064 513108
rect 311942 512468 312200 512564
rect 311942 511476 312038 512468
rect 370968 512020 371064 513012
rect 370436 511924 371064 512020
rect 311942 511380 312200 511476
rect 311942 510388 312038 511380
rect 370968 510932 371064 511924
rect 370436 510836 371064 510932
rect 311942 510292 312200 510388
rect 311942 509300 312038 510292
rect 370968 509844 371064 510836
rect 370436 509748 371064 509844
rect 311942 509204 312200 509300
rect 311942 508212 312038 509204
rect 370968 508756 371064 509748
rect 370436 508660 371064 508756
rect 311942 508116 312200 508212
rect 311942 507124 312038 508116
rect 370968 507668 371064 508660
rect 370436 507572 371064 507668
rect 311942 507028 312200 507124
rect 311942 506036 312038 507028
rect 370968 506580 371064 507572
rect 370436 506484 371064 506580
rect 311942 505940 312200 506036
rect 311942 504948 312038 505940
rect 370968 505492 371064 506484
rect 370436 505396 371064 505492
rect 311942 504852 312296 504948
rect 309839 498868 309915 503960
rect 311942 503860 312038 504852
rect 370968 504404 371064 505396
rect 370436 504308 371064 504404
rect 311942 503857 312296 503860
rect 311936 503761 311942 503857
rect 312038 503764 312296 503857
rect 312038 503761 312044 503764
rect 370968 503316 371064 504308
rect 376448 528984 376544 529953
rect 435474 529528 435570 530520
rect 435312 529432 435570 529528
rect 376448 528888 377076 528984
rect 376448 527896 376544 528888
rect 435474 528866 435570 529432
rect 437262 560436 437358 560570
rect 496288 560881 497171 560884
rect 437262 560340 437520 560436
rect 437262 559348 437358 560340
rect 496288 559892 496384 560881
rect 495756 559796 496384 559892
rect 437262 559252 437520 559348
rect 437262 558260 437358 559252
rect 496288 558804 496384 559796
rect 495756 558708 496384 558804
rect 437262 558164 437520 558260
rect 437262 557172 437358 558164
rect 496288 557716 496384 558708
rect 495756 557620 496384 557716
rect 437262 557076 437520 557172
rect 437262 556084 437358 557076
rect 496288 556628 496384 557620
rect 495756 556532 496384 556628
rect 437262 555988 437520 556084
rect 437262 554996 437358 555988
rect 496288 555540 496384 556532
rect 495756 555444 496384 555540
rect 437262 554900 437520 554996
rect 437262 553908 437358 554900
rect 496288 554452 496384 555444
rect 495756 554356 496384 554452
rect 437262 553812 437520 553908
rect 437262 552820 437358 553812
rect 496288 553364 496384 554356
rect 495756 553268 496384 553364
rect 437262 552724 437520 552820
rect 437262 551732 437358 552724
rect 496288 552276 496384 553268
rect 495756 552180 496384 552276
rect 437262 551636 437520 551732
rect 437262 550644 437358 551636
rect 496288 551188 496384 552180
rect 495756 551092 496384 551188
rect 437262 550548 437520 550644
rect 437262 549556 437358 550548
rect 496288 550100 496384 551092
rect 495756 550004 496384 550100
rect 437262 549460 437520 549556
rect 437262 548468 437358 549460
rect 496288 549012 496384 550004
rect 495756 548916 496384 549012
rect 437262 548372 437520 548468
rect 437262 547380 437358 548372
rect 496288 547924 496384 548916
rect 495756 547828 496384 547924
rect 437262 547284 437520 547380
rect 437262 546292 437358 547284
rect 496288 546836 496384 547828
rect 495756 546740 496384 546836
rect 437262 546196 437520 546292
rect 437262 545204 437358 546196
rect 496288 545748 496384 546740
rect 495756 545652 496384 545748
rect 437262 545108 437520 545204
rect 437262 544116 437358 545108
rect 496288 544660 496384 545652
rect 495756 544564 496384 544660
rect 437262 544020 437520 544116
rect 437262 543028 437358 544020
rect 496288 543572 496384 544564
rect 495756 543476 496384 543572
rect 437262 542932 437520 543028
rect 437262 541940 437358 542932
rect 496288 542484 496384 543476
rect 495756 542388 496384 542484
rect 437262 541844 437520 541940
rect 437262 540852 437358 541844
rect 496288 541396 496384 542388
rect 495756 541300 496384 541396
rect 437262 540756 437520 540852
rect 437262 539764 437358 540756
rect 496288 540308 496384 541300
rect 495756 540212 496384 540308
rect 437262 539668 437520 539764
rect 437262 538676 437358 539668
rect 496288 539220 496384 540212
rect 495756 539124 496384 539220
rect 437262 538580 437520 538676
rect 437262 537588 437358 538580
rect 496288 538132 496384 539124
rect 495756 538036 496384 538132
rect 437262 537492 437520 537588
rect 437262 536500 437358 537492
rect 496288 537044 496384 538036
rect 495756 536948 496384 537044
rect 437262 536404 437520 536500
rect 437262 535412 437358 536404
rect 496288 535956 496384 536948
rect 495756 535860 496384 535956
rect 437262 535316 437520 535412
rect 437262 534324 437358 535316
rect 496288 534868 496384 535860
rect 495756 534772 496384 534868
rect 437262 534228 437520 534324
rect 437262 533236 437358 534228
rect 496288 533780 496384 534772
rect 495756 533684 496384 533780
rect 437262 533140 437520 533236
rect 437262 532148 437358 533140
rect 496288 532692 496384 533684
rect 495756 532596 496384 532692
rect 437262 532052 437520 532148
rect 437262 531060 437358 532052
rect 496288 531604 496384 532596
rect 495756 531508 496384 531604
rect 437262 530964 437520 531060
rect 496288 530977 496384 531508
rect 501768 560536 501864 561528
rect 560794 561392 560888 561420
rect 560536 561001 560888 561080
rect 560536 560984 560786 561001
rect 560780 560905 560786 560984
rect 560894 560905 560900 561001
rect 560794 560781 560888 560905
rect 501768 560440 502396 560536
rect 501768 559448 501864 560440
rect 560794 559992 560890 560781
rect 560536 559896 560890 559992
rect 501768 559352 502396 559448
rect 501768 558360 501864 559352
rect 560794 558904 560890 559896
rect 560632 558808 560890 558904
rect 501768 558264 502396 558360
rect 501768 557272 501864 558264
rect 560794 557816 560890 558808
rect 560632 557720 560890 557816
rect 501768 557176 502396 557272
rect 501768 556184 501864 557176
rect 560794 556728 560890 557720
rect 560632 556632 560890 556728
rect 501768 556088 502396 556184
rect 501768 555096 501864 556088
rect 560794 555640 560890 556632
rect 560632 555544 560890 555640
rect 501768 555000 502396 555096
rect 501768 554008 501864 555000
rect 560794 554552 560890 555544
rect 560632 554456 560890 554552
rect 501768 553912 502396 554008
rect 501768 552920 501864 553912
rect 560794 553464 560890 554456
rect 560632 553368 560890 553464
rect 501768 552824 502396 552920
rect 501768 551832 501864 552824
rect 560794 552376 560890 553368
rect 560632 552280 560890 552376
rect 501768 551736 502396 551832
rect 501768 550744 501864 551736
rect 560794 551288 560890 552280
rect 560632 551192 560890 551288
rect 501768 550648 502396 550744
rect 501768 549656 501864 550648
rect 560794 550200 560890 551192
rect 560632 550104 560890 550200
rect 501768 549560 502396 549656
rect 501768 548568 501864 549560
rect 560794 549112 560890 550104
rect 560632 549016 560890 549112
rect 501768 548472 502396 548568
rect 501768 547480 501864 548472
rect 560794 548024 560890 549016
rect 560632 547928 560890 548024
rect 501768 547384 502396 547480
rect 501768 546392 501864 547384
rect 560794 546936 560890 547928
rect 560632 546840 560890 546936
rect 501768 546296 502396 546392
rect 501768 545304 501864 546296
rect 560794 545848 560890 546840
rect 560632 545752 560890 545848
rect 501768 545208 502396 545304
rect 501768 544216 501864 545208
rect 560794 544760 560890 545752
rect 560632 544664 560890 544760
rect 501768 544120 502396 544216
rect 501768 543128 501864 544120
rect 560794 543672 560890 544664
rect 560632 543576 560890 543672
rect 501768 543032 502396 543128
rect 501768 542040 501864 543032
rect 560794 542584 560890 543576
rect 560632 542488 560890 542584
rect 501768 541944 502396 542040
rect 501768 540952 501864 541944
rect 560794 541496 560890 542488
rect 560632 541400 560890 541496
rect 501768 540856 502396 540952
rect 501768 539864 501864 540856
rect 560794 540408 560890 541400
rect 560632 540312 560890 540408
rect 501768 539768 502396 539864
rect 501768 538776 501864 539768
rect 560794 539320 560890 540312
rect 560632 539224 560890 539320
rect 501768 538680 502396 538776
rect 501768 537688 501864 538680
rect 560794 538232 560890 539224
rect 560632 538136 560890 538232
rect 501768 537592 502396 537688
rect 501768 536600 501864 537592
rect 560794 537144 560890 538136
rect 560632 537048 560890 537144
rect 501768 536504 502396 536600
rect 501768 535512 501864 536504
rect 560794 536056 560890 537048
rect 560632 535960 560890 536056
rect 501768 535416 502396 535512
rect 501768 534424 501864 535416
rect 560794 534968 560890 535960
rect 560632 534872 560890 534968
rect 501768 534328 502396 534424
rect 501768 533336 501864 534328
rect 560794 533880 560890 534872
rect 560632 533784 560890 533880
rect 501768 533240 502396 533336
rect 501768 532248 501864 533240
rect 560794 532792 560890 533784
rect 560632 532696 560890 532792
rect 501768 532152 502396 532248
rect 501768 531160 501864 532152
rect 560794 531704 560890 532696
rect 560632 531608 560890 531704
rect 501768 531064 502396 531160
rect 501768 530977 501864 531064
rect 437262 529972 437358 530964
rect 496288 530929 501864 530977
rect 496288 530516 498496 530929
rect 495756 530420 498496 530516
rect 496288 530001 498496 530420
rect 499520 530072 501864 530929
rect 560794 530977 560890 531608
rect 560794 530929 566821 530977
rect 560794 530616 564289 530929
rect 560632 530520 564289 530616
rect 499520 530001 502396 530072
rect 496288 529976 502396 530001
rect 560794 530001 564289 530520
rect 565313 530001 566821 530929
rect 437262 529876 437520 529972
rect 496288 529953 501864 529976
rect 437262 528884 437358 529876
rect 496288 529428 496384 529953
rect 495756 529332 496384 529428
rect 436432 528866 437075 528869
rect 435474 528863 437075 528866
rect 437262 528863 437520 528884
rect 435474 528815 437520 528863
rect 435474 528440 436583 528815
rect 435312 528344 436583 528440
rect 435474 528143 436583 528344
rect 437273 528788 437520 528815
rect 437273 528143 437358 528788
rect 496288 528340 496384 529332
rect 495756 528244 496384 528340
rect 435474 528071 437358 528143
rect 435474 528058 437075 528071
rect 376448 527800 377076 527896
rect 376448 526808 376544 527800
rect 435474 527352 435570 528058
rect 435312 527256 435570 527352
rect 376448 526712 377076 526808
rect 376448 525720 376544 526712
rect 435474 526264 435570 527256
rect 435312 526168 435570 526264
rect 376448 525624 377076 525720
rect 376448 524632 376544 525624
rect 435474 525176 435570 526168
rect 435312 525080 435570 525176
rect 376448 524536 377076 524632
rect 376448 523544 376544 524536
rect 435474 524088 435570 525080
rect 435312 523992 435570 524088
rect 376448 523448 377076 523544
rect 376448 522456 376544 523448
rect 435474 523000 435570 523992
rect 435312 522904 435570 523000
rect 376448 522360 377076 522456
rect 376448 521368 376544 522360
rect 435474 521912 435570 522904
rect 435312 521816 435570 521912
rect 376448 521272 377076 521368
rect 376448 520280 376544 521272
rect 435474 520824 435570 521816
rect 435312 520728 435570 520824
rect 376448 520184 377076 520280
rect 376448 519192 376544 520184
rect 435474 519736 435570 520728
rect 435312 519640 435570 519736
rect 376448 519096 377076 519192
rect 376448 518104 376544 519096
rect 435474 518648 435570 519640
rect 435312 518552 435570 518648
rect 376448 518008 377076 518104
rect 376448 517016 376544 518008
rect 435474 517560 435570 518552
rect 435312 517464 435570 517560
rect 376448 516920 377076 517016
rect 376448 515928 376544 516920
rect 435474 516472 435570 517464
rect 435312 516376 435570 516472
rect 376448 515832 377076 515928
rect 376448 514840 376544 515832
rect 435474 515384 435570 516376
rect 435312 515288 435570 515384
rect 376448 514744 377076 514840
rect 376448 513752 376544 514744
rect 435474 514296 435570 515288
rect 435312 514200 435570 514296
rect 376448 513656 377076 513752
rect 376448 512664 376544 513656
rect 435474 513208 435570 514200
rect 435312 513112 435570 513208
rect 376448 512568 377076 512664
rect 376448 511576 376544 512568
rect 435474 512120 435570 513112
rect 435312 512024 435570 512120
rect 376448 511480 377076 511576
rect 376448 510488 376544 511480
rect 435474 511032 435570 512024
rect 435312 510936 435570 511032
rect 376448 510392 377076 510488
rect 376448 509400 376544 510392
rect 435474 509944 435570 510936
rect 435312 509848 435570 509944
rect 376448 509304 377076 509400
rect 376448 508312 376544 509304
rect 435474 508856 435570 509848
rect 435312 508760 435570 508856
rect 376448 508216 377076 508312
rect 376448 507224 376544 508216
rect 435474 507768 435570 508760
rect 435312 507672 435570 507768
rect 376448 507128 377076 507224
rect 376448 506136 376544 507128
rect 435474 506680 435570 507672
rect 435312 506584 435570 506680
rect 376448 506040 377076 506136
rect 376448 505048 376544 506040
rect 435474 505592 435570 506584
rect 435312 505496 435570 505592
rect 376448 504952 377076 505048
rect 376448 503960 376544 504952
rect 435474 504504 435570 505496
rect 435312 504408 435570 504504
rect 375632 503864 377076 503960
rect 370340 503220 371880 503316
rect 311936 503007 311942 503103
rect 312038 503007 312044 503103
rect 311942 498864 312038 503007
rect 311942 498768 312200 498864
rect 311942 497776 312038 498768
rect 371784 498320 371880 503220
rect 375632 498964 375728 503864
rect 435474 503416 435570 504408
rect 437262 527796 437358 528071
rect 437262 527700 437520 527796
rect 437262 526708 437358 527700
rect 496288 527252 496384 528244
rect 495756 527156 496384 527252
rect 437262 526612 437520 526708
rect 437262 525620 437358 526612
rect 496288 526164 496384 527156
rect 495756 526068 496384 526164
rect 437262 525524 437520 525620
rect 437262 524532 437358 525524
rect 496288 525076 496384 526068
rect 495756 524980 496384 525076
rect 437262 524436 437520 524532
rect 437262 523444 437358 524436
rect 496288 523988 496384 524980
rect 495756 523892 496384 523988
rect 437262 523348 437520 523444
rect 437262 522356 437358 523348
rect 496288 522900 496384 523892
rect 495756 522804 496384 522900
rect 437262 522260 437520 522356
rect 437262 521268 437358 522260
rect 496288 521812 496384 522804
rect 495756 521716 496384 521812
rect 437262 521172 437520 521268
rect 437262 520180 437358 521172
rect 496288 520724 496384 521716
rect 495756 520628 496384 520724
rect 437262 520084 437520 520180
rect 437262 519092 437358 520084
rect 496288 519636 496384 520628
rect 495756 519540 496384 519636
rect 437262 518996 437520 519092
rect 437262 518004 437358 518996
rect 496288 518548 496384 519540
rect 495756 518452 496384 518548
rect 437262 517908 437520 518004
rect 437262 516916 437358 517908
rect 496288 517460 496384 518452
rect 495756 517364 496384 517460
rect 437262 516820 437520 516916
rect 437262 515828 437358 516820
rect 496288 516372 496384 517364
rect 495756 516276 496384 516372
rect 437262 515732 437520 515828
rect 437262 514740 437358 515732
rect 496288 515284 496384 516276
rect 495756 515188 496384 515284
rect 437262 514644 437520 514740
rect 437262 513652 437358 514644
rect 496288 514196 496384 515188
rect 495756 514100 496384 514196
rect 437262 513556 437520 513652
rect 437262 512564 437358 513556
rect 496288 513108 496384 514100
rect 495756 513012 496384 513108
rect 437262 512468 437520 512564
rect 437262 511476 437358 512468
rect 496288 512020 496384 513012
rect 495756 511924 496384 512020
rect 437262 511380 437520 511476
rect 437262 510388 437358 511380
rect 496288 510932 496384 511924
rect 495756 510836 496384 510932
rect 437262 510292 437520 510388
rect 437262 509300 437358 510292
rect 496288 509844 496384 510836
rect 495756 509748 496384 509844
rect 437262 509204 437520 509300
rect 437262 508212 437358 509204
rect 496288 508756 496384 509748
rect 495756 508660 496384 508756
rect 437262 508116 437520 508212
rect 437262 507124 437358 508116
rect 496288 507668 496384 508660
rect 495756 507572 496384 507668
rect 437262 507028 437520 507124
rect 437262 506036 437358 507028
rect 496288 506580 496384 507572
rect 495756 506484 496384 506580
rect 437262 505940 437520 506036
rect 437262 504948 437358 505940
rect 496288 505492 496384 506484
rect 495756 505396 496384 505492
rect 437262 504852 437616 504948
rect 437262 503860 437358 504852
rect 496288 504404 496384 505396
rect 495756 504308 496384 504404
rect 437262 503857 437616 503860
rect 437256 503761 437262 503857
rect 437358 503764 437616 503857
rect 437358 503761 437364 503764
rect 435312 503320 435570 503416
rect 435474 499177 435570 503320
rect 496288 503316 496384 504308
rect 501768 528984 501864 529953
rect 560794 529953 566821 530001
rect 560794 529528 560890 529953
rect 560632 529432 560890 529528
rect 501768 528888 502396 528984
rect 501768 527896 501864 528888
rect 560794 528440 560890 529432
rect 560632 528344 560890 528440
rect 501768 527800 502396 527896
rect 501768 526808 501864 527800
rect 560794 527352 560890 528344
rect 560632 527256 560890 527352
rect 501768 526712 502396 526808
rect 501768 525720 501864 526712
rect 560794 526264 560890 527256
rect 560632 526168 560890 526264
rect 501768 525624 502396 525720
rect 501768 524632 501864 525624
rect 560794 525176 560890 526168
rect 560632 525080 560890 525176
rect 501768 524536 502396 524632
rect 501768 523544 501864 524536
rect 560794 524088 560890 525080
rect 560632 523992 560890 524088
rect 501768 523448 502396 523544
rect 501768 522456 501864 523448
rect 560794 523000 560890 523992
rect 560632 522904 560890 523000
rect 501768 522360 502396 522456
rect 501768 521368 501864 522360
rect 560794 521912 560890 522904
rect 560632 521816 560890 521912
rect 501768 521272 502396 521368
rect 501768 520280 501864 521272
rect 560794 520824 560890 521816
rect 560632 520728 560890 520824
rect 501768 520184 502396 520280
rect 501768 519192 501864 520184
rect 560794 519736 560890 520728
rect 560632 519640 560890 519736
rect 501768 519096 502396 519192
rect 501768 518104 501864 519096
rect 560794 518648 560890 519640
rect 560632 518552 560890 518648
rect 501768 518008 502396 518104
rect 501768 517016 501864 518008
rect 560794 517560 560890 518552
rect 560632 517464 560890 517560
rect 501768 516920 502396 517016
rect 501768 515928 501864 516920
rect 560794 516472 560890 517464
rect 560632 516376 560890 516472
rect 501768 515832 502396 515928
rect 501768 514840 501864 515832
rect 560794 515384 560890 516376
rect 560632 515288 560890 515384
rect 501768 514744 502396 514840
rect 501768 513752 501864 514744
rect 560794 514296 560890 515288
rect 560632 514200 560890 514296
rect 501768 513656 502396 513752
rect 501768 512664 501864 513656
rect 560794 513208 560890 514200
rect 560632 513112 560890 513208
rect 501768 512568 502396 512664
rect 501768 511576 501864 512568
rect 560794 512120 560890 513112
rect 560632 512024 560890 512120
rect 501768 511480 502396 511576
rect 501768 510488 501864 511480
rect 560794 511032 560890 512024
rect 560632 510936 560890 511032
rect 501768 510392 502396 510488
rect 501768 509400 501864 510392
rect 560794 509944 560890 510936
rect 560632 509848 560890 509944
rect 501768 509304 502396 509400
rect 501768 508312 501864 509304
rect 560794 508856 560890 509848
rect 560632 508760 560890 508856
rect 501768 508216 502396 508312
rect 501768 507224 501864 508216
rect 560794 507768 560890 508760
rect 560632 507672 560890 507768
rect 501768 507128 502396 507224
rect 501768 506136 501864 507128
rect 560794 506680 560890 507672
rect 560632 506584 560890 506680
rect 501768 506040 502396 506136
rect 501768 505048 501864 506040
rect 560794 505592 560890 506584
rect 560632 505496 560890 505592
rect 501768 504952 502396 505048
rect 501768 503960 501864 504952
rect 560794 504504 560890 505496
rect 560632 504408 560890 504504
rect 500952 503864 502396 503960
rect 495660 503220 497200 503316
rect 437256 503007 437262 503103
rect 437358 503007 437364 503103
rect 435468 499081 435474 499177
rect 435570 499081 435576 499177
rect 375632 498868 377172 498964
rect 370436 498224 371880 498320
rect 311942 497680 312200 497776
rect 311942 496688 312038 497680
rect 370968 497232 371064 498224
rect 370436 497136 371064 497232
rect 311942 496592 312200 496688
rect 311942 495600 312038 496592
rect 370968 496144 371064 497136
rect 370436 496048 371064 496144
rect 311942 495504 312200 495600
rect 311942 494512 312038 495504
rect 370968 495056 371064 496048
rect 370436 494960 371064 495056
rect 311942 494416 312200 494512
rect 311942 493424 312038 494416
rect 370968 493968 371064 494960
rect 370436 493872 371064 493968
rect 311942 493328 312200 493424
rect 311942 492336 312038 493328
rect 370968 492880 371064 493872
rect 370436 492784 371064 492880
rect 311942 492240 312200 492336
rect 311942 491248 312038 492240
rect 370968 491792 371064 492784
rect 370436 491696 371064 491792
rect 311942 491152 312200 491248
rect 311942 490160 312038 491152
rect 370968 490704 371064 491696
rect 370436 490608 371064 490704
rect 311942 490064 312200 490160
rect 311942 489072 312038 490064
rect 370968 489616 371064 490608
rect 370436 489520 371064 489616
rect 311942 488976 312200 489072
rect 311942 487984 312038 488976
rect 370968 488528 371064 489520
rect 370436 488432 371064 488528
rect 311942 487888 312200 487984
rect 311942 486896 312038 487888
rect 370968 487440 371064 488432
rect 370436 487344 371064 487440
rect 311942 486800 312200 486896
rect 311942 485808 312038 486800
rect 370968 486352 371064 487344
rect 370436 486256 371064 486352
rect 311942 485712 312200 485808
rect 311942 484720 312038 485712
rect 370968 485264 371064 486256
rect 370436 485168 371064 485264
rect 311942 484624 312200 484720
rect 311942 483632 312038 484624
rect 370968 484176 371064 485168
rect 370436 484080 371064 484176
rect 311942 483536 312200 483632
rect 311942 482544 312038 483536
rect 370968 483088 371064 484080
rect 370436 482992 371064 483088
rect 311942 482448 312200 482544
rect 311942 481456 312038 482448
rect 370968 482000 371064 482992
rect 370436 481904 371064 482000
rect 311942 481360 312200 481456
rect 311942 480368 312038 481360
rect 370968 480912 371064 481904
rect 370436 480816 371064 480912
rect 311942 480272 312200 480368
rect 311942 479280 312038 480272
rect 370968 479824 371064 480816
rect 370436 479728 371064 479824
rect 311942 479184 312200 479280
rect 311942 478192 312038 479184
rect 370968 478736 371064 479728
rect 370436 478640 371064 478736
rect 311942 478096 312200 478192
rect 311942 477104 312038 478096
rect 370968 477648 371064 478640
rect 370436 477552 371064 477648
rect 311942 477008 312200 477104
rect 311942 476016 312038 477008
rect 370968 476560 371064 477552
rect 370436 476464 371064 476560
rect 311942 475920 312200 476016
rect 311942 474928 312038 475920
rect 370968 475472 371064 476464
rect 370436 475376 371064 475472
rect 311942 474832 312200 474928
rect 311942 473840 312038 474832
rect 370968 474384 371064 475376
rect 370436 474288 371064 474384
rect 311942 473744 312200 473840
rect 311942 472752 312038 473744
rect 370968 473296 371064 474288
rect 370436 473200 371064 473296
rect 311942 472656 312200 472752
rect 311942 471664 312038 472656
rect 370968 472208 371064 473200
rect 370436 472112 371064 472208
rect 311942 471568 312200 471664
rect 311942 470576 312038 471568
rect 370968 471120 371064 472112
rect 370436 471024 371064 471120
rect 311942 470480 312200 470576
rect 311942 469488 312038 470480
rect 370968 470032 371064 471024
rect 370436 469936 371064 470032
rect 311942 469392 312200 469488
rect 311942 468400 312038 469392
rect 370968 468944 371064 469936
rect 370436 468848 371064 468944
rect 311942 468317 312200 468400
rect 306149 468304 312200 468317
rect 370968 468317 371064 468848
rect 376448 497876 376544 498868
rect 437262 498864 437358 503007
rect 437262 498768 437520 498864
rect 435468 498420 435474 498423
rect 435216 498327 435474 498420
rect 435570 498327 435576 498423
rect 435216 498324 435570 498327
rect 376448 497780 377076 497876
rect 376448 496788 376544 497780
rect 435474 497332 435570 498324
rect 435216 497236 435570 497332
rect 376448 496692 377076 496788
rect 376448 495700 376544 496692
rect 435474 496244 435570 497236
rect 435312 496148 435570 496244
rect 376448 495604 377076 495700
rect 376448 494612 376544 495604
rect 435474 495156 435570 496148
rect 435312 495060 435570 495156
rect 376448 494516 377076 494612
rect 376448 493524 376544 494516
rect 435474 494068 435570 495060
rect 435312 493972 435570 494068
rect 376448 493428 377076 493524
rect 376448 492436 376544 493428
rect 435474 492980 435570 493972
rect 435312 492884 435570 492980
rect 376448 492340 377076 492436
rect 376448 491348 376544 492340
rect 435474 491892 435570 492884
rect 435312 491796 435570 491892
rect 376448 491252 377076 491348
rect 376448 490260 376544 491252
rect 435474 490804 435570 491796
rect 435312 490708 435570 490804
rect 376448 490164 377076 490260
rect 376448 489172 376544 490164
rect 435474 489716 435570 490708
rect 435312 489620 435570 489716
rect 376448 489076 377076 489172
rect 376448 488084 376544 489076
rect 435474 488628 435570 489620
rect 435312 488532 435570 488628
rect 376448 487988 377076 488084
rect 376448 486996 376544 487988
rect 435474 487540 435570 488532
rect 435312 487444 435570 487540
rect 376448 486900 377076 486996
rect 376448 485908 376544 486900
rect 435474 486452 435570 487444
rect 435312 486356 435570 486452
rect 376448 485812 377076 485908
rect 376448 484820 376544 485812
rect 435474 485364 435570 486356
rect 435312 485268 435570 485364
rect 376448 484724 377076 484820
rect 376448 483732 376544 484724
rect 435474 484276 435570 485268
rect 435312 484180 435570 484276
rect 376448 483636 377076 483732
rect 376448 482644 376544 483636
rect 435474 483188 435570 484180
rect 435312 483092 435570 483188
rect 376448 482548 377076 482644
rect 376448 481556 376544 482548
rect 435474 482100 435570 483092
rect 435312 482004 435570 482100
rect 376448 481460 377076 481556
rect 376448 480468 376544 481460
rect 435474 481012 435570 482004
rect 435312 480916 435570 481012
rect 376448 480372 377076 480468
rect 376448 479380 376544 480372
rect 435474 479924 435570 480916
rect 435312 479828 435570 479924
rect 376448 479284 377076 479380
rect 376448 478292 376544 479284
rect 435474 478836 435570 479828
rect 435312 478740 435570 478836
rect 376448 478196 377076 478292
rect 376448 477204 376544 478196
rect 435474 477748 435570 478740
rect 435312 477652 435570 477748
rect 376448 477108 377076 477204
rect 376448 476116 376544 477108
rect 435474 476660 435570 477652
rect 435312 476564 435570 476660
rect 376448 476020 377076 476116
rect 376448 475028 376544 476020
rect 435474 475572 435570 476564
rect 435312 475476 435570 475572
rect 376448 474932 377076 475028
rect 376448 473940 376544 474932
rect 435474 474484 435570 475476
rect 435312 474388 435570 474484
rect 376448 473844 377076 473940
rect 376448 472852 376544 473844
rect 435474 473396 435570 474388
rect 435312 473300 435570 473396
rect 376448 472756 377076 472852
rect 376448 471764 376544 472756
rect 435474 472308 435570 473300
rect 435312 472212 435570 472308
rect 376448 471668 377076 471764
rect 376448 470676 376544 471668
rect 435474 471220 435570 472212
rect 435312 471124 435570 471220
rect 376448 470580 377076 470676
rect 376448 469588 376544 470580
rect 435474 470132 435570 471124
rect 435312 470036 435570 470132
rect 376448 469492 377076 469588
rect 376448 468500 376544 469492
rect 435474 469044 435570 470036
rect 435312 468948 435570 469044
rect 376448 468404 377076 468500
rect 376448 468317 376544 468404
rect 306149 468269 312038 468304
rect 306149 467341 307383 468269
rect 308407 467341 312038 468269
rect 370968 468269 376544 468317
rect 370968 467856 373176 468269
rect 370436 467760 373176 467856
rect 306149 467312 312038 467341
rect 370968 467341 373176 467760
rect 374200 467412 376544 468269
rect 435474 467956 435570 468948
rect 435312 467860 435570 467956
rect 374200 467341 377076 467412
rect 370968 467316 377076 467341
rect 306149 467293 312200 467312
rect 311942 467216 312200 467293
rect 370968 467293 376544 467316
rect 311942 466224 312038 467216
rect 370968 466768 371064 467293
rect 370436 466672 371064 466768
rect 311942 466128 312200 466224
rect 311942 465136 312038 466128
rect 370968 465680 371064 466672
rect 370436 465584 371064 465680
rect 311942 465040 312200 465136
rect 311942 464048 312038 465040
rect 370968 464592 371064 465584
rect 370436 464496 371064 464592
rect 311942 463952 312200 464048
rect 311942 462960 312038 463952
rect 370968 463504 371064 464496
rect 370436 463408 371064 463504
rect 311942 462864 312200 462960
rect 311942 461872 312038 462864
rect 370968 462416 371064 463408
rect 370436 462320 371064 462416
rect 311942 461776 312200 461872
rect 311942 460784 312038 461776
rect 370968 461328 371064 462320
rect 370436 461232 371064 461328
rect 311942 460688 312200 460784
rect 311942 459696 312038 460688
rect 370968 460240 371064 461232
rect 370436 460144 371064 460240
rect 311942 459600 312200 459696
rect 311942 458608 312038 459600
rect 370968 459152 371064 460144
rect 370436 459056 371064 459152
rect 311942 458512 312200 458608
rect 311942 457520 312038 458512
rect 370968 458064 371064 459056
rect 370436 457968 371064 458064
rect 311942 457424 312200 457520
rect 311942 456432 312038 457424
rect 370968 456976 371064 457968
rect 370436 456880 371064 456976
rect 311942 456336 312200 456432
rect 311942 455344 312038 456336
rect 370968 455888 371064 456880
rect 370436 455792 371064 455888
rect 311942 455248 312200 455344
rect 311942 454256 312038 455248
rect 370968 454800 371064 455792
rect 370436 454704 371064 454800
rect 311942 454160 312200 454256
rect 311942 453168 312038 454160
rect 370968 453712 371064 454704
rect 370436 453616 371064 453712
rect 311942 453072 312200 453168
rect 311942 452080 312038 453072
rect 370968 452624 371064 453616
rect 370436 452528 371064 452624
rect 311942 451984 312200 452080
rect 311942 450992 312038 451984
rect 370968 451536 371064 452528
rect 370436 451440 371064 451536
rect 311942 450896 312200 450992
rect 311942 449904 312038 450896
rect 370968 450448 371064 451440
rect 370436 450352 371064 450448
rect 311942 449808 312200 449904
rect 311942 448816 312038 449808
rect 370968 449360 371064 450352
rect 370436 449264 371064 449360
rect 311942 448720 312200 448816
rect 311942 447728 312038 448720
rect 370968 448272 371064 449264
rect 370436 448176 371064 448272
rect 311942 447632 312200 447728
rect 311942 446640 312038 447632
rect 370968 447184 371064 448176
rect 370436 447088 371064 447184
rect 311942 446544 312200 446640
rect 311942 445552 312038 446544
rect 370968 446096 371064 447088
rect 370436 446000 371064 446096
rect 311942 445456 312200 445552
rect 311942 444464 312038 445456
rect 370968 445008 371064 446000
rect 370436 444912 371064 445008
rect 311942 444368 312200 444464
rect 311942 443376 312038 444368
rect 370968 443920 371064 444912
rect 370436 443824 371064 443920
rect 311942 443280 312200 443376
rect 311942 442288 312038 443280
rect 370968 442832 371064 443824
rect 370436 442736 371064 442832
rect 311942 442192 312296 442288
rect 311942 441403 312038 442192
rect 370968 441744 371064 442736
rect 370436 441648 371064 441744
rect 309868 436219 309915 441303
rect 311944 441279 312038 441403
rect 311932 441183 311938 441279
rect 312046 441200 312052 441279
rect 312046 441183 312296 441200
rect 311944 441104 312296 441183
rect 311944 440764 312038 440792
rect 370968 440656 371064 441648
rect 376448 466324 376544 467293
rect 435474 466868 435570 467860
rect 435312 466772 435570 466868
rect 376448 466228 377076 466324
rect 376448 465236 376544 466228
rect 435474 466211 435570 466772
rect 437262 497776 437358 498768
rect 497104 498320 497200 503220
rect 500952 498964 501048 503864
rect 560794 503416 560890 504408
rect 560632 503320 560890 503416
rect 560794 499177 560890 503320
rect 560788 499081 560794 499177
rect 560890 499081 560896 499177
rect 500952 498868 502492 498964
rect 566745 498868 566821 503960
rect 495756 498224 497200 498320
rect 437262 497680 437520 497776
rect 437262 496688 437358 497680
rect 496288 497232 496384 498224
rect 495756 497136 496384 497232
rect 437262 496592 437520 496688
rect 437262 495600 437358 496592
rect 496288 496144 496384 497136
rect 495756 496048 496384 496144
rect 437262 495504 437520 495600
rect 437262 494512 437358 495504
rect 496288 495056 496384 496048
rect 495756 494960 496384 495056
rect 437262 494416 437520 494512
rect 437262 493424 437358 494416
rect 496288 493968 496384 494960
rect 495756 493872 496384 493968
rect 437262 493328 437520 493424
rect 437262 492336 437358 493328
rect 496288 492880 496384 493872
rect 495756 492784 496384 492880
rect 437262 492240 437520 492336
rect 437262 491248 437358 492240
rect 496288 491792 496384 492784
rect 495756 491696 496384 491792
rect 437262 491152 437520 491248
rect 437262 490160 437358 491152
rect 496288 490704 496384 491696
rect 495756 490608 496384 490704
rect 437262 490064 437520 490160
rect 437262 489072 437358 490064
rect 496288 489616 496384 490608
rect 495756 489520 496384 489616
rect 437262 488976 437520 489072
rect 437262 487984 437358 488976
rect 496288 488528 496384 489520
rect 495756 488432 496384 488528
rect 437262 487888 437520 487984
rect 437262 486896 437358 487888
rect 496288 487440 496384 488432
rect 495756 487344 496384 487440
rect 437262 486800 437520 486896
rect 437262 485808 437358 486800
rect 496288 486352 496384 487344
rect 495756 486256 496384 486352
rect 437262 485712 437520 485808
rect 437262 484720 437358 485712
rect 496288 485264 496384 486256
rect 495756 485168 496384 485264
rect 437262 484624 437520 484720
rect 437262 483632 437358 484624
rect 496288 484176 496384 485168
rect 495756 484080 496384 484176
rect 437262 483536 437520 483632
rect 437262 482544 437358 483536
rect 496288 483088 496384 484080
rect 495756 482992 496384 483088
rect 437262 482448 437520 482544
rect 437262 481456 437358 482448
rect 496288 482000 496384 482992
rect 495756 481904 496384 482000
rect 437262 481360 437520 481456
rect 437262 480368 437358 481360
rect 496288 480912 496384 481904
rect 495756 480816 496384 480912
rect 437262 480272 437520 480368
rect 437262 479280 437358 480272
rect 496288 479824 496384 480816
rect 495756 479728 496384 479824
rect 437262 479184 437520 479280
rect 437262 478192 437358 479184
rect 496288 478736 496384 479728
rect 495756 478640 496384 478736
rect 437262 478096 437520 478192
rect 437262 477104 437358 478096
rect 496288 477648 496384 478640
rect 495756 477552 496384 477648
rect 437262 477008 437520 477104
rect 437262 476016 437358 477008
rect 496288 476560 496384 477552
rect 495756 476464 496384 476560
rect 437262 475920 437520 476016
rect 437262 474928 437358 475920
rect 496288 475472 496384 476464
rect 495756 475376 496384 475472
rect 437262 474832 437520 474928
rect 437262 473840 437358 474832
rect 496288 474384 496384 475376
rect 495756 474288 496384 474384
rect 437262 473744 437520 473840
rect 437262 472752 437358 473744
rect 496288 473296 496384 474288
rect 495756 473200 496384 473296
rect 437262 472656 437520 472752
rect 437262 471664 437358 472656
rect 496288 472208 496384 473200
rect 495756 472112 496384 472208
rect 437262 471568 437520 471664
rect 437262 470576 437358 471568
rect 496288 471120 496384 472112
rect 495756 471024 496384 471120
rect 437262 470480 437520 470576
rect 437262 469488 437358 470480
rect 496288 470032 496384 471024
rect 495756 469936 496384 470032
rect 437262 469392 437520 469488
rect 437262 468400 437358 469392
rect 496288 468944 496384 469936
rect 495756 468848 496384 468944
rect 437262 468304 437520 468400
rect 496288 468317 496384 468848
rect 501768 497876 501864 498868
rect 560788 498420 560794 498423
rect 560536 498327 560794 498420
rect 560890 498327 560896 498423
rect 560536 498324 560890 498327
rect 501768 497780 502396 497876
rect 501768 496788 501864 497780
rect 560794 497332 560890 498324
rect 560536 497236 560890 497332
rect 501768 496692 502396 496788
rect 501768 495700 501864 496692
rect 560794 496244 560890 497236
rect 560632 496148 560890 496244
rect 501768 495604 502396 495700
rect 501768 494612 501864 495604
rect 560794 495156 560890 496148
rect 560632 495060 560890 495156
rect 501768 494516 502396 494612
rect 501768 493524 501864 494516
rect 560794 494068 560890 495060
rect 560632 493972 560890 494068
rect 501768 493428 502396 493524
rect 501768 492436 501864 493428
rect 560794 492980 560890 493972
rect 560632 492884 560890 492980
rect 501768 492340 502396 492436
rect 501768 491348 501864 492340
rect 560794 491892 560890 492884
rect 560632 491796 560890 491892
rect 501768 491252 502396 491348
rect 501768 490260 501864 491252
rect 560794 490804 560890 491796
rect 560632 490708 560890 490804
rect 501768 490164 502396 490260
rect 501768 489172 501864 490164
rect 560794 489716 560890 490708
rect 560632 489620 560890 489716
rect 501768 489076 502396 489172
rect 501768 488084 501864 489076
rect 560794 488628 560890 489620
rect 560632 488532 560890 488628
rect 501768 487988 502396 488084
rect 501768 486996 501864 487988
rect 560794 487540 560890 488532
rect 560632 487444 560890 487540
rect 501768 486900 502396 486996
rect 501768 485908 501864 486900
rect 560794 486452 560890 487444
rect 560632 486356 560890 486452
rect 501768 485812 502396 485908
rect 501768 484820 501864 485812
rect 560794 485364 560890 486356
rect 560632 485268 560890 485364
rect 501768 484724 502396 484820
rect 501768 483732 501864 484724
rect 560794 484276 560890 485268
rect 560632 484180 560890 484276
rect 501768 483636 502396 483732
rect 501768 482644 501864 483636
rect 560794 483188 560890 484180
rect 560632 483092 560890 483188
rect 501768 482548 502396 482644
rect 501768 481556 501864 482548
rect 560794 482100 560890 483092
rect 560632 482004 560890 482100
rect 501768 481460 502396 481556
rect 501768 480468 501864 481460
rect 560794 481012 560890 482004
rect 560632 480916 560890 481012
rect 501768 480372 502396 480468
rect 501768 479380 501864 480372
rect 560794 479924 560890 480916
rect 560632 479828 560890 479924
rect 501768 479284 502396 479380
rect 501768 478292 501864 479284
rect 560794 478836 560890 479828
rect 560632 478740 560890 478836
rect 501768 478196 502396 478292
rect 501768 477204 501864 478196
rect 560794 477748 560890 478740
rect 560632 477652 560890 477748
rect 501768 477108 502396 477204
rect 501768 476116 501864 477108
rect 560794 476660 560890 477652
rect 560632 476564 560890 476660
rect 501768 476020 502396 476116
rect 501768 475028 501864 476020
rect 560794 475572 560890 476564
rect 560632 475476 560890 475572
rect 501768 474932 502396 475028
rect 501768 473940 501864 474932
rect 560794 474484 560890 475476
rect 560632 474388 560890 474484
rect 501768 473844 502396 473940
rect 501768 472852 501864 473844
rect 560794 473396 560890 474388
rect 560632 473300 560890 473396
rect 501768 472756 502396 472852
rect 501768 471764 501864 472756
rect 560794 472308 560890 473300
rect 560632 472212 560890 472308
rect 501768 471668 502396 471764
rect 501768 470676 501864 471668
rect 560794 471220 560890 472212
rect 560632 471124 560890 471220
rect 501768 470580 502396 470676
rect 501768 469588 501864 470580
rect 560794 470132 560890 471124
rect 560632 470036 560890 470132
rect 501768 469492 502396 469588
rect 501768 468500 501864 469492
rect 560794 469044 560890 470036
rect 560632 468948 560890 469044
rect 501768 468404 502396 468500
rect 501768 468317 501864 468404
rect 437262 467312 437358 468304
rect 496288 468269 501864 468317
rect 496288 467856 498496 468269
rect 495756 467760 498496 467856
rect 496288 467341 498496 467760
rect 499520 467412 501864 468269
rect 560794 468317 560890 468948
rect 560794 468269 566821 468317
rect 560794 467956 564289 468269
rect 560632 467860 564289 467956
rect 499520 467341 502396 467412
rect 496288 467316 502396 467341
rect 560794 467341 564289 467860
rect 565313 467341 566821 468269
rect 437262 467216 437520 467312
rect 496288 467293 501864 467316
rect 437262 466224 437358 467216
rect 496288 466768 496384 467293
rect 495756 466672 496384 466768
rect 435474 466209 436462 466211
rect 435474 466203 437075 466209
rect 437262 466203 437520 466224
rect 435474 466155 437520 466203
rect 435474 465780 436583 466155
rect 435312 465684 436583 465780
rect 435474 465483 436583 465684
rect 437273 466128 437520 466155
rect 437273 465483 437358 466128
rect 496288 465680 496384 466672
rect 495756 465584 496384 465680
rect 435474 465411 437358 465483
rect 435474 465403 437075 465411
rect 376448 465140 377076 465236
rect 376448 464148 376544 465140
rect 435474 464692 435570 465403
rect 436432 465398 437075 465403
rect 435312 464596 435570 464692
rect 376448 464052 377076 464148
rect 376448 463060 376544 464052
rect 435474 463604 435570 464596
rect 435312 463508 435570 463604
rect 376448 462964 377076 463060
rect 376448 461972 376544 462964
rect 435474 462516 435570 463508
rect 435312 462420 435570 462516
rect 376448 461876 377076 461972
rect 376448 460884 376544 461876
rect 435474 461428 435570 462420
rect 435312 461332 435570 461428
rect 376448 460788 377076 460884
rect 376448 459796 376544 460788
rect 435474 460340 435570 461332
rect 435312 460244 435570 460340
rect 376448 459700 377076 459796
rect 376448 458708 376544 459700
rect 435474 459252 435570 460244
rect 435312 459156 435570 459252
rect 376448 458612 377076 458708
rect 376448 457620 376544 458612
rect 435474 458164 435570 459156
rect 435312 458068 435570 458164
rect 376448 457524 377076 457620
rect 376448 456532 376544 457524
rect 435474 457076 435570 458068
rect 435312 456980 435570 457076
rect 376448 456436 377076 456532
rect 376448 455444 376544 456436
rect 435474 455988 435570 456980
rect 435312 455892 435570 455988
rect 376448 455348 377076 455444
rect 376448 454356 376544 455348
rect 435474 454900 435570 455892
rect 435312 454804 435570 454900
rect 376448 454260 377076 454356
rect 376448 453268 376544 454260
rect 435474 453812 435570 454804
rect 435312 453716 435570 453812
rect 376448 453172 377076 453268
rect 376448 452180 376544 453172
rect 435474 452724 435570 453716
rect 435312 452628 435570 452724
rect 376448 452084 377076 452180
rect 376448 451092 376544 452084
rect 435474 451636 435570 452628
rect 435312 451540 435570 451636
rect 376448 450996 377076 451092
rect 376448 450004 376544 450996
rect 435474 450548 435570 451540
rect 435312 450452 435570 450548
rect 376448 449908 377076 450004
rect 376448 448916 376544 449908
rect 435474 449460 435570 450452
rect 435312 449364 435570 449460
rect 376448 448820 377076 448916
rect 376448 447828 376544 448820
rect 435474 448372 435570 449364
rect 435312 448276 435570 448372
rect 376448 447732 377076 447828
rect 376448 446740 376544 447732
rect 435474 447284 435570 448276
rect 435312 447188 435570 447284
rect 376448 446644 377076 446740
rect 376448 445652 376544 446644
rect 435474 446196 435570 447188
rect 435312 446100 435570 446196
rect 376448 445556 377076 445652
rect 376448 444564 376544 445556
rect 435474 445108 435570 446100
rect 435312 445012 435570 445108
rect 376448 444468 377076 444564
rect 376448 443476 376544 444468
rect 435474 444020 435570 445012
rect 435312 443924 435570 444020
rect 376448 443380 377076 443476
rect 376448 442388 376544 443380
rect 435474 442932 435570 443924
rect 435312 442836 435570 442932
rect 376448 442292 377076 442388
rect 376448 441303 376544 442292
rect 435474 441844 435570 442836
rect 435312 441748 435570 441844
rect 375661 441300 376544 441303
rect 435474 441614 435570 441748
rect 437262 465136 437358 465411
rect 437262 465040 437520 465136
rect 437262 464048 437358 465040
rect 496288 464592 496384 465584
rect 495756 464496 496384 464592
rect 437262 463952 437520 464048
rect 437262 462960 437358 463952
rect 496288 463504 496384 464496
rect 495756 463408 496384 463504
rect 437262 462864 437520 462960
rect 437262 461872 437358 462864
rect 496288 462416 496384 463408
rect 495756 462320 496384 462416
rect 437262 461776 437520 461872
rect 437262 460784 437358 461776
rect 496288 461328 496384 462320
rect 495756 461232 496384 461328
rect 437262 460688 437520 460784
rect 437262 459696 437358 460688
rect 496288 460240 496384 461232
rect 495756 460144 496384 460240
rect 437262 459600 437520 459696
rect 437262 458608 437358 459600
rect 496288 459152 496384 460144
rect 495756 459056 496384 459152
rect 437262 458512 437520 458608
rect 437262 457520 437358 458512
rect 496288 458064 496384 459056
rect 495756 457968 496384 458064
rect 437262 457424 437520 457520
rect 437262 456432 437358 457424
rect 496288 456976 496384 457968
rect 495756 456880 496384 456976
rect 437262 456336 437520 456432
rect 437262 455344 437358 456336
rect 496288 455888 496384 456880
rect 495756 455792 496384 455888
rect 437262 455248 437520 455344
rect 437262 454256 437358 455248
rect 496288 454800 496384 455792
rect 495756 454704 496384 454800
rect 437262 454160 437520 454256
rect 437262 453168 437358 454160
rect 496288 453712 496384 454704
rect 495756 453616 496384 453712
rect 437262 453072 437520 453168
rect 437262 452080 437358 453072
rect 496288 452624 496384 453616
rect 495756 452528 496384 452624
rect 437262 451984 437520 452080
rect 437262 450992 437358 451984
rect 496288 451536 496384 452528
rect 495756 451440 496384 451536
rect 437262 450896 437520 450992
rect 437262 449904 437358 450896
rect 496288 450448 496384 451440
rect 495756 450352 496384 450448
rect 437262 449808 437520 449904
rect 437262 448816 437358 449808
rect 496288 449360 496384 450352
rect 495756 449264 496384 449360
rect 437262 448720 437520 448816
rect 437262 447728 437358 448720
rect 496288 448272 496384 449264
rect 495756 448176 496384 448272
rect 437262 447632 437520 447728
rect 437262 446640 437358 447632
rect 496288 447184 496384 448176
rect 495756 447088 496384 447184
rect 437262 446544 437520 446640
rect 437262 445552 437358 446544
rect 496288 446096 496384 447088
rect 495756 446000 496384 446096
rect 437262 445456 437520 445552
rect 437262 444464 437358 445456
rect 496288 445008 496384 446000
rect 495756 444912 496384 445008
rect 437262 444368 437520 444464
rect 437262 443376 437358 444368
rect 496288 443920 496384 444912
rect 495756 443824 496384 443920
rect 437262 443280 437520 443376
rect 437262 442288 437358 443280
rect 496288 442832 496384 443824
rect 495756 442736 496384 442832
rect 437262 442192 437616 442288
rect 375661 441207 377076 441300
rect 370340 440645 371850 440656
rect 370340 440560 371851 440645
rect 309869 436208 309915 436219
rect 311944 440355 312040 440367
rect 311944 436204 312040 440259
rect 311944 436108 312200 436204
rect 311944 435250 312038 436108
rect 370436 435657 371064 435660
rect 371755 435657 371851 440560
rect 375661 436304 375757 441207
rect 376448 441204 377076 441207
rect 435474 440756 435568 441614
rect 437262 441403 437358 442192
rect 496288 441744 496384 442736
rect 495756 441648 496384 441744
rect 437264 441279 437358 441403
rect 437252 441183 437258 441279
rect 437366 441200 437372 441279
rect 437366 441183 437616 441200
rect 437264 441104 437616 441183
rect 437264 440764 437358 440792
rect 435312 440660 435568 440756
rect 435472 436605 435568 440660
rect 496288 440656 496384 441648
rect 501768 466324 501864 467293
rect 560794 467293 566821 467341
rect 560794 466868 560890 467293
rect 560632 466772 560890 466868
rect 501768 466228 502396 466324
rect 501768 465236 501864 466228
rect 560794 465780 560890 466772
rect 560632 465684 560890 465780
rect 501768 465140 502396 465236
rect 501768 464148 501864 465140
rect 560794 464692 560890 465684
rect 560632 464596 560890 464692
rect 501768 464052 502396 464148
rect 501768 463060 501864 464052
rect 560794 463604 560890 464596
rect 560632 463508 560890 463604
rect 501768 462964 502396 463060
rect 501768 461972 501864 462964
rect 560794 462516 560890 463508
rect 560632 462420 560890 462516
rect 501768 461876 502396 461972
rect 501768 460884 501864 461876
rect 560794 461428 560890 462420
rect 560632 461332 560890 461428
rect 501768 460788 502396 460884
rect 501768 459796 501864 460788
rect 560794 460340 560890 461332
rect 560632 460244 560890 460340
rect 501768 459700 502396 459796
rect 501768 458708 501864 459700
rect 560794 459252 560890 460244
rect 560632 459156 560890 459252
rect 501768 458612 502396 458708
rect 501768 457620 501864 458612
rect 560794 458164 560890 459156
rect 560632 458068 560890 458164
rect 501768 457524 502396 457620
rect 501768 456532 501864 457524
rect 560794 457076 560890 458068
rect 560632 456980 560890 457076
rect 501768 456436 502396 456532
rect 501768 455444 501864 456436
rect 560794 455988 560890 456980
rect 560632 455892 560890 455988
rect 501768 455348 502396 455444
rect 501768 454356 501864 455348
rect 560794 454900 560890 455892
rect 560632 454804 560890 454900
rect 501768 454260 502396 454356
rect 501768 453268 501864 454260
rect 560794 453812 560890 454804
rect 560632 453716 560890 453812
rect 501768 453172 502396 453268
rect 501768 452180 501864 453172
rect 560794 452724 560890 453716
rect 560632 452628 560890 452724
rect 501768 452084 502396 452180
rect 501768 451092 501864 452084
rect 560794 451636 560890 452628
rect 560632 451540 560890 451636
rect 501768 450996 502396 451092
rect 501768 450004 501864 450996
rect 560794 450548 560890 451540
rect 560632 450452 560890 450548
rect 501768 449908 502396 450004
rect 501768 448916 501864 449908
rect 560794 449460 560890 450452
rect 560632 449364 560890 449460
rect 501768 448820 502396 448916
rect 501768 447828 501864 448820
rect 560794 448372 560890 449364
rect 560632 448276 560890 448372
rect 501768 447732 502396 447828
rect 501768 446740 501864 447732
rect 560794 447284 560890 448276
rect 560632 447188 560890 447284
rect 501768 446644 502396 446740
rect 501768 445652 501864 446644
rect 560794 446196 560890 447188
rect 560632 446100 560890 446196
rect 501768 445556 502396 445652
rect 501768 444564 501864 445556
rect 560794 445108 560890 446100
rect 560632 445012 560890 445108
rect 501768 444468 502396 444564
rect 501768 443476 501864 444468
rect 560794 444020 560890 445012
rect 560632 443924 560890 444020
rect 501768 443380 502396 443476
rect 501768 442388 501864 443380
rect 560794 442932 560890 443924
rect 560632 442836 560890 442932
rect 501768 442292 502396 442388
rect 501768 441303 501864 442292
rect 560794 441844 560890 442836
rect 560632 441748 560890 441844
rect 500981 441300 501864 441303
rect 560794 441614 560890 441748
rect 500981 441207 502396 441300
rect 495660 440645 497170 440656
rect 495660 440560 497171 440645
rect 435472 436497 435568 436509
rect 437264 440355 437360 440367
rect 375661 436219 377172 436304
rect 375662 436208 377172 436219
rect 370436 435564 371851 435657
rect 311942 435116 312038 435250
rect 370968 435561 371851 435564
rect 311942 435020 312200 435116
rect 311942 434028 312038 435020
rect 370968 434572 371064 435561
rect 370436 434476 371064 434572
rect 311942 433932 312200 434028
rect 311942 432940 312038 433932
rect 370968 433484 371064 434476
rect 370436 433388 371064 433484
rect 311942 432844 312200 432940
rect 311942 431852 312038 432844
rect 370968 432396 371064 433388
rect 370436 432300 371064 432396
rect 311942 431756 312200 431852
rect 311942 430764 312038 431756
rect 370968 431308 371064 432300
rect 370436 431212 371064 431308
rect 311942 430668 312200 430764
rect 311942 429676 312038 430668
rect 370968 430220 371064 431212
rect 370436 430124 371064 430220
rect 311942 429580 312200 429676
rect 311942 428588 312038 429580
rect 370968 429132 371064 430124
rect 370436 429036 371064 429132
rect 311942 428492 312200 428588
rect 311942 427500 312038 428492
rect 370968 428044 371064 429036
rect 370436 427948 371064 428044
rect 311942 427404 312200 427500
rect 311942 426412 312038 427404
rect 370968 426956 371064 427948
rect 370436 426860 371064 426956
rect 311942 426316 312200 426412
rect 311942 425324 312038 426316
rect 370968 425868 371064 426860
rect 370436 425772 371064 425868
rect 311942 425228 312200 425324
rect 311942 424236 312038 425228
rect 370968 424780 371064 425772
rect 370436 424684 371064 424780
rect 311942 424140 312200 424236
rect 311942 423148 312038 424140
rect 370968 423692 371064 424684
rect 370436 423596 371064 423692
rect 311942 423052 312200 423148
rect 311942 422060 312038 423052
rect 370968 422604 371064 423596
rect 370436 422508 371064 422604
rect 311942 421964 312200 422060
rect 311942 420972 312038 421964
rect 370968 421516 371064 422508
rect 370436 421420 371064 421516
rect 311942 420876 312200 420972
rect 311942 419884 312038 420876
rect 370968 420428 371064 421420
rect 370436 420332 371064 420428
rect 311942 419788 312200 419884
rect 311942 418796 312038 419788
rect 370968 419340 371064 420332
rect 370436 419244 371064 419340
rect 311942 418700 312200 418796
rect 311942 417708 312038 418700
rect 370968 418252 371064 419244
rect 370436 418156 371064 418252
rect 311942 417612 312200 417708
rect 311942 416620 312038 417612
rect 370968 417164 371064 418156
rect 370436 417068 371064 417164
rect 311942 416524 312200 416620
rect 311942 415532 312038 416524
rect 370968 416076 371064 417068
rect 370436 415980 371064 416076
rect 311942 415436 312200 415532
rect 311942 414444 312038 415436
rect 370968 414988 371064 415980
rect 370436 414892 371064 414988
rect 311942 414348 312200 414444
rect 311942 413356 312038 414348
rect 370968 413900 371064 414892
rect 370436 413804 371064 413900
rect 311942 413260 312200 413356
rect 311942 412268 312038 413260
rect 370968 412812 371064 413804
rect 370436 412716 371064 412812
rect 311942 412172 312200 412268
rect 311942 411180 312038 412172
rect 370968 411724 371064 412716
rect 370436 411628 371064 411724
rect 311942 411084 312200 411180
rect 311942 410092 312038 411084
rect 370968 410636 371064 411628
rect 370436 410540 371064 410636
rect 311942 409996 312200 410092
rect 311942 409004 312038 409996
rect 370968 409548 371064 410540
rect 370436 409452 371064 409548
rect 311942 408908 312200 409004
rect 311942 407916 312038 408908
rect 370968 408460 371064 409452
rect 370436 408364 371064 408460
rect 311942 407820 312200 407916
rect 311942 406828 312038 407820
rect 370968 407372 371064 408364
rect 370436 407276 371064 407372
rect 311942 406732 312200 406828
rect 311942 405740 312038 406732
rect 370968 406284 371064 407276
rect 370436 406188 371064 406284
rect 311942 405657 312200 405740
rect 306149 405644 312200 405657
rect 370968 405657 371064 406188
rect 376448 435216 376544 436208
rect 437264 436204 437360 440259
rect 437264 436108 437520 436204
rect 435474 436072 435568 436100
rect 435216 435681 435568 435760
rect 435216 435664 435466 435681
rect 435460 435585 435466 435664
rect 435574 435585 435580 435681
rect 435474 435461 435568 435585
rect 376448 435120 377076 435216
rect 376448 434128 376544 435120
rect 435474 434672 435570 435461
rect 437264 435250 437358 436108
rect 495756 435657 496384 435660
rect 497075 435657 497171 440560
rect 500981 436304 501077 441207
rect 501768 441204 502396 441207
rect 560794 440756 560888 441614
rect 560632 440660 560888 440756
rect 560792 436605 560888 440660
rect 560792 436497 560888 436509
rect 500981 436219 502492 436304
rect 566774 436219 566821 441303
rect 500982 436208 502492 436219
rect 566775 436208 566821 436219
rect 495756 435564 497171 435657
rect 435216 434576 435570 434672
rect 376448 434032 377076 434128
rect 376448 433040 376544 434032
rect 435474 433584 435570 434576
rect 435312 433488 435570 433584
rect 376448 432944 377076 433040
rect 376448 431952 376544 432944
rect 435474 432496 435570 433488
rect 435312 432400 435570 432496
rect 376448 431856 377076 431952
rect 376448 430864 376544 431856
rect 435474 431408 435570 432400
rect 435312 431312 435570 431408
rect 376448 430768 377076 430864
rect 376448 429776 376544 430768
rect 435474 430320 435570 431312
rect 435312 430224 435570 430320
rect 376448 429680 377076 429776
rect 376448 428688 376544 429680
rect 435474 429232 435570 430224
rect 435312 429136 435570 429232
rect 376448 428592 377076 428688
rect 376448 427600 376544 428592
rect 435474 428144 435570 429136
rect 435312 428048 435570 428144
rect 376448 427504 377076 427600
rect 376448 426512 376544 427504
rect 435474 427056 435570 428048
rect 435312 426960 435570 427056
rect 376448 426416 377076 426512
rect 376448 425424 376544 426416
rect 435474 425968 435570 426960
rect 435312 425872 435570 425968
rect 376448 425328 377076 425424
rect 376448 424336 376544 425328
rect 435474 424880 435570 425872
rect 435312 424784 435570 424880
rect 376448 424240 377076 424336
rect 376448 423248 376544 424240
rect 435474 423792 435570 424784
rect 435312 423696 435570 423792
rect 376448 423152 377076 423248
rect 376448 422160 376544 423152
rect 435474 422704 435570 423696
rect 435312 422608 435570 422704
rect 376448 422064 377076 422160
rect 376448 421072 376544 422064
rect 435474 421616 435570 422608
rect 435312 421520 435570 421616
rect 376448 420976 377076 421072
rect 376448 419984 376544 420976
rect 435474 420528 435570 421520
rect 435312 420432 435570 420528
rect 376448 419888 377076 419984
rect 376448 418896 376544 419888
rect 435474 419440 435570 420432
rect 435312 419344 435570 419440
rect 376448 418800 377076 418896
rect 376448 417808 376544 418800
rect 435474 418352 435570 419344
rect 435312 418256 435570 418352
rect 376448 417712 377076 417808
rect 376448 416720 376544 417712
rect 435474 417264 435570 418256
rect 435312 417168 435570 417264
rect 376448 416624 377076 416720
rect 376448 415632 376544 416624
rect 435474 416176 435570 417168
rect 435312 416080 435570 416176
rect 376448 415536 377076 415632
rect 376448 414544 376544 415536
rect 435474 415088 435570 416080
rect 435312 414992 435570 415088
rect 376448 414448 377076 414544
rect 376448 413456 376544 414448
rect 435474 414000 435570 414992
rect 435312 413904 435570 414000
rect 376448 413360 377076 413456
rect 376448 412368 376544 413360
rect 435474 412912 435570 413904
rect 435312 412816 435570 412912
rect 376448 412272 377076 412368
rect 376448 411280 376544 412272
rect 435474 411824 435570 412816
rect 435312 411728 435570 411824
rect 376448 411184 377076 411280
rect 376448 410192 376544 411184
rect 435474 410736 435570 411728
rect 435312 410640 435570 410736
rect 376448 410096 377076 410192
rect 376448 409104 376544 410096
rect 435474 409648 435570 410640
rect 435312 409552 435570 409648
rect 376448 409008 377076 409104
rect 376448 408016 376544 409008
rect 435474 408560 435570 409552
rect 435312 408464 435570 408560
rect 376448 407920 377076 408016
rect 376448 406928 376544 407920
rect 435474 407472 435570 408464
rect 435312 407376 435570 407472
rect 376448 406832 377076 406928
rect 376448 405840 376544 406832
rect 435474 406384 435570 407376
rect 435312 406288 435570 406384
rect 376448 405744 377076 405840
rect 376448 405657 376544 405744
rect 306149 405609 312038 405644
rect 306149 404681 307383 405609
rect 308407 404681 312038 405609
rect 370968 405609 376544 405657
rect 370968 405196 373176 405609
rect 370436 405100 373176 405196
rect 306149 404652 312038 404681
rect 370968 404681 373176 405100
rect 374200 404752 376544 405609
rect 435474 405296 435570 406288
rect 435312 405200 435570 405296
rect 374200 404681 377076 404752
rect 370968 404656 377076 404681
rect 306149 404633 312200 404652
rect 311942 404556 312200 404633
rect 370968 404633 376544 404656
rect 311942 403564 312038 404556
rect 370968 404108 371064 404633
rect 370436 404012 371064 404108
rect 311942 403468 312200 403564
rect 311942 402476 312038 403468
rect 370968 403020 371064 404012
rect 370436 402924 371064 403020
rect 311942 402380 312200 402476
rect 311942 401388 312038 402380
rect 370968 401932 371064 402924
rect 370436 401836 371064 401932
rect 311942 401292 312200 401388
rect 311942 400300 312038 401292
rect 370968 400844 371064 401836
rect 370436 400748 371064 400844
rect 311942 400204 312200 400300
rect 311942 399212 312038 400204
rect 370968 399756 371064 400748
rect 370436 399660 371064 399756
rect 311942 399116 312200 399212
rect 311942 398124 312038 399116
rect 370968 398668 371064 399660
rect 370436 398572 371064 398668
rect 311942 398028 312200 398124
rect 311942 397036 312038 398028
rect 370968 397580 371064 398572
rect 370436 397484 371064 397580
rect 311942 396940 312200 397036
rect 311942 395948 312038 396940
rect 370968 396492 371064 397484
rect 370436 396396 371064 396492
rect 311942 395852 312200 395948
rect 311942 394860 312038 395852
rect 370968 395404 371064 396396
rect 370436 395308 371064 395404
rect 311942 394764 312200 394860
rect 311942 393772 312038 394764
rect 370968 394316 371064 395308
rect 370436 394220 371064 394316
rect 311942 393676 312200 393772
rect 311942 392684 312038 393676
rect 370968 393228 371064 394220
rect 370436 393132 371064 393228
rect 311942 392588 312200 392684
rect 311942 391596 312038 392588
rect 370968 392140 371064 393132
rect 370436 392044 371064 392140
rect 311942 391500 312200 391596
rect 311942 390508 312038 391500
rect 370968 391052 371064 392044
rect 370436 390956 371064 391052
rect 311942 390412 312200 390508
rect 311942 389420 312038 390412
rect 370968 389964 371064 390956
rect 370436 389868 371064 389964
rect 311942 389324 312200 389420
rect 311942 388332 312038 389324
rect 370968 388876 371064 389868
rect 370436 388780 371064 388876
rect 311942 388236 312200 388332
rect 311942 387244 312038 388236
rect 370968 387788 371064 388780
rect 370436 387692 371064 387788
rect 311942 387148 312200 387244
rect 311942 386156 312038 387148
rect 370968 386700 371064 387692
rect 370436 386604 371064 386700
rect 311942 386060 312200 386156
rect 311942 385068 312038 386060
rect 370968 385612 371064 386604
rect 370436 385516 371064 385612
rect 311942 384972 312200 385068
rect 311942 383980 312038 384972
rect 370968 384524 371064 385516
rect 370436 384428 371064 384524
rect 311942 383884 312200 383980
rect 311942 382892 312038 383884
rect 370968 383436 371064 384428
rect 370436 383340 371064 383436
rect 311942 382796 312200 382892
rect 311942 381804 312038 382796
rect 370968 382348 371064 383340
rect 370436 382252 371064 382348
rect 311942 381708 312200 381804
rect 311942 380716 312038 381708
rect 370968 381260 371064 382252
rect 370436 381164 371064 381260
rect 311942 380620 312200 380716
rect 311942 379628 312038 380620
rect 370968 380172 371064 381164
rect 370436 380076 371064 380172
rect 311942 379532 312296 379628
rect 309839 373548 309915 378640
rect 311942 378540 312038 379532
rect 370968 379084 371064 380076
rect 370436 378988 371064 379084
rect 311942 378537 312296 378540
rect 311936 378441 311942 378537
rect 312038 378444 312296 378537
rect 312038 378441 312044 378444
rect 370968 377996 371064 378988
rect 376448 403664 376544 404633
rect 435474 404208 435570 405200
rect 435312 404112 435570 404208
rect 376448 403568 377076 403664
rect 376448 402576 376544 403568
rect 435474 403550 435570 404112
rect 437262 435116 437358 435250
rect 496288 435561 497171 435564
rect 437262 435020 437520 435116
rect 437262 434028 437358 435020
rect 496288 434572 496384 435561
rect 495756 434476 496384 434572
rect 437262 433932 437520 434028
rect 437262 432940 437358 433932
rect 496288 433484 496384 434476
rect 495756 433388 496384 433484
rect 437262 432844 437520 432940
rect 437262 431852 437358 432844
rect 496288 432396 496384 433388
rect 495756 432300 496384 432396
rect 437262 431756 437520 431852
rect 437262 430764 437358 431756
rect 496288 431308 496384 432300
rect 495756 431212 496384 431308
rect 437262 430668 437520 430764
rect 437262 429676 437358 430668
rect 496288 430220 496384 431212
rect 495756 430124 496384 430220
rect 437262 429580 437520 429676
rect 437262 428588 437358 429580
rect 496288 429132 496384 430124
rect 495756 429036 496384 429132
rect 437262 428492 437520 428588
rect 437262 427500 437358 428492
rect 496288 428044 496384 429036
rect 495756 427948 496384 428044
rect 437262 427404 437520 427500
rect 437262 426412 437358 427404
rect 496288 426956 496384 427948
rect 495756 426860 496384 426956
rect 437262 426316 437520 426412
rect 437262 425324 437358 426316
rect 496288 425868 496384 426860
rect 495756 425772 496384 425868
rect 437262 425228 437520 425324
rect 437262 424236 437358 425228
rect 496288 424780 496384 425772
rect 495756 424684 496384 424780
rect 437262 424140 437520 424236
rect 437262 423148 437358 424140
rect 496288 423692 496384 424684
rect 495756 423596 496384 423692
rect 437262 423052 437520 423148
rect 437262 422060 437358 423052
rect 496288 422604 496384 423596
rect 495756 422508 496384 422604
rect 437262 421964 437520 422060
rect 437262 420972 437358 421964
rect 496288 421516 496384 422508
rect 495756 421420 496384 421516
rect 437262 420876 437520 420972
rect 437262 419884 437358 420876
rect 496288 420428 496384 421420
rect 495756 420332 496384 420428
rect 437262 419788 437520 419884
rect 437262 418796 437358 419788
rect 496288 419340 496384 420332
rect 495756 419244 496384 419340
rect 437262 418700 437520 418796
rect 437262 417708 437358 418700
rect 496288 418252 496384 419244
rect 495756 418156 496384 418252
rect 437262 417612 437520 417708
rect 437262 416620 437358 417612
rect 496288 417164 496384 418156
rect 495756 417068 496384 417164
rect 437262 416524 437520 416620
rect 437262 415532 437358 416524
rect 496288 416076 496384 417068
rect 495756 415980 496384 416076
rect 437262 415436 437520 415532
rect 437262 414444 437358 415436
rect 496288 414988 496384 415980
rect 495756 414892 496384 414988
rect 437262 414348 437520 414444
rect 437262 413356 437358 414348
rect 496288 413900 496384 414892
rect 495756 413804 496384 413900
rect 437262 413260 437520 413356
rect 437262 412268 437358 413260
rect 496288 412812 496384 413804
rect 495756 412716 496384 412812
rect 437262 412172 437520 412268
rect 437262 411180 437358 412172
rect 496288 411724 496384 412716
rect 495756 411628 496384 411724
rect 437262 411084 437520 411180
rect 437262 410092 437358 411084
rect 496288 410636 496384 411628
rect 495756 410540 496384 410636
rect 437262 409996 437520 410092
rect 437262 409004 437358 409996
rect 496288 409548 496384 410540
rect 495756 409452 496384 409548
rect 437262 408908 437520 409004
rect 437262 407916 437358 408908
rect 496288 408460 496384 409452
rect 495756 408364 496384 408460
rect 437262 407820 437520 407916
rect 437262 406828 437358 407820
rect 496288 407372 496384 408364
rect 495756 407276 496384 407372
rect 437262 406732 437520 406828
rect 437262 405740 437358 406732
rect 496288 406284 496384 407276
rect 495756 406188 496384 406284
rect 437262 405644 437520 405740
rect 496288 405657 496384 406188
rect 501768 435216 501864 436208
rect 560794 436072 560888 436100
rect 560536 435681 560888 435760
rect 560536 435664 560786 435681
rect 560780 435585 560786 435664
rect 560894 435585 560900 435681
rect 560794 435461 560888 435585
rect 501768 435120 502396 435216
rect 501768 434128 501864 435120
rect 560794 434672 560890 435461
rect 560536 434576 560890 434672
rect 501768 434032 502396 434128
rect 501768 433040 501864 434032
rect 560794 433584 560890 434576
rect 560632 433488 560890 433584
rect 501768 432944 502396 433040
rect 501768 431952 501864 432944
rect 560794 432496 560890 433488
rect 560632 432400 560890 432496
rect 501768 431856 502396 431952
rect 501768 430864 501864 431856
rect 560794 431408 560890 432400
rect 560632 431312 560890 431408
rect 501768 430768 502396 430864
rect 501768 429776 501864 430768
rect 560794 430320 560890 431312
rect 560632 430224 560890 430320
rect 501768 429680 502396 429776
rect 501768 428688 501864 429680
rect 560794 429232 560890 430224
rect 560632 429136 560890 429232
rect 501768 428592 502396 428688
rect 501768 427600 501864 428592
rect 560794 428144 560890 429136
rect 560632 428048 560890 428144
rect 501768 427504 502396 427600
rect 501768 426512 501864 427504
rect 560794 427056 560890 428048
rect 560632 426960 560890 427056
rect 501768 426416 502396 426512
rect 501768 425424 501864 426416
rect 560794 425968 560890 426960
rect 560632 425872 560890 425968
rect 501768 425328 502396 425424
rect 501768 424336 501864 425328
rect 560794 424880 560890 425872
rect 560632 424784 560890 424880
rect 501768 424240 502396 424336
rect 501768 423248 501864 424240
rect 560794 423792 560890 424784
rect 560632 423696 560890 423792
rect 501768 423152 502396 423248
rect 501768 422160 501864 423152
rect 560794 422704 560890 423696
rect 560632 422608 560890 422704
rect 501768 422064 502396 422160
rect 501768 421072 501864 422064
rect 560794 421616 560890 422608
rect 560632 421520 560890 421616
rect 501768 420976 502396 421072
rect 501768 419984 501864 420976
rect 560794 420528 560890 421520
rect 560632 420432 560890 420528
rect 501768 419888 502396 419984
rect 501768 418896 501864 419888
rect 560794 419440 560890 420432
rect 560632 419344 560890 419440
rect 501768 418800 502396 418896
rect 501768 417808 501864 418800
rect 560794 418352 560890 419344
rect 560632 418256 560890 418352
rect 501768 417712 502396 417808
rect 501768 416720 501864 417712
rect 560794 417264 560890 418256
rect 560632 417168 560890 417264
rect 501768 416624 502396 416720
rect 501768 415632 501864 416624
rect 560794 416176 560890 417168
rect 560632 416080 560890 416176
rect 501768 415536 502396 415632
rect 501768 414544 501864 415536
rect 560794 415088 560890 416080
rect 560632 414992 560890 415088
rect 501768 414448 502396 414544
rect 501768 413456 501864 414448
rect 560794 414000 560890 414992
rect 560632 413904 560890 414000
rect 501768 413360 502396 413456
rect 501768 412368 501864 413360
rect 560794 412912 560890 413904
rect 560632 412816 560890 412912
rect 501768 412272 502396 412368
rect 501768 411280 501864 412272
rect 560794 411824 560890 412816
rect 560632 411728 560890 411824
rect 501768 411184 502396 411280
rect 501768 410192 501864 411184
rect 560794 410736 560890 411728
rect 560632 410640 560890 410736
rect 501768 410096 502396 410192
rect 501768 409104 501864 410096
rect 560794 409648 560890 410640
rect 560632 409552 560890 409648
rect 501768 409008 502396 409104
rect 501768 408016 501864 409008
rect 560794 408560 560890 409552
rect 560632 408464 560890 408560
rect 501768 407920 502396 408016
rect 501768 406928 501864 407920
rect 560794 407472 560890 408464
rect 560632 407376 560890 407472
rect 501768 406832 502396 406928
rect 501768 405840 501864 406832
rect 560794 406384 560890 407376
rect 560632 406288 560890 406384
rect 501768 405744 502396 405840
rect 501768 405657 501864 405744
rect 437262 404652 437358 405644
rect 496288 405609 501864 405657
rect 496288 405196 498496 405609
rect 495756 405100 498496 405196
rect 496288 404681 498496 405100
rect 499520 404752 501864 405609
rect 560794 405657 560890 406288
rect 560794 405609 566821 405657
rect 560794 405296 564289 405609
rect 560632 405200 564289 405296
rect 499520 404681 502396 404752
rect 496288 404656 502396 404681
rect 560794 404681 564289 405200
rect 565313 404681 566821 405609
rect 437262 404556 437520 404652
rect 496288 404633 501864 404656
rect 437262 403564 437358 404556
rect 496288 404108 496384 404633
rect 495756 404012 496384 404108
rect 435474 403549 436461 403550
rect 435474 403543 437075 403549
rect 437262 403543 437520 403564
rect 435474 403495 437520 403543
rect 435474 403120 436583 403495
rect 435312 403024 436583 403120
rect 435474 402823 436583 403024
rect 437273 403468 437520 403495
rect 437273 402823 437358 403468
rect 496288 403020 496384 404012
rect 495756 402924 496384 403020
rect 435474 402751 437358 402823
rect 435474 402742 437075 402751
rect 376448 402480 377076 402576
rect 376448 401488 376544 402480
rect 435474 402032 435570 402742
rect 436432 402738 437075 402742
rect 435312 401936 435570 402032
rect 376448 401392 377076 401488
rect 376448 400400 376544 401392
rect 435474 400944 435570 401936
rect 435312 400848 435570 400944
rect 376448 400304 377076 400400
rect 376448 399312 376544 400304
rect 435474 399856 435570 400848
rect 435312 399760 435570 399856
rect 376448 399216 377076 399312
rect 376448 398224 376544 399216
rect 435474 398768 435570 399760
rect 435312 398672 435570 398768
rect 376448 398128 377076 398224
rect 376448 397136 376544 398128
rect 435474 397680 435570 398672
rect 435312 397584 435570 397680
rect 376448 397040 377076 397136
rect 376448 396048 376544 397040
rect 435474 396592 435570 397584
rect 435312 396496 435570 396592
rect 376448 395952 377076 396048
rect 376448 394960 376544 395952
rect 435474 395504 435570 396496
rect 435312 395408 435570 395504
rect 376448 394864 377076 394960
rect 376448 393872 376544 394864
rect 435474 394416 435570 395408
rect 435312 394320 435570 394416
rect 376448 393776 377076 393872
rect 376448 392784 376544 393776
rect 435474 393328 435570 394320
rect 435312 393232 435570 393328
rect 376448 392688 377076 392784
rect 376448 391696 376544 392688
rect 435474 392240 435570 393232
rect 435312 392144 435570 392240
rect 376448 391600 377076 391696
rect 376448 390608 376544 391600
rect 435474 391152 435570 392144
rect 435312 391056 435570 391152
rect 376448 390512 377076 390608
rect 376448 389520 376544 390512
rect 435474 390064 435570 391056
rect 435312 389968 435570 390064
rect 376448 389424 377076 389520
rect 376448 388432 376544 389424
rect 435474 388976 435570 389968
rect 435312 388880 435570 388976
rect 376448 388336 377076 388432
rect 376448 387344 376544 388336
rect 435474 387888 435570 388880
rect 435312 387792 435570 387888
rect 376448 387248 377076 387344
rect 376448 386256 376544 387248
rect 435474 386800 435570 387792
rect 435312 386704 435570 386800
rect 376448 386160 377076 386256
rect 376448 385168 376544 386160
rect 435474 385712 435570 386704
rect 435312 385616 435570 385712
rect 376448 385072 377076 385168
rect 376448 384080 376544 385072
rect 435474 384624 435570 385616
rect 435312 384528 435570 384624
rect 376448 383984 377076 384080
rect 376448 382992 376544 383984
rect 435474 383536 435570 384528
rect 435312 383440 435570 383536
rect 376448 382896 377076 382992
rect 376448 381904 376544 382896
rect 435474 382448 435570 383440
rect 435312 382352 435570 382448
rect 376448 381808 377076 381904
rect 376448 380816 376544 381808
rect 435474 381360 435570 382352
rect 435312 381264 435570 381360
rect 376448 380720 377076 380816
rect 376448 379728 376544 380720
rect 435474 380272 435570 381264
rect 435312 380176 435570 380272
rect 376448 379632 377076 379728
rect 376448 378640 376544 379632
rect 435474 379184 435570 380176
rect 435312 379088 435570 379184
rect 375632 378544 377076 378640
rect 370340 377900 371880 377996
rect 311936 377687 311942 377783
rect 312038 377687 312044 377783
rect 311942 373544 312038 377687
rect 311942 373448 312200 373544
rect 311942 372456 312038 373448
rect 371784 373000 371880 377900
rect 375632 373644 375728 378544
rect 435474 378096 435570 379088
rect 437262 402476 437358 402751
rect 437262 402380 437520 402476
rect 437262 401388 437358 402380
rect 496288 401932 496384 402924
rect 495756 401836 496384 401932
rect 437262 401292 437520 401388
rect 437262 400300 437358 401292
rect 496288 400844 496384 401836
rect 495756 400748 496384 400844
rect 437262 400204 437520 400300
rect 437262 399212 437358 400204
rect 496288 399756 496384 400748
rect 495756 399660 496384 399756
rect 437262 399116 437520 399212
rect 437262 398124 437358 399116
rect 496288 398668 496384 399660
rect 495756 398572 496384 398668
rect 437262 398028 437520 398124
rect 437262 397036 437358 398028
rect 496288 397580 496384 398572
rect 495756 397484 496384 397580
rect 437262 396940 437520 397036
rect 437262 395948 437358 396940
rect 496288 396492 496384 397484
rect 495756 396396 496384 396492
rect 437262 395852 437520 395948
rect 437262 394860 437358 395852
rect 496288 395404 496384 396396
rect 495756 395308 496384 395404
rect 437262 394764 437520 394860
rect 437262 393772 437358 394764
rect 496288 394316 496384 395308
rect 495756 394220 496384 394316
rect 437262 393676 437520 393772
rect 437262 392684 437358 393676
rect 496288 393228 496384 394220
rect 495756 393132 496384 393228
rect 437262 392588 437520 392684
rect 437262 391596 437358 392588
rect 496288 392140 496384 393132
rect 495756 392044 496384 392140
rect 437262 391500 437520 391596
rect 437262 390508 437358 391500
rect 496288 391052 496384 392044
rect 495756 390956 496384 391052
rect 437262 390412 437520 390508
rect 437262 389420 437358 390412
rect 496288 389964 496384 390956
rect 495756 389868 496384 389964
rect 437262 389324 437520 389420
rect 437262 388332 437358 389324
rect 496288 388876 496384 389868
rect 495756 388780 496384 388876
rect 437262 388236 437520 388332
rect 437262 387244 437358 388236
rect 496288 387788 496384 388780
rect 495756 387692 496384 387788
rect 437262 387148 437520 387244
rect 437262 386156 437358 387148
rect 496288 386700 496384 387692
rect 495756 386604 496384 386700
rect 437262 386060 437520 386156
rect 437262 385068 437358 386060
rect 496288 385612 496384 386604
rect 495756 385516 496384 385612
rect 437262 384972 437520 385068
rect 437262 383980 437358 384972
rect 496288 384524 496384 385516
rect 495756 384428 496384 384524
rect 437262 383884 437520 383980
rect 437262 382892 437358 383884
rect 496288 383436 496384 384428
rect 495756 383340 496384 383436
rect 437262 382796 437520 382892
rect 437262 381804 437358 382796
rect 496288 382348 496384 383340
rect 495756 382252 496384 382348
rect 437262 381708 437520 381804
rect 437262 380716 437358 381708
rect 496288 381260 496384 382252
rect 495756 381164 496384 381260
rect 437262 380620 437520 380716
rect 437262 379628 437358 380620
rect 496288 380172 496384 381164
rect 495756 380076 496384 380172
rect 437262 379532 437616 379628
rect 437262 378540 437358 379532
rect 496288 379084 496384 380076
rect 495756 378988 496384 379084
rect 437262 378537 437616 378540
rect 437256 378441 437262 378537
rect 437358 378444 437616 378537
rect 437358 378441 437364 378444
rect 435312 378000 435570 378096
rect 435474 373857 435570 378000
rect 496288 377996 496384 378988
rect 501768 403664 501864 404633
rect 560794 404633 566821 404681
rect 560794 404208 560890 404633
rect 560632 404112 560890 404208
rect 501768 403568 502396 403664
rect 501768 402576 501864 403568
rect 560794 403120 560890 404112
rect 560632 403024 560890 403120
rect 501768 402480 502396 402576
rect 501768 401488 501864 402480
rect 560794 402032 560890 403024
rect 560632 401936 560890 402032
rect 501768 401392 502396 401488
rect 501768 400400 501864 401392
rect 560794 400944 560890 401936
rect 560632 400848 560890 400944
rect 501768 400304 502396 400400
rect 501768 399312 501864 400304
rect 560794 399856 560890 400848
rect 560632 399760 560890 399856
rect 501768 399216 502396 399312
rect 501768 398224 501864 399216
rect 560794 398768 560890 399760
rect 560632 398672 560890 398768
rect 501768 398128 502396 398224
rect 501768 397136 501864 398128
rect 560794 397680 560890 398672
rect 560632 397584 560890 397680
rect 501768 397040 502396 397136
rect 501768 396048 501864 397040
rect 560794 396592 560890 397584
rect 560632 396496 560890 396592
rect 501768 395952 502396 396048
rect 501768 394960 501864 395952
rect 560794 395504 560890 396496
rect 560632 395408 560890 395504
rect 501768 394864 502396 394960
rect 501768 393872 501864 394864
rect 560794 394416 560890 395408
rect 560632 394320 560890 394416
rect 501768 393776 502396 393872
rect 501768 392784 501864 393776
rect 560794 393328 560890 394320
rect 560632 393232 560890 393328
rect 501768 392688 502396 392784
rect 501768 391696 501864 392688
rect 560794 392240 560890 393232
rect 560632 392144 560890 392240
rect 501768 391600 502396 391696
rect 501768 390608 501864 391600
rect 560794 391152 560890 392144
rect 560632 391056 560890 391152
rect 501768 390512 502396 390608
rect 501768 389520 501864 390512
rect 560794 390064 560890 391056
rect 560632 389968 560890 390064
rect 501768 389424 502396 389520
rect 501768 388432 501864 389424
rect 560794 388976 560890 389968
rect 560632 388880 560890 388976
rect 501768 388336 502396 388432
rect 501768 387344 501864 388336
rect 560794 387888 560890 388880
rect 560632 387792 560890 387888
rect 501768 387248 502396 387344
rect 501768 386256 501864 387248
rect 560794 386800 560890 387792
rect 560632 386704 560890 386800
rect 501768 386160 502396 386256
rect 501768 385168 501864 386160
rect 560794 385712 560890 386704
rect 560632 385616 560890 385712
rect 501768 385072 502396 385168
rect 501768 384080 501864 385072
rect 560794 384624 560890 385616
rect 560632 384528 560890 384624
rect 501768 383984 502396 384080
rect 501768 382992 501864 383984
rect 560794 383536 560890 384528
rect 560632 383440 560890 383536
rect 501768 382896 502396 382992
rect 501768 381904 501864 382896
rect 560794 382448 560890 383440
rect 560632 382352 560890 382448
rect 501768 381808 502396 381904
rect 501768 380816 501864 381808
rect 560794 381360 560890 382352
rect 560632 381264 560890 381360
rect 501768 380720 502396 380816
rect 501768 379728 501864 380720
rect 560794 380272 560890 381264
rect 560632 380176 560890 380272
rect 501768 379632 502396 379728
rect 501768 378640 501864 379632
rect 560794 379184 560890 380176
rect 560632 379088 560890 379184
rect 500952 378544 502396 378640
rect 495660 377900 497200 377996
rect 437256 377687 437262 377783
rect 437358 377687 437364 377783
rect 435468 373761 435474 373857
rect 435570 373761 435576 373857
rect 375632 373548 377172 373644
rect 370436 372904 371880 373000
rect 311942 372360 312200 372456
rect 311942 371368 312038 372360
rect 370968 371912 371064 372904
rect 370436 371816 371064 371912
rect 311942 371272 312200 371368
rect 311942 370280 312038 371272
rect 370968 370824 371064 371816
rect 370436 370728 371064 370824
rect 311942 370184 312200 370280
rect 311942 369192 312038 370184
rect 370968 369736 371064 370728
rect 370436 369640 371064 369736
rect 311942 369096 312200 369192
rect 311942 368104 312038 369096
rect 370968 368648 371064 369640
rect 370436 368552 371064 368648
rect 311942 368008 312200 368104
rect 311942 367016 312038 368008
rect 370968 367560 371064 368552
rect 370436 367464 371064 367560
rect 311942 366920 312200 367016
rect 311942 365928 312038 366920
rect 370968 366472 371064 367464
rect 370436 366376 371064 366472
rect 311942 365832 312200 365928
rect 311942 364840 312038 365832
rect 370968 365384 371064 366376
rect 370436 365288 371064 365384
rect 311942 364744 312200 364840
rect 311942 363752 312038 364744
rect 370968 364296 371064 365288
rect 370436 364200 371064 364296
rect 311942 363656 312200 363752
rect 311942 362664 312038 363656
rect 370968 363208 371064 364200
rect 370436 363112 371064 363208
rect 311942 362568 312200 362664
rect 311942 361576 312038 362568
rect 370968 362120 371064 363112
rect 370436 362024 371064 362120
rect 311942 361480 312200 361576
rect 311942 360488 312038 361480
rect 370968 361032 371064 362024
rect 370436 360936 371064 361032
rect 311942 360392 312200 360488
rect 311942 359400 312038 360392
rect 370968 359944 371064 360936
rect 370436 359848 371064 359944
rect 311942 359304 312200 359400
rect 311942 358312 312038 359304
rect 370968 358856 371064 359848
rect 370436 358760 371064 358856
rect 311942 358216 312200 358312
rect 311942 357224 312038 358216
rect 370968 357768 371064 358760
rect 370436 357672 371064 357768
rect 311942 357128 312200 357224
rect 311942 356136 312038 357128
rect 370968 356680 371064 357672
rect 370436 356584 371064 356680
rect 311942 356040 312200 356136
rect 311942 355048 312038 356040
rect 370968 355592 371064 356584
rect 370436 355496 371064 355592
rect 311942 354952 312200 355048
rect 311942 353960 312038 354952
rect 370968 354504 371064 355496
rect 370436 354408 371064 354504
rect 311942 353864 312200 353960
rect 311942 352872 312038 353864
rect 370968 353416 371064 354408
rect 370436 353320 371064 353416
rect 311942 352776 312200 352872
rect 311942 351784 312038 352776
rect 370968 352328 371064 353320
rect 370436 352232 371064 352328
rect 311942 351688 312200 351784
rect 311942 350696 312038 351688
rect 370968 351240 371064 352232
rect 370436 351144 371064 351240
rect 311942 350600 312200 350696
rect 311942 349608 312038 350600
rect 370968 350152 371064 351144
rect 370436 350056 371064 350152
rect 311942 349512 312200 349608
rect 311942 348520 312038 349512
rect 370968 349064 371064 350056
rect 370436 348968 371064 349064
rect 311942 348424 312200 348520
rect 311942 347432 312038 348424
rect 370968 347976 371064 348968
rect 370436 347880 371064 347976
rect 311942 347336 312200 347432
rect 311942 346344 312038 347336
rect 370968 346888 371064 347880
rect 370436 346792 371064 346888
rect 311942 346248 312200 346344
rect 311942 345256 312038 346248
rect 370968 345800 371064 346792
rect 370436 345704 371064 345800
rect 311942 345160 312200 345256
rect 311942 344168 312038 345160
rect 370968 344712 371064 345704
rect 370436 344616 371064 344712
rect 311942 344072 312200 344168
rect 311942 343080 312038 344072
rect 370968 343624 371064 344616
rect 370436 343528 371064 343624
rect 311942 342997 312200 343080
rect 306149 342984 312200 342997
rect 370968 342997 371064 343528
rect 376448 372556 376544 373548
rect 437262 373544 437358 377687
rect 437262 373448 437520 373544
rect 435468 373100 435474 373103
rect 435216 373007 435474 373100
rect 435570 373007 435576 373103
rect 435216 373004 435570 373007
rect 376448 372460 377076 372556
rect 376448 371468 376544 372460
rect 435474 372012 435570 373004
rect 435216 371916 435570 372012
rect 376448 371372 377076 371468
rect 376448 370380 376544 371372
rect 435474 370924 435570 371916
rect 435312 370828 435570 370924
rect 376448 370284 377076 370380
rect 376448 369292 376544 370284
rect 435474 369836 435570 370828
rect 435312 369740 435570 369836
rect 376448 369196 377076 369292
rect 376448 368204 376544 369196
rect 435474 368748 435570 369740
rect 435312 368652 435570 368748
rect 376448 368108 377076 368204
rect 376448 367116 376544 368108
rect 435474 367660 435570 368652
rect 435312 367564 435570 367660
rect 376448 367020 377076 367116
rect 376448 366028 376544 367020
rect 435474 366572 435570 367564
rect 435312 366476 435570 366572
rect 376448 365932 377076 366028
rect 376448 364940 376544 365932
rect 435474 365484 435570 366476
rect 435312 365388 435570 365484
rect 376448 364844 377076 364940
rect 376448 363852 376544 364844
rect 435474 364396 435570 365388
rect 435312 364300 435570 364396
rect 376448 363756 377076 363852
rect 376448 362764 376544 363756
rect 435474 363308 435570 364300
rect 435312 363212 435570 363308
rect 376448 362668 377076 362764
rect 376448 361676 376544 362668
rect 435474 362220 435570 363212
rect 435312 362124 435570 362220
rect 376448 361580 377076 361676
rect 376448 360588 376544 361580
rect 435474 361132 435570 362124
rect 435312 361036 435570 361132
rect 376448 360492 377076 360588
rect 376448 359500 376544 360492
rect 435474 360044 435570 361036
rect 435312 359948 435570 360044
rect 376448 359404 377076 359500
rect 376448 358412 376544 359404
rect 435474 358956 435570 359948
rect 435312 358860 435570 358956
rect 376448 358316 377076 358412
rect 376448 357324 376544 358316
rect 435474 357868 435570 358860
rect 435312 357772 435570 357868
rect 376448 357228 377076 357324
rect 376448 356236 376544 357228
rect 435474 356780 435570 357772
rect 435312 356684 435570 356780
rect 376448 356140 377076 356236
rect 376448 355148 376544 356140
rect 435474 355692 435570 356684
rect 435312 355596 435570 355692
rect 376448 355052 377076 355148
rect 376448 354060 376544 355052
rect 435474 354604 435570 355596
rect 435312 354508 435570 354604
rect 376448 353964 377076 354060
rect 376448 352972 376544 353964
rect 435474 353516 435570 354508
rect 435312 353420 435570 353516
rect 376448 352876 377076 352972
rect 376448 351884 376544 352876
rect 435474 352428 435570 353420
rect 435312 352332 435570 352428
rect 376448 351788 377076 351884
rect 376448 350796 376544 351788
rect 435474 351340 435570 352332
rect 435312 351244 435570 351340
rect 376448 350700 377076 350796
rect 376448 349708 376544 350700
rect 435474 350252 435570 351244
rect 435312 350156 435570 350252
rect 376448 349612 377076 349708
rect 376448 348620 376544 349612
rect 435474 349164 435570 350156
rect 435312 349068 435570 349164
rect 376448 348524 377076 348620
rect 376448 347532 376544 348524
rect 435474 348076 435570 349068
rect 435312 347980 435570 348076
rect 376448 347436 377076 347532
rect 376448 346444 376544 347436
rect 435474 346988 435570 347980
rect 435312 346892 435570 346988
rect 376448 346348 377076 346444
rect 376448 345356 376544 346348
rect 435474 345900 435570 346892
rect 435312 345804 435570 345900
rect 376448 345260 377076 345356
rect 376448 344268 376544 345260
rect 435474 344812 435570 345804
rect 435312 344716 435570 344812
rect 376448 344172 377076 344268
rect 376448 343180 376544 344172
rect 435474 343724 435570 344716
rect 435312 343628 435570 343724
rect 376448 343084 377076 343180
rect 376448 342997 376544 343084
rect 306149 342949 312038 342984
rect 306149 342021 307383 342949
rect 308407 342021 312038 342949
rect 370968 342949 376544 342997
rect 370968 342536 373176 342949
rect 370436 342440 373176 342536
rect 306149 341992 312038 342021
rect 370968 342021 373176 342440
rect 374200 342092 376544 342949
rect 435474 342636 435570 343628
rect 435312 342540 435570 342636
rect 374200 342021 377076 342092
rect 370968 341996 377076 342021
rect 306149 341973 312200 341992
rect 311942 341896 312200 341973
rect 370968 341973 376544 341996
rect 311942 340904 312038 341896
rect 370968 341448 371064 341973
rect 370436 341352 371064 341448
rect 311942 340808 312200 340904
rect 311942 339816 312038 340808
rect 370968 340360 371064 341352
rect 370436 340264 371064 340360
rect 311942 339720 312200 339816
rect 311942 338728 312038 339720
rect 370968 339272 371064 340264
rect 370436 339176 371064 339272
rect 311942 338632 312200 338728
rect 311942 337640 312038 338632
rect 370968 338184 371064 339176
rect 370436 338088 371064 338184
rect 311942 337544 312200 337640
rect 311942 336552 312038 337544
rect 370968 337096 371064 338088
rect 370436 337000 371064 337096
rect 311942 336456 312200 336552
rect 311942 335464 312038 336456
rect 370968 336008 371064 337000
rect 370436 335912 371064 336008
rect 311942 335368 312200 335464
rect 311942 334376 312038 335368
rect 370968 334920 371064 335912
rect 370436 334824 371064 334920
rect 311942 334280 312200 334376
rect 311942 333288 312038 334280
rect 370968 333832 371064 334824
rect 370436 333736 371064 333832
rect 311942 333192 312200 333288
rect 311942 332200 312038 333192
rect 370968 332744 371064 333736
rect 370436 332648 371064 332744
rect 311942 332104 312200 332200
rect 311942 331112 312038 332104
rect 370968 331656 371064 332648
rect 370436 331560 371064 331656
rect 311942 331016 312200 331112
rect 311942 330024 312038 331016
rect 370968 330568 371064 331560
rect 370436 330472 371064 330568
rect 311942 329928 312200 330024
rect 311942 328936 312038 329928
rect 370968 329480 371064 330472
rect 370436 329384 371064 329480
rect 311942 328840 312200 328936
rect 311942 327848 312038 328840
rect 370968 328392 371064 329384
rect 370436 328296 371064 328392
rect 311942 327752 312200 327848
rect 311942 326760 312038 327752
rect 370968 327304 371064 328296
rect 370436 327208 371064 327304
rect 311942 326664 312200 326760
rect 311942 325672 312038 326664
rect 370968 326216 371064 327208
rect 370436 326120 371064 326216
rect 311942 325576 312200 325672
rect 311942 324584 312038 325576
rect 370968 325128 371064 326120
rect 370436 325032 371064 325128
rect 311942 324488 312200 324584
rect 311942 323496 312038 324488
rect 370968 324040 371064 325032
rect 370436 323944 371064 324040
rect 311942 323400 312200 323496
rect 311942 322408 312038 323400
rect 370968 322952 371064 323944
rect 370436 322856 371064 322952
rect 311942 322312 312200 322408
rect 311942 321320 312038 322312
rect 370968 321864 371064 322856
rect 370436 321768 371064 321864
rect 311942 321224 312200 321320
rect 311942 320232 312038 321224
rect 370968 320776 371064 321768
rect 370436 320680 371064 320776
rect 311942 320136 312200 320232
rect 311942 319144 312038 320136
rect 370968 319688 371064 320680
rect 370436 319592 371064 319688
rect 311942 319048 312200 319144
rect 311942 318056 312038 319048
rect 370968 318600 371064 319592
rect 370436 318504 371064 318600
rect 311942 317960 312200 318056
rect 311942 316968 312038 317960
rect 370968 317512 371064 318504
rect 370436 317416 371064 317512
rect 311942 316872 312296 316968
rect 311942 316083 312038 316872
rect 370968 316424 371064 317416
rect 370436 316328 371064 316424
rect 309868 310899 309915 315983
rect 311944 315959 312038 316083
rect 311932 315863 311938 315959
rect 312046 315880 312052 315959
rect 312046 315863 312296 315880
rect 311944 315784 312296 315863
rect 311944 315444 312038 315472
rect 370968 315336 371064 316328
rect 376448 341004 376544 341973
rect 435474 341548 435570 342540
rect 435312 341452 435570 341548
rect 376448 340908 377076 341004
rect 376448 339916 376544 340908
rect 435474 340882 435570 341452
rect 437262 372456 437358 373448
rect 497104 373000 497200 377900
rect 500952 373644 501048 378544
rect 560794 378096 560890 379088
rect 560632 378000 560890 378096
rect 560794 373857 560890 378000
rect 560788 373761 560794 373857
rect 560890 373761 560896 373857
rect 500952 373548 502492 373644
rect 566745 373548 566821 378640
rect 495756 372904 497200 373000
rect 437262 372360 437520 372456
rect 437262 371368 437358 372360
rect 496288 371912 496384 372904
rect 495756 371816 496384 371912
rect 437262 371272 437520 371368
rect 437262 370280 437358 371272
rect 496288 370824 496384 371816
rect 495756 370728 496384 370824
rect 437262 370184 437520 370280
rect 437262 369192 437358 370184
rect 496288 369736 496384 370728
rect 495756 369640 496384 369736
rect 437262 369096 437520 369192
rect 437262 368104 437358 369096
rect 496288 368648 496384 369640
rect 495756 368552 496384 368648
rect 437262 368008 437520 368104
rect 437262 367016 437358 368008
rect 496288 367560 496384 368552
rect 495756 367464 496384 367560
rect 437262 366920 437520 367016
rect 437262 365928 437358 366920
rect 496288 366472 496384 367464
rect 495756 366376 496384 366472
rect 437262 365832 437520 365928
rect 437262 364840 437358 365832
rect 496288 365384 496384 366376
rect 495756 365288 496384 365384
rect 437262 364744 437520 364840
rect 437262 363752 437358 364744
rect 496288 364296 496384 365288
rect 495756 364200 496384 364296
rect 437262 363656 437520 363752
rect 437262 362664 437358 363656
rect 496288 363208 496384 364200
rect 495756 363112 496384 363208
rect 437262 362568 437520 362664
rect 437262 361576 437358 362568
rect 496288 362120 496384 363112
rect 495756 362024 496384 362120
rect 437262 361480 437520 361576
rect 437262 360488 437358 361480
rect 496288 361032 496384 362024
rect 495756 360936 496384 361032
rect 437262 360392 437520 360488
rect 437262 359400 437358 360392
rect 496288 359944 496384 360936
rect 495756 359848 496384 359944
rect 437262 359304 437520 359400
rect 437262 358312 437358 359304
rect 496288 358856 496384 359848
rect 495756 358760 496384 358856
rect 437262 358216 437520 358312
rect 437262 357224 437358 358216
rect 496288 357768 496384 358760
rect 495756 357672 496384 357768
rect 437262 357128 437520 357224
rect 437262 356136 437358 357128
rect 496288 356680 496384 357672
rect 495756 356584 496384 356680
rect 437262 356040 437520 356136
rect 437262 355048 437358 356040
rect 496288 355592 496384 356584
rect 495756 355496 496384 355592
rect 437262 354952 437520 355048
rect 437262 353960 437358 354952
rect 496288 354504 496384 355496
rect 495756 354408 496384 354504
rect 437262 353864 437520 353960
rect 437262 352872 437358 353864
rect 496288 353416 496384 354408
rect 495756 353320 496384 353416
rect 437262 352776 437520 352872
rect 437262 351784 437358 352776
rect 496288 352328 496384 353320
rect 495756 352232 496384 352328
rect 437262 351688 437520 351784
rect 437262 350696 437358 351688
rect 496288 351240 496384 352232
rect 495756 351144 496384 351240
rect 437262 350600 437520 350696
rect 437262 349608 437358 350600
rect 496288 350152 496384 351144
rect 495756 350056 496384 350152
rect 437262 349512 437520 349608
rect 437262 348520 437358 349512
rect 496288 349064 496384 350056
rect 495756 348968 496384 349064
rect 437262 348424 437520 348520
rect 437262 347432 437358 348424
rect 496288 347976 496384 348968
rect 495756 347880 496384 347976
rect 437262 347336 437520 347432
rect 437262 346344 437358 347336
rect 496288 346888 496384 347880
rect 495756 346792 496384 346888
rect 437262 346248 437520 346344
rect 437262 345256 437358 346248
rect 496288 345800 496384 346792
rect 495756 345704 496384 345800
rect 437262 345160 437520 345256
rect 437262 344168 437358 345160
rect 496288 344712 496384 345704
rect 495756 344616 496384 344712
rect 437262 344072 437520 344168
rect 437262 343080 437358 344072
rect 496288 343624 496384 344616
rect 495756 343528 496384 343624
rect 437262 342984 437520 343080
rect 496288 342997 496384 343528
rect 501768 372556 501864 373548
rect 560788 373100 560794 373103
rect 560536 373007 560794 373100
rect 560890 373007 560896 373103
rect 560536 373004 560890 373007
rect 501768 372460 502396 372556
rect 501768 371468 501864 372460
rect 560794 372012 560890 373004
rect 560536 371916 560890 372012
rect 501768 371372 502396 371468
rect 501768 370380 501864 371372
rect 560794 370924 560890 371916
rect 560632 370828 560890 370924
rect 501768 370284 502396 370380
rect 501768 369292 501864 370284
rect 560794 369836 560890 370828
rect 560632 369740 560890 369836
rect 501768 369196 502396 369292
rect 501768 368204 501864 369196
rect 560794 368748 560890 369740
rect 560632 368652 560890 368748
rect 501768 368108 502396 368204
rect 501768 367116 501864 368108
rect 560794 367660 560890 368652
rect 560632 367564 560890 367660
rect 501768 367020 502396 367116
rect 501768 366028 501864 367020
rect 560794 366572 560890 367564
rect 560632 366476 560890 366572
rect 501768 365932 502396 366028
rect 501768 364940 501864 365932
rect 560794 365484 560890 366476
rect 560632 365388 560890 365484
rect 501768 364844 502396 364940
rect 501768 363852 501864 364844
rect 560794 364396 560890 365388
rect 560632 364300 560890 364396
rect 501768 363756 502396 363852
rect 501768 362764 501864 363756
rect 560794 363308 560890 364300
rect 560632 363212 560890 363308
rect 501768 362668 502396 362764
rect 501768 361676 501864 362668
rect 560794 362220 560890 363212
rect 560632 362124 560890 362220
rect 501768 361580 502396 361676
rect 501768 360588 501864 361580
rect 560794 361132 560890 362124
rect 560632 361036 560890 361132
rect 501768 360492 502396 360588
rect 501768 359500 501864 360492
rect 560794 360044 560890 361036
rect 560632 359948 560890 360044
rect 501768 359404 502396 359500
rect 501768 358412 501864 359404
rect 560794 358956 560890 359948
rect 560632 358860 560890 358956
rect 501768 358316 502396 358412
rect 501768 357324 501864 358316
rect 560794 357868 560890 358860
rect 560632 357772 560890 357868
rect 501768 357228 502396 357324
rect 501768 356236 501864 357228
rect 560794 356780 560890 357772
rect 560632 356684 560890 356780
rect 501768 356140 502396 356236
rect 501768 355148 501864 356140
rect 560794 355692 560890 356684
rect 560632 355596 560890 355692
rect 501768 355052 502396 355148
rect 501768 354060 501864 355052
rect 560794 354604 560890 355596
rect 560632 354508 560890 354604
rect 501768 353964 502396 354060
rect 501768 352972 501864 353964
rect 560794 353516 560890 354508
rect 560632 353420 560890 353516
rect 501768 352876 502396 352972
rect 501768 351884 501864 352876
rect 560794 352428 560890 353420
rect 560632 352332 560890 352428
rect 501768 351788 502396 351884
rect 501768 350796 501864 351788
rect 560794 351340 560890 352332
rect 560632 351244 560890 351340
rect 501768 350700 502396 350796
rect 501768 349708 501864 350700
rect 560794 350252 560890 351244
rect 560632 350156 560890 350252
rect 501768 349612 502396 349708
rect 501768 348620 501864 349612
rect 560794 349164 560890 350156
rect 560632 349068 560890 349164
rect 501768 348524 502396 348620
rect 501768 347532 501864 348524
rect 560794 348076 560890 349068
rect 560632 347980 560890 348076
rect 501768 347436 502396 347532
rect 501768 346444 501864 347436
rect 560794 346988 560890 347980
rect 560632 346892 560890 346988
rect 501768 346348 502396 346444
rect 501768 345356 501864 346348
rect 560794 345900 560890 346892
rect 560632 345804 560890 345900
rect 501768 345260 502396 345356
rect 501768 344268 501864 345260
rect 560794 344812 560890 345804
rect 560632 344716 560890 344812
rect 501768 344172 502396 344268
rect 501768 343180 501864 344172
rect 560794 343724 560890 344716
rect 560632 343628 560890 343724
rect 501768 343084 502396 343180
rect 501768 342997 501864 343084
rect 437262 341992 437358 342984
rect 496288 342949 501864 342997
rect 496288 342536 498496 342949
rect 495756 342440 498496 342536
rect 496288 342021 498496 342440
rect 499520 342092 501864 342949
rect 560794 342997 560890 343628
rect 560794 342949 566821 342997
rect 560794 342636 564289 342949
rect 560632 342540 564289 342636
rect 499520 342021 502396 342092
rect 496288 341996 502396 342021
rect 560794 342021 564289 342540
rect 565313 342021 566821 342949
rect 437262 341896 437520 341992
rect 496288 341973 501864 341996
rect 437262 340904 437358 341896
rect 496288 341448 496384 341973
rect 495756 341352 496384 341448
rect 436432 340883 437075 340889
rect 437262 340883 437520 340904
rect 436432 340882 437520 340883
rect 435474 340835 437520 340882
rect 435474 340460 436583 340835
rect 435312 340364 436583 340460
rect 435474 340163 436583 340364
rect 437273 340808 437520 340835
rect 437273 340163 437358 340808
rect 496288 340360 496384 341352
rect 495756 340264 496384 340360
rect 435474 340091 437358 340163
rect 435474 340078 437075 340091
rect 435474 340074 436468 340078
rect 376448 339820 377076 339916
rect 376448 338828 376544 339820
rect 435474 339372 435570 340074
rect 435312 339276 435570 339372
rect 376448 338732 377076 338828
rect 376448 337740 376544 338732
rect 435474 338284 435570 339276
rect 435312 338188 435570 338284
rect 376448 337644 377076 337740
rect 376448 336652 376544 337644
rect 435474 337196 435570 338188
rect 435312 337100 435570 337196
rect 376448 336556 377076 336652
rect 376448 335564 376544 336556
rect 435474 336108 435570 337100
rect 435312 336012 435570 336108
rect 376448 335468 377076 335564
rect 376448 334476 376544 335468
rect 435474 335020 435570 336012
rect 435312 334924 435570 335020
rect 376448 334380 377076 334476
rect 376448 333388 376544 334380
rect 435474 333932 435570 334924
rect 435312 333836 435570 333932
rect 376448 333292 377076 333388
rect 376448 332300 376544 333292
rect 435474 332844 435570 333836
rect 435312 332748 435570 332844
rect 376448 332204 377076 332300
rect 376448 331212 376544 332204
rect 435474 331756 435570 332748
rect 435312 331660 435570 331756
rect 376448 331116 377076 331212
rect 376448 330124 376544 331116
rect 435474 330668 435570 331660
rect 435312 330572 435570 330668
rect 376448 330028 377076 330124
rect 376448 329036 376544 330028
rect 435474 329580 435570 330572
rect 435312 329484 435570 329580
rect 376448 328940 377076 329036
rect 376448 327948 376544 328940
rect 435474 328492 435570 329484
rect 435312 328396 435570 328492
rect 376448 327852 377076 327948
rect 376448 326860 376544 327852
rect 435474 327404 435570 328396
rect 435312 327308 435570 327404
rect 376448 326764 377076 326860
rect 376448 325772 376544 326764
rect 435474 326316 435570 327308
rect 435312 326220 435570 326316
rect 376448 325676 377076 325772
rect 376448 324684 376544 325676
rect 435474 325228 435570 326220
rect 435312 325132 435570 325228
rect 376448 324588 377076 324684
rect 376448 323596 376544 324588
rect 435474 324140 435570 325132
rect 435312 324044 435570 324140
rect 376448 323500 377076 323596
rect 376448 322508 376544 323500
rect 435474 323052 435570 324044
rect 435312 322956 435570 323052
rect 376448 322412 377076 322508
rect 376448 321420 376544 322412
rect 435474 321964 435570 322956
rect 435312 321868 435570 321964
rect 376448 321324 377076 321420
rect 376448 320332 376544 321324
rect 435474 320876 435570 321868
rect 435312 320780 435570 320876
rect 376448 320236 377076 320332
rect 376448 319244 376544 320236
rect 435474 319788 435570 320780
rect 435312 319692 435570 319788
rect 376448 319148 377076 319244
rect 376448 318156 376544 319148
rect 435474 318700 435570 319692
rect 435312 318604 435570 318700
rect 376448 318060 377076 318156
rect 376448 317068 376544 318060
rect 435474 317612 435570 318604
rect 435312 317516 435570 317612
rect 376448 316972 377076 317068
rect 376448 315983 376544 316972
rect 435474 316524 435570 317516
rect 435312 316428 435570 316524
rect 375661 315980 376544 315983
rect 435474 316294 435570 316428
rect 437262 339816 437358 340091
rect 437262 339720 437520 339816
rect 437262 338728 437358 339720
rect 496288 339272 496384 340264
rect 495756 339176 496384 339272
rect 437262 338632 437520 338728
rect 437262 337640 437358 338632
rect 496288 338184 496384 339176
rect 495756 338088 496384 338184
rect 437262 337544 437520 337640
rect 437262 336552 437358 337544
rect 496288 337096 496384 338088
rect 495756 337000 496384 337096
rect 437262 336456 437520 336552
rect 437262 335464 437358 336456
rect 496288 336008 496384 337000
rect 495756 335912 496384 336008
rect 437262 335368 437520 335464
rect 437262 334376 437358 335368
rect 496288 334920 496384 335912
rect 495756 334824 496384 334920
rect 437262 334280 437520 334376
rect 437262 333288 437358 334280
rect 496288 333832 496384 334824
rect 495756 333736 496384 333832
rect 437262 333192 437520 333288
rect 437262 332200 437358 333192
rect 496288 332744 496384 333736
rect 495756 332648 496384 332744
rect 437262 332104 437520 332200
rect 437262 331112 437358 332104
rect 496288 331656 496384 332648
rect 495756 331560 496384 331656
rect 437262 331016 437520 331112
rect 437262 330024 437358 331016
rect 496288 330568 496384 331560
rect 495756 330472 496384 330568
rect 437262 329928 437520 330024
rect 437262 328936 437358 329928
rect 496288 329480 496384 330472
rect 495756 329384 496384 329480
rect 437262 328840 437520 328936
rect 437262 327848 437358 328840
rect 496288 328392 496384 329384
rect 495756 328296 496384 328392
rect 437262 327752 437520 327848
rect 437262 326760 437358 327752
rect 496288 327304 496384 328296
rect 495756 327208 496384 327304
rect 437262 326664 437520 326760
rect 437262 325672 437358 326664
rect 496288 326216 496384 327208
rect 495756 326120 496384 326216
rect 437262 325576 437520 325672
rect 437262 324584 437358 325576
rect 496288 325128 496384 326120
rect 495756 325032 496384 325128
rect 437262 324488 437520 324584
rect 437262 323496 437358 324488
rect 496288 324040 496384 325032
rect 495756 323944 496384 324040
rect 437262 323400 437520 323496
rect 437262 322408 437358 323400
rect 496288 322952 496384 323944
rect 495756 322856 496384 322952
rect 437262 322312 437520 322408
rect 437262 321320 437358 322312
rect 496288 321864 496384 322856
rect 495756 321768 496384 321864
rect 437262 321224 437520 321320
rect 437262 320232 437358 321224
rect 496288 320776 496384 321768
rect 495756 320680 496384 320776
rect 437262 320136 437520 320232
rect 437262 319144 437358 320136
rect 496288 319688 496384 320680
rect 495756 319592 496384 319688
rect 437262 319048 437520 319144
rect 437262 318056 437358 319048
rect 496288 318600 496384 319592
rect 495756 318504 496384 318600
rect 437262 317960 437520 318056
rect 437262 316968 437358 317960
rect 496288 317512 496384 318504
rect 495756 317416 496384 317512
rect 437262 316872 437616 316968
rect 375661 315887 377076 315980
rect 370340 315325 371850 315336
rect 370340 315240 371851 315325
rect 309869 310888 309915 310899
rect 311944 315035 312040 315047
rect 311944 310884 312040 314939
rect 311944 310788 312200 310884
rect 311944 309930 312038 310788
rect 370436 310337 371064 310340
rect 371755 310337 371851 315240
rect 375661 310984 375757 315887
rect 376448 315884 377076 315887
rect 435474 315436 435568 316294
rect 437262 316083 437358 316872
rect 496288 316424 496384 317416
rect 495756 316328 496384 316424
rect 437264 315959 437358 316083
rect 437252 315863 437258 315959
rect 437366 315880 437372 315959
rect 437366 315863 437616 315880
rect 437264 315784 437616 315863
rect 437264 315444 437358 315472
rect 435312 315340 435568 315436
rect 435472 311285 435568 315340
rect 496288 315336 496384 316328
rect 501768 341004 501864 341973
rect 560794 341973 566821 342021
rect 560794 341548 560890 341973
rect 560632 341452 560890 341548
rect 501768 340908 502396 341004
rect 501768 339916 501864 340908
rect 560794 340460 560890 341452
rect 560632 340364 560890 340460
rect 501768 339820 502396 339916
rect 501768 338828 501864 339820
rect 560794 339372 560890 340364
rect 560632 339276 560890 339372
rect 501768 338732 502396 338828
rect 501768 337740 501864 338732
rect 560794 338284 560890 339276
rect 560632 338188 560890 338284
rect 501768 337644 502396 337740
rect 501768 336652 501864 337644
rect 560794 337196 560890 338188
rect 560632 337100 560890 337196
rect 501768 336556 502396 336652
rect 501768 335564 501864 336556
rect 560794 336108 560890 337100
rect 560632 336012 560890 336108
rect 501768 335468 502396 335564
rect 501768 334476 501864 335468
rect 560794 335020 560890 336012
rect 560632 334924 560890 335020
rect 501768 334380 502396 334476
rect 501768 333388 501864 334380
rect 560794 333932 560890 334924
rect 560632 333836 560890 333932
rect 501768 333292 502396 333388
rect 501768 332300 501864 333292
rect 560794 332844 560890 333836
rect 560632 332748 560890 332844
rect 501768 332204 502396 332300
rect 501768 331212 501864 332204
rect 560794 331756 560890 332748
rect 560632 331660 560890 331756
rect 501768 331116 502396 331212
rect 501768 330124 501864 331116
rect 560794 330668 560890 331660
rect 560632 330572 560890 330668
rect 501768 330028 502396 330124
rect 501768 329036 501864 330028
rect 560794 329580 560890 330572
rect 560632 329484 560890 329580
rect 501768 328940 502396 329036
rect 501768 327948 501864 328940
rect 560794 328492 560890 329484
rect 560632 328396 560890 328492
rect 501768 327852 502396 327948
rect 501768 326860 501864 327852
rect 560794 327404 560890 328396
rect 560632 327308 560890 327404
rect 501768 326764 502396 326860
rect 501768 325772 501864 326764
rect 560794 326316 560890 327308
rect 560632 326220 560890 326316
rect 501768 325676 502396 325772
rect 501768 324684 501864 325676
rect 560794 325228 560890 326220
rect 560632 325132 560890 325228
rect 501768 324588 502396 324684
rect 501768 323596 501864 324588
rect 560794 324140 560890 325132
rect 560632 324044 560890 324140
rect 501768 323500 502396 323596
rect 501768 322508 501864 323500
rect 560794 323052 560890 324044
rect 560632 322956 560890 323052
rect 501768 322412 502396 322508
rect 501768 321420 501864 322412
rect 560794 321964 560890 322956
rect 560632 321868 560890 321964
rect 501768 321324 502396 321420
rect 501768 320332 501864 321324
rect 560794 320876 560890 321868
rect 560632 320780 560890 320876
rect 501768 320236 502396 320332
rect 501768 319244 501864 320236
rect 560794 319788 560890 320780
rect 560632 319692 560890 319788
rect 501768 319148 502396 319244
rect 501768 318156 501864 319148
rect 560794 318700 560890 319692
rect 560632 318604 560890 318700
rect 501768 318060 502396 318156
rect 501768 317068 501864 318060
rect 560794 317612 560890 318604
rect 560632 317516 560890 317612
rect 501768 316972 502396 317068
rect 501768 315983 501864 316972
rect 560794 316524 560890 317516
rect 560632 316428 560890 316524
rect 500981 315980 501864 315983
rect 560794 316294 560890 316428
rect 500981 315887 502396 315980
rect 495660 315325 497170 315336
rect 495660 315240 497171 315325
rect 435472 311177 435568 311189
rect 437264 315035 437360 315047
rect 375661 310899 377172 310984
rect 375662 310888 377172 310899
rect 370436 310244 371851 310337
rect 311942 309796 312038 309930
rect 370968 310241 371851 310244
rect 311942 309700 312200 309796
rect 311942 308708 312038 309700
rect 370968 309252 371064 310241
rect 370436 309156 371064 309252
rect 311942 308612 312200 308708
rect 311942 307620 312038 308612
rect 370968 308164 371064 309156
rect 370436 308068 371064 308164
rect 311942 307524 312200 307620
rect 311942 306532 312038 307524
rect 370968 307076 371064 308068
rect 370436 306980 371064 307076
rect 311942 306436 312200 306532
rect 311942 305444 312038 306436
rect 370968 305988 371064 306980
rect 370436 305892 371064 305988
rect 311942 305348 312200 305444
rect 311942 304356 312038 305348
rect 370968 304900 371064 305892
rect 370436 304804 371064 304900
rect 311942 304260 312200 304356
rect 311942 303268 312038 304260
rect 370968 303812 371064 304804
rect 370436 303716 371064 303812
rect 311942 303172 312200 303268
rect 311942 302180 312038 303172
rect 370968 302724 371064 303716
rect 370436 302628 371064 302724
rect 311942 302084 312200 302180
rect 311942 301092 312038 302084
rect 370968 301636 371064 302628
rect 370436 301540 371064 301636
rect 311942 300996 312200 301092
rect 311942 300004 312038 300996
rect 370968 300548 371064 301540
rect 370436 300452 371064 300548
rect 311942 299908 312200 300004
rect 311942 298916 312038 299908
rect 370968 299460 371064 300452
rect 370436 299364 371064 299460
rect 311942 298820 312200 298916
rect 311942 297828 312038 298820
rect 370968 298372 371064 299364
rect 370436 298276 371064 298372
rect 311942 297732 312200 297828
rect 311942 296740 312038 297732
rect 370968 297284 371064 298276
rect 370436 297188 371064 297284
rect 311942 296644 312200 296740
rect 311942 295652 312038 296644
rect 370968 296196 371064 297188
rect 370436 296100 371064 296196
rect 311942 295556 312200 295652
rect 311942 294564 312038 295556
rect 370968 295108 371064 296100
rect 370436 295012 371064 295108
rect 311942 294468 312200 294564
rect 311942 293476 312038 294468
rect 370968 294020 371064 295012
rect 370436 293924 371064 294020
rect 311942 293380 312200 293476
rect 311942 292388 312038 293380
rect 370968 292932 371064 293924
rect 370436 292836 371064 292932
rect 311942 292292 312200 292388
rect 311942 291300 312038 292292
rect 370968 291844 371064 292836
rect 370436 291748 371064 291844
rect 311942 291204 312200 291300
rect 311942 290212 312038 291204
rect 370968 290756 371064 291748
rect 370436 290660 371064 290756
rect 311942 290116 312200 290212
rect 311942 289124 312038 290116
rect 370968 289668 371064 290660
rect 370436 289572 371064 289668
rect 311942 289028 312200 289124
rect 311942 288036 312038 289028
rect 370968 288580 371064 289572
rect 370436 288484 371064 288580
rect 311942 287940 312200 288036
rect 311942 286948 312038 287940
rect 370968 287492 371064 288484
rect 370436 287396 371064 287492
rect 311942 286852 312200 286948
rect 311942 285860 312038 286852
rect 370968 286404 371064 287396
rect 370436 286308 371064 286404
rect 311942 285764 312200 285860
rect 311942 284772 312038 285764
rect 370968 285316 371064 286308
rect 370436 285220 371064 285316
rect 311942 284676 312200 284772
rect 311942 283684 312038 284676
rect 370968 284228 371064 285220
rect 370436 284132 371064 284228
rect 311942 283588 312200 283684
rect 311942 282596 312038 283588
rect 370968 283140 371064 284132
rect 370436 283044 371064 283140
rect 311942 282500 312200 282596
rect 311942 281508 312038 282500
rect 370968 282052 371064 283044
rect 370436 281956 371064 282052
rect 311942 281412 312200 281508
rect 311942 280420 312038 281412
rect 370968 280964 371064 281956
rect 370436 280868 371064 280964
rect 311942 280337 312200 280420
rect 306149 280324 312200 280337
rect 370968 280337 371064 280868
rect 376448 309896 376544 310888
rect 437264 310884 437360 314939
rect 437264 310788 437520 310884
rect 435474 310752 435568 310780
rect 435216 310361 435568 310440
rect 435216 310344 435466 310361
rect 435460 310265 435466 310344
rect 435574 310265 435580 310361
rect 435474 310141 435568 310265
rect 376448 309800 377076 309896
rect 376448 308808 376544 309800
rect 435474 309352 435570 310141
rect 437264 309930 437358 310788
rect 495756 310337 496384 310340
rect 497075 310337 497171 315240
rect 500981 310984 501077 315887
rect 501768 315884 502396 315887
rect 560794 315436 560888 316294
rect 560632 315340 560888 315436
rect 560792 311285 560888 315340
rect 560792 311177 560888 311189
rect 500981 310899 502492 310984
rect 566774 310899 566821 315983
rect 500982 310888 502492 310899
rect 566775 310888 566821 310899
rect 495756 310244 497171 310337
rect 435216 309256 435570 309352
rect 376448 308712 377076 308808
rect 376448 307720 376544 308712
rect 435474 308264 435570 309256
rect 435312 308168 435570 308264
rect 376448 307624 377076 307720
rect 376448 306632 376544 307624
rect 435474 307176 435570 308168
rect 435312 307080 435570 307176
rect 376448 306536 377076 306632
rect 376448 305544 376544 306536
rect 435474 306088 435570 307080
rect 435312 305992 435570 306088
rect 376448 305448 377076 305544
rect 376448 304456 376544 305448
rect 435474 305000 435570 305992
rect 435312 304904 435570 305000
rect 376448 304360 377076 304456
rect 376448 303368 376544 304360
rect 435474 303912 435570 304904
rect 435312 303816 435570 303912
rect 376448 303272 377076 303368
rect 376448 302280 376544 303272
rect 435474 302824 435570 303816
rect 435312 302728 435570 302824
rect 376448 302184 377076 302280
rect 376448 301192 376544 302184
rect 435474 301736 435570 302728
rect 435312 301640 435570 301736
rect 376448 301096 377076 301192
rect 376448 300104 376544 301096
rect 435474 300648 435570 301640
rect 435312 300552 435570 300648
rect 376448 300008 377076 300104
rect 376448 299016 376544 300008
rect 435474 299560 435570 300552
rect 435312 299464 435570 299560
rect 376448 298920 377076 299016
rect 376448 297928 376544 298920
rect 435474 298472 435570 299464
rect 435312 298376 435570 298472
rect 376448 297832 377076 297928
rect 376448 296840 376544 297832
rect 435474 297384 435570 298376
rect 435312 297288 435570 297384
rect 376448 296744 377076 296840
rect 376448 295752 376544 296744
rect 435474 296296 435570 297288
rect 435312 296200 435570 296296
rect 376448 295656 377076 295752
rect 376448 294664 376544 295656
rect 435474 295208 435570 296200
rect 435312 295112 435570 295208
rect 376448 294568 377076 294664
rect 376448 293576 376544 294568
rect 435474 294120 435570 295112
rect 435312 294024 435570 294120
rect 376448 293480 377076 293576
rect 376448 292488 376544 293480
rect 435474 293032 435570 294024
rect 435312 292936 435570 293032
rect 376448 292392 377076 292488
rect 376448 291400 376544 292392
rect 435474 291944 435570 292936
rect 435312 291848 435570 291944
rect 376448 291304 377076 291400
rect 376448 290312 376544 291304
rect 435474 290856 435570 291848
rect 435312 290760 435570 290856
rect 376448 290216 377076 290312
rect 376448 289224 376544 290216
rect 435474 289768 435570 290760
rect 435312 289672 435570 289768
rect 376448 289128 377076 289224
rect 376448 288136 376544 289128
rect 435474 288680 435570 289672
rect 435312 288584 435570 288680
rect 376448 288040 377076 288136
rect 376448 287048 376544 288040
rect 435474 287592 435570 288584
rect 435312 287496 435570 287592
rect 376448 286952 377076 287048
rect 376448 285960 376544 286952
rect 435474 286504 435570 287496
rect 435312 286408 435570 286504
rect 376448 285864 377076 285960
rect 376448 284872 376544 285864
rect 435474 285416 435570 286408
rect 435312 285320 435570 285416
rect 376448 284776 377076 284872
rect 376448 283784 376544 284776
rect 435474 284328 435570 285320
rect 435312 284232 435570 284328
rect 376448 283688 377076 283784
rect 376448 282696 376544 283688
rect 435474 283240 435570 284232
rect 435312 283144 435570 283240
rect 376448 282600 377076 282696
rect 376448 281608 376544 282600
rect 435474 282152 435570 283144
rect 435312 282056 435570 282152
rect 376448 281512 377076 281608
rect 376448 280520 376544 281512
rect 435474 281064 435570 282056
rect 435312 280968 435570 281064
rect 376448 280424 377076 280520
rect 376448 280337 376544 280424
rect 306149 280289 312038 280324
rect 306149 279361 307383 280289
rect 308407 279361 312038 280289
rect 370968 280289 376544 280337
rect 370968 279876 373176 280289
rect 370436 279780 373176 279876
rect 306149 279332 312038 279361
rect 370968 279361 373176 279780
rect 374200 279432 376544 280289
rect 435474 279976 435570 280968
rect 435312 279880 435570 279976
rect 374200 279361 377076 279432
rect 370968 279336 377076 279361
rect 306149 279313 312200 279332
rect 311942 279236 312200 279313
rect 370968 279313 376544 279336
rect 311942 278244 312038 279236
rect 370968 278788 371064 279313
rect 370436 278692 371064 278788
rect 311942 278148 312200 278244
rect 311942 277156 312038 278148
rect 370968 277700 371064 278692
rect 370436 277604 371064 277700
rect 311942 277060 312200 277156
rect 311942 276068 312038 277060
rect 370968 276612 371064 277604
rect 370436 276516 371064 276612
rect 311942 275972 312200 276068
rect 311942 274980 312038 275972
rect 370968 275524 371064 276516
rect 370436 275428 371064 275524
rect 311942 274884 312200 274980
rect 311942 273892 312038 274884
rect 370968 274436 371064 275428
rect 370436 274340 371064 274436
rect 311942 273796 312200 273892
rect 311942 272804 312038 273796
rect 370968 273348 371064 274340
rect 370436 273252 371064 273348
rect 311942 272708 312200 272804
rect 311942 271716 312038 272708
rect 370968 272260 371064 273252
rect 370436 272164 371064 272260
rect 311942 271620 312200 271716
rect 311942 270628 312038 271620
rect 370968 271172 371064 272164
rect 370436 271076 371064 271172
rect 311942 270532 312200 270628
rect 311942 269540 312038 270532
rect 370968 270084 371064 271076
rect 370436 269988 371064 270084
rect 311942 269444 312200 269540
rect 311942 268452 312038 269444
rect 370968 268996 371064 269988
rect 370436 268900 371064 268996
rect 311942 268356 312200 268452
rect 311942 267364 312038 268356
rect 370968 267908 371064 268900
rect 370436 267812 371064 267908
rect 311942 267268 312200 267364
rect 311942 266276 312038 267268
rect 370968 266820 371064 267812
rect 370436 266724 371064 266820
rect 311942 266180 312200 266276
rect 311942 265188 312038 266180
rect 370968 265732 371064 266724
rect 370436 265636 371064 265732
rect 311942 265092 312200 265188
rect 311942 264100 312038 265092
rect 370968 264644 371064 265636
rect 370436 264548 371064 264644
rect 311942 264004 312200 264100
rect 311942 263012 312038 264004
rect 370968 263556 371064 264548
rect 370436 263460 371064 263556
rect 311942 262916 312200 263012
rect 311942 261924 312038 262916
rect 370968 262468 371064 263460
rect 370436 262372 371064 262468
rect 311942 261828 312200 261924
rect 311942 260836 312038 261828
rect 370968 261380 371064 262372
rect 370436 261284 371064 261380
rect 311942 260740 312200 260836
rect 311942 259748 312038 260740
rect 370968 260292 371064 261284
rect 370436 260196 371064 260292
rect 311942 259652 312200 259748
rect 311942 258660 312038 259652
rect 370968 259204 371064 260196
rect 370436 259108 371064 259204
rect 311942 258564 312200 258660
rect 311942 257572 312038 258564
rect 370968 258116 371064 259108
rect 370436 258020 371064 258116
rect 311942 257476 312200 257572
rect 311942 256484 312038 257476
rect 370968 257028 371064 258020
rect 370436 256932 371064 257028
rect 311942 256388 312200 256484
rect 311942 255396 312038 256388
rect 370968 255940 371064 256932
rect 370436 255844 371064 255940
rect 311942 255300 312200 255396
rect 311942 254308 312038 255300
rect 370968 254852 371064 255844
rect 370436 254756 371064 254852
rect 311942 254212 312296 254308
rect 309839 248228 309915 253320
rect 311942 253220 312038 254212
rect 370968 253764 371064 254756
rect 370436 253668 371064 253764
rect 311942 253217 312296 253220
rect 311936 253121 311942 253217
rect 312038 253124 312296 253217
rect 312038 253121 312044 253124
rect 370968 252676 371064 253668
rect 376448 278344 376544 279313
rect 435474 278888 435570 279880
rect 435312 278792 435570 278888
rect 376448 278248 377076 278344
rect 376448 277256 376544 278248
rect 435474 278228 435570 278792
rect 437262 309796 437358 309930
rect 496288 310241 497171 310244
rect 437262 309700 437520 309796
rect 437262 308708 437358 309700
rect 496288 309252 496384 310241
rect 495756 309156 496384 309252
rect 437262 308612 437520 308708
rect 437262 307620 437358 308612
rect 496288 308164 496384 309156
rect 495756 308068 496384 308164
rect 437262 307524 437520 307620
rect 437262 306532 437358 307524
rect 496288 307076 496384 308068
rect 495756 306980 496384 307076
rect 437262 306436 437520 306532
rect 437262 305444 437358 306436
rect 496288 305988 496384 306980
rect 495756 305892 496384 305988
rect 437262 305348 437520 305444
rect 437262 304356 437358 305348
rect 496288 304900 496384 305892
rect 495756 304804 496384 304900
rect 437262 304260 437520 304356
rect 437262 303268 437358 304260
rect 496288 303812 496384 304804
rect 495756 303716 496384 303812
rect 437262 303172 437520 303268
rect 437262 302180 437358 303172
rect 496288 302724 496384 303716
rect 495756 302628 496384 302724
rect 437262 302084 437520 302180
rect 437262 301092 437358 302084
rect 496288 301636 496384 302628
rect 495756 301540 496384 301636
rect 437262 300996 437520 301092
rect 437262 300004 437358 300996
rect 496288 300548 496384 301540
rect 495756 300452 496384 300548
rect 437262 299908 437520 300004
rect 437262 298916 437358 299908
rect 496288 299460 496384 300452
rect 495756 299364 496384 299460
rect 437262 298820 437520 298916
rect 437262 297828 437358 298820
rect 496288 298372 496384 299364
rect 495756 298276 496384 298372
rect 437262 297732 437520 297828
rect 437262 296740 437358 297732
rect 496288 297284 496384 298276
rect 495756 297188 496384 297284
rect 437262 296644 437520 296740
rect 437262 295652 437358 296644
rect 496288 296196 496384 297188
rect 495756 296100 496384 296196
rect 437262 295556 437520 295652
rect 437262 294564 437358 295556
rect 496288 295108 496384 296100
rect 495756 295012 496384 295108
rect 437262 294468 437520 294564
rect 437262 293476 437358 294468
rect 496288 294020 496384 295012
rect 495756 293924 496384 294020
rect 437262 293380 437520 293476
rect 437262 292388 437358 293380
rect 496288 292932 496384 293924
rect 495756 292836 496384 292932
rect 437262 292292 437520 292388
rect 437262 291300 437358 292292
rect 496288 291844 496384 292836
rect 495756 291748 496384 291844
rect 437262 291204 437520 291300
rect 437262 290212 437358 291204
rect 496288 290756 496384 291748
rect 495756 290660 496384 290756
rect 437262 290116 437520 290212
rect 437262 289124 437358 290116
rect 496288 289668 496384 290660
rect 495756 289572 496384 289668
rect 437262 289028 437520 289124
rect 437262 288036 437358 289028
rect 496288 288580 496384 289572
rect 495756 288484 496384 288580
rect 437262 287940 437520 288036
rect 437262 286948 437358 287940
rect 496288 287492 496384 288484
rect 495756 287396 496384 287492
rect 437262 286852 437520 286948
rect 437262 285860 437358 286852
rect 496288 286404 496384 287396
rect 495756 286308 496384 286404
rect 437262 285764 437520 285860
rect 437262 284772 437358 285764
rect 496288 285316 496384 286308
rect 495756 285220 496384 285316
rect 437262 284676 437520 284772
rect 437262 283684 437358 284676
rect 496288 284228 496384 285220
rect 495756 284132 496384 284228
rect 437262 283588 437520 283684
rect 437262 282596 437358 283588
rect 496288 283140 496384 284132
rect 495756 283044 496384 283140
rect 437262 282500 437520 282596
rect 437262 281508 437358 282500
rect 496288 282052 496384 283044
rect 495756 281956 496384 282052
rect 437262 281412 437520 281508
rect 437262 280420 437358 281412
rect 496288 280964 496384 281956
rect 495756 280868 496384 280964
rect 437262 280324 437520 280420
rect 496288 280337 496384 280868
rect 501768 309896 501864 310888
rect 560794 310752 560888 310780
rect 560536 310361 560888 310440
rect 560536 310344 560786 310361
rect 560780 310265 560786 310344
rect 560894 310265 560900 310361
rect 560794 310141 560888 310265
rect 501768 309800 502396 309896
rect 501768 308808 501864 309800
rect 560794 309352 560890 310141
rect 560536 309256 560890 309352
rect 501768 308712 502396 308808
rect 501768 307720 501864 308712
rect 560794 308264 560890 309256
rect 560632 308168 560890 308264
rect 501768 307624 502396 307720
rect 501768 306632 501864 307624
rect 560794 307176 560890 308168
rect 560632 307080 560890 307176
rect 501768 306536 502396 306632
rect 501768 305544 501864 306536
rect 560794 306088 560890 307080
rect 560632 305992 560890 306088
rect 501768 305448 502396 305544
rect 501768 304456 501864 305448
rect 560794 305000 560890 305992
rect 560632 304904 560890 305000
rect 501768 304360 502396 304456
rect 501768 303368 501864 304360
rect 560794 303912 560890 304904
rect 560632 303816 560890 303912
rect 501768 303272 502396 303368
rect 501768 302280 501864 303272
rect 560794 302824 560890 303816
rect 560632 302728 560890 302824
rect 501768 302184 502396 302280
rect 501768 301192 501864 302184
rect 560794 301736 560890 302728
rect 560632 301640 560890 301736
rect 501768 301096 502396 301192
rect 501768 300104 501864 301096
rect 560794 300648 560890 301640
rect 560632 300552 560890 300648
rect 501768 300008 502396 300104
rect 501768 299016 501864 300008
rect 560794 299560 560890 300552
rect 560632 299464 560890 299560
rect 501768 298920 502396 299016
rect 501768 297928 501864 298920
rect 560794 298472 560890 299464
rect 560632 298376 560890 298472
rect 501768 297832 502396 297928
rect 501768 296840 501864 297832
rect 560794 297384 560890 298376
rect 560632 297288 560890 297384
rect 501768 296744 502396 296840
rect 501768 295752 501864 296744
rect 560794 296296 560890 297288
rect 560632 296200 560890 296296
rect 501768 295656 502396 295752
rect 501768 294664 501864 295656
rect 560794 295208 560890 296200
rect 560632 295112 560890 295208
rect 501768 294568 502396 294664
rect 501768 293576 501864 294568
rect 560794 294120 560890 295112
rect 560632 294024 560890 294120
rect 501768 293480 502396 293576
rect 501768 292488 501864 293480
rect 560794 293032 560890 294024
rect 560632 292936 560890 293032
rect 501768 292392 502396 292488
rect 501768 291400 501864 292392
rect 560794 291944 560890 292936
rect 560632 291848 560890 291944
rect 501768 291304 502396 291400
rect 501768 290312 501864 291304
rect 560794 290856 560890 291848
rect 560632 290760 560890 290856
rect 501768 290216 502396 290312
rect 501768 289224 501864 290216
rect 560794 289768 560890 290760
rect 560632 289672 560890 289768
rect 501768 289128 502396 289224
rect 501768 288136 501864 289128
rect 560794 288680 560890 289672
rect 560632 288584 560890 288680
rect 501768 288040 502396 288136
rect 501768 287048 501864 288040
rect 560794 287592 560890 288584
rect 560632 287496 560890 287592
rect 501768 286952 502396 287048
rect 501768 285960 501864 286952
rect 560794 286504 560890 287496
rect 560632 286408 560890 286504
rect 501768 285864 502396 285960
rect 501768 284872 501864 285864
rect 560794 285416 560890 286408
rect 560632 285320 560890 285416
rect 501768 284776 502396 284872
rect 501768 283784 501864 284776
rect 560794 284328 560890 285320
rect 560632 284232 560890 284328
rect 501768 283688 502396 283784
rect 501768 282696 501864 283688
rect 560794 283240 560890 284232
rect 560632 283144 560890 283240
rect 501768 282600 502396 282696
rect 501768 281608 501864 282600
rect 560794 282152 560890 283144
rect 560632 282056 560890 282152
rect 501768 281512 502396 281608
rect 501768 280520 501864 281512
rect 560794 281064 560890 282056
rect 560632 280968 560890 281064
rect 501768 280424 502396 280520
rect 501768 280337 501864 280424
rect 437262 279332 437358 280324
rect 496288 280289 501864 280337
rect 496288 279876 498496 280289
rect 495756 279780 498496 279876
rect 496288 279361 498496 279780
rect 499520 279432 501864 280289
rect 560794 280337 560890 280968
rect 560794 280289 566821 280337
rect 560794 279976 564289 280289
rect 560632 279880 564289 279976
rect 499520 279361 502396 279432
rect 496288 279336 502396 279361
rect 560794 279361 564289 279880
rect 565313 279361 566821 280289
rect 437262 279236 437520 279332
rect 496288 279313 501864 279336
rect 437262 278244 437358 279236
rect 496288 278788 496384 279313
rect 495756 278692 496384 278788
rect 436432 278228 437075 278229
rect 435474 278223 437075 278228
rect 437262 278223 437520 278244
rect 435474 278175 437520 278223
rect 435474 277800 436583 278175
rect 435312 277704 436583 277800
rect 435474 277503 436583 277704
rect 437273 278148 437520 278175
rect 437273 277503 437358 278148
rect 496288 277700 496384 278692
rect 495756 277604 496384 277700
rect 435474 277431 437358 277503
rect 435474 277420 437075 277431
rect 376448 277160 377076 277256
rect 376448 276168 376544 277160
rect 435474 276712 435570 277420
rect 436432 277418 437075 277420
rect 435312 276616 435570 276712
rect 376448 276072 377076 276168
rect 376448 275080 376544 276072
rect 435474 275624 435570 276616
rect 435312 275528 435570 275624
rect 376448 274984 377076 275080
rect 376448 273992 376544 274984
rect 435474 274536 435570 275528
rect 435312 274440 435570 274536
rect 376448 273896 377076 273992
rect 376448 272904 376544 273896
rect 435474 273448 435570 274440
rect 435312 273352 435570 273448
rect 376448 272808 377076 272904
rect 376448 271816 376544 272808
rect 435474 272360 435570 273352
rect 435312 272264 435570 272360
rect 376448 271720 377076 271816
rect 376448 270728 376544 271720
rect 435474 271272 435570 272264
rect 435312 271176 435570 271272
rect 376448 270632 377076 270728
rect 376448 269640 376544 270632
rect 435474 270184 435570 271176
rect 435312 270088 435570 270184
rect 376448 269544 377076 269640
rect 376448 268552 376544 269544
rect 435474 269096 435570 270088
rect 435312 269000 435570 269096
rect 376448 268456 377076 268552
rect 376448 267464 376544 268456
rect 435474 268008 435570 269000
rect 435312 267912 435570 268008
rect 376448 267368 377076 267464
rect 376448 266376 376544 267368
rect 435474 266920 435570 267912
rect 435312 266824 435570 266920
rect 376448 266280 377076 266376
rect 376448 265288 376544 266280
rect 435474 265832 435570 266824
rect 435312 265736 435570 265832
rect 376448 265192 377076 265288
rect 376448 264200 376544 265192
rect 435474 264744 435570 265736
rect 435312 264648 435570 264744
rect 376448 264104 377076 264200
rect 376448 263112 376544 264104
rect 435474 263656 435570 264648
rect 435312 263560 435570 263656
rect 376448 263016 377076 263112
rect 376448 262024 376544 263016
rect 435474 262568 435570 263560
rect 435312 262472 435570 262568
rect 376448 261928 377076 262024
rect 376448 260936 376544 261928
rect 435474 261480 435570 262472
rect 435312 261384 435570 261480
rect 376448 260840 377076 260936
rect 376448 259848 376544 260840
rect 435474 260392 435570 261384
rect 435312 260296 435570 260392
rect 376448 259752 377076 259848
rect 376448 258760 376544 259752
rect 435474 259304 435570 260296
rect 435312 259208 435570 259304
rect 376448 258664 377076 258760
rect 376448 257672 376544 258664
rect 435474 258216 435570 259208
rect 435312 258120 435570 258216
rect 376448 257576 377076 257672
rect 376448 256584 376544 257576
rect 435474 257128 435570 258120
rect 435312 257032 435570 257128
rect 376448 256488 377076 256584
rect 376448 255496 376544 256488
rect 435474 256040 435570 257032
rect 435312 255944 435570 256040
rect 376448 255400 377076 255496
rect 376448 254408 376544 255400
rect 435474 254952 435570 255944
rect 435312 254856 435570 254952
rect 376448 254312 377076 254408
rect 376448 253320 376544 254312
rect 435474 253864 435570 254856
rect 435312 253768 435570 253864
rect 375632 253224 377076 253320
rect 370340 252580 371880 252676
rect 311936 252367 311942 252463
rect 312038 252367 312044 252463
rect 311942 248224 312038 252367
rect 311942 248128 312200 248224
rect 311942 247136 312038 248128
rect 371784 247680 371880 252580
rect 375632 248324 375728 253224
rect 435474 252776 435570 253768
rect 437262 277156 437358 277431
rect 437262 277060 437520 277156
rect 437262 276068 437358 277060
rect 496288 276612 496384 277604
rect 495756 276516 496384 276612
rect 437262 275972 437520 276068
rect 437262 274980 437358 275972
rect 496288 275524 496384 276516
rect 495756 275428 496384 275524
rect 437262 274884 437520 274980
rect 437262 273892 437358 274884
rect 496288 274436 496384 275428
rect 495756 274340 496384 274436
rect 437262 273796 437520 273892
rect 437262 272804 437358 273796
rect 496288 273348 496384 274340
rect 495756 273252 496384 273348
rect 437262 272708 437520 272804
rect 437262 271716 437358 272708
rect 496288 272260 496384 273252
rect 495756 272164 496384 272260
rect 437262 271620 437520 271716
rect 437262 270628 437358 271620
rect 496288 271172 496384 272164
rect 495756 271076 496384 271172
rect 437262 270532 437520 270628
rect 437262 269540 437358 270532
rect 496288 270084 496384 271076
rect 495756 269988 496384 270084
rect 437262 269444 437520 269540
rect 437262 268452 437358 269444
rect 496288 268996 496384 269988
rect 495756 268900 496384 268996
rect 437262 268356 437520 268452
rect 437262 267364 437358 268356
rect 496288 267908 496384 268900
rect 495756 267812 496384 267908
rect 437262 267268 437520 267364
rect 437262 266276 437358 267268
rect 496288 266820 496384 267812
rect 495756 266724 496384 266820
rect 437262 266180 437520 266276
rect 437262 265188 437358 266180
rect 496288 265732 496384 266724
rect 495756 265636 496384 265732
rect 437262 265092 437520 265188
rect 437262 264100 437358 265092
rect 496288 264644 496384 265636
rect 495756 264548 496384 264644
rect 437262 264004 437520 264100
rect 437262 263012 437358 264004
rect 496288 263556 496384 264548
rect 495756 263460 496384 263556
rect 437262 262916 437520 263012
rect 437262 261924 437358 262916
rect 496288 262468 496384 263460
rect 495756 262372 496384 262468
rect 437262 261828 437520 261924
rect 437262 260836 437358 261828
rect 496288 261380 496384 262372
rect 495756 261284 496384 261380
rect 437262 260740 437520 260836
rect 437262 259748 437358 260740
rect 496288 260292 496384 261284
rect 495756 260196 496384 260292
rect 437262 259652 437520 259748
rect 437262 258660 437358 259652
rect 496288 259204 496384 260196
rect 495756 259108 496384 259204
rect 437262 258564 437520 258660
rect 437262 257572 437358 258564
rect 496288 258116 496384 259108
rect 495756 258020 496384 258116
rect 437262 257476 437520 257572
rect 437262 256484 437358 257476
rect 496288 257028 496384 258020
rect 495756 256932 496384 257028
rect 437262 256388 437520 256484
rect 437262 255396 437358 256388
rect 496288 255940 496384 256932
rect 495756 255844 496384 255940
rect 437262 255300 437520 255396
rect 437262 254308 437358 255300
rect 496288 254852 496384 255844
rect 495756 254756 496384 254852
rect 437262 254212 437616 254308
rect 437262 253220 437358 254212
rect 496288 253764 496384 254756
rect 495756 253668 496384 253764
rect 437262 253217 437616 253220
rect 437256 253121 437262 253217
rect 437358 253124 437616 253217
rect 437358 253121 437364 253124
rect 435312 252680 435570 252776
rect 435474 248537 435570 252680
rect 496288 252676 496384 253668
rect 501768 278344 501864 279313
rect 560794 279313 566821 279361
rect 560794 278888 560890 279313
rect 560632 278792 560890 278888
rect 501768 278248 502396 278344
rect 501768 277256 501864 278248
rect 560794 277800 560890 278792
rect 560632 277704 560890 277800
rect 501768 277160 502396 277256
rect 501768 276168 501864 277160
rect 560794 276712 560890 277704
rect 560632 276616 560890 276712
rect 501768 276072 502396 276168
rect 501768 275080 501864 276072
rect 560794 275624 560890 276616
rect 560632 275528 560890 275624
rect 501768 274984 502396 275080
rect 501768 273992 501864 274984
rect 560794 274536 560890 275528
rect 560632 274440 560890 274536
rect 501768 273896 502396 273992
rect 501768 272904 501864 273896
rect 560794 273448 560890 274440
rect 560632 273352 560890 273448
rect 501768 272808 502396 272904
rect 501768 271816 501864 272808
rect 560794 272360 560890 273352
rect 560632 272264 560890 272360
rect 501768 271720 502396 271816
rect 501768 270728 501864 271720
rect 560794 271272 560890 272264
rect 560632 271176 560890 271272
rect 501768 270632 502396 270728
rect 501768 269640 501864 270632
rect 560794 270184 560890 271176
rect 560632 270088 560890 270184
rect 501768 269544 502396 269640
rect 501768 268552 501864 269544
rect 560794 269096 560890 270088
rect 560632 269000 560890 269096
rect 501768 268456 502396 268552
rect 501768 267464 501864 268456
rect 560794 268008 560890 269000
rect 560632 267912 560890 268008
rect 501768 267368 502396 267464
rect 501768 266376 501864 267368
rect 560794 266920 560890 267912
rect 560632 266824 560890 266920
rect 501768 266280 502396 266376
rect 501768 265288 501864 266280
rect 560794 265832 560890 266824
rect 560632 265736 560890 265832
rect 501768 265192 502396 265288
rect 501768 264200 501864 265192
rect 560794 264744 560890 265736
rect 560632 264648 560890 264744
rect 501768 264104 502396 264200
rect 501768 263112 501864 264104
rect 560794 263656 560890 264648
rect 560632 263560 560890 263656
rect 501768 263016 502396 263112
rect 501768 262024 501864 263016
rect 560794 262568 560890 263560
rect 560632 262472 560890 262568
rect 501768 261928 502396 262024
rect 501768 260936 501864 261928
rect 560794 261480 560890 262472
rect 560632 261384 560890 261480
rect 501768 260840 502396 260936
rect 501768 259848 501864 260840
rect 560794 260392 560890 261384
rect 560632 260296 560890 260392
rect 501768 259752 502396 259848
rect 501768 258760 501864 259752
rect 560794 259304 560890 260296
rect 560632 259208 560890 259304
rect 501768 258664 502396 258760
rect 501768 257672 501864 258664
rect 560794 258216 560890 259208
rect 560632 258120 560890 258216
rect 501768 257576 502396 257672
rect 501768 256584 501864 257576
rect 560794 257128 560890 258120
rect 560632 257032 560890 257128
rect 501768 256488 502396 256584
rect 501768 255496 501864 256488
rect 560794 256040 560890 257032
rect 560632 255944 560890 256040
rect 501768 255400 502396 255496
rect 501768 254408 501864 255400
rect 560794 254952 560890 255944
rect 560632 254856 560890 254952
rect 501768 254312 502396 254408
rect 501768 253320 501864 254312
rect 560794 253864 560890 254856
rect 560632 253768 560890 253864
rect 500952 253224 502396 253320
rect 495660 252580 497200 252676
rect 437256 252367 437262 252463
rect 437358 252367 437364 252463
rect 435468 248441 435474 248537
rect 435570 248441 435576 248537
rect 375632 248228 377172 248324
rect 370436 247584 371880 247680
rect 311942 247040 312200 247136
rect 311942 246048 312038 247040
rect 370968 246592 371064 247584
rect 370436 246496 371064 246592
rect 311942 245952 312200 246048
rect 311942 244960 312038 245952
rect 370968 245504 371064 246496
rect 370436 245408 371064 245504
rect 311942 244864 312200 244960
rect 311942 243872 312038 244864
rect 370968 244416 371064 245408
rect 370436 244320 371064 244416
rect 311942 243776 312200 243872
rect 311942 242784 312038 243776
rect 370968 243328 371064 244320
rect 370436 243232 371064 243328
rect 311942 242688 312200 242784
rect 311942 241696 312038 242688
rect 370968 242240 371064 243232
rect 370436 242144 371064 242240
rect 311942 241600 312200 241696
rect 311942 240608 312038 241600
rect 370968 241152 371064 242144
rect 370436 241056 371064 241152
rect 311942 240512 312200 240608
rect 311942 239520 312038 240512
rect 370968 240064 371064 241056
rect 370436 239968 371064 240064
rect 311942 239424 312200 239520
rect 311942 238432 312038 239424
rect 370968 238976 371064 239968
rect 370436 238880 371064 238976
rect 311942 238336 312200 238432
rect 311942 237344 312038 238336
rect 370968 237888 371064 238880
rect 370436 237792 371064 237888
rect 311942 237248 312200 237344
rect 311942 236256 312038 237248
rect 370968 236800 371064 237792
rect 370436 236704 371064 236800
rect 311942 236160 312200 236256
rect 311942 235168 312038 236160
rect 370968 235712 371064 236704
rect 370436 235616 371064 235712
rect 311942 235072 312200 235168
rect 311942 234080 312038 235072
rect 370968 234624 371064 235616
rect 370436 234528 371064 234624
rect 311942 233984 312200 234080
rect 311942 232992 312038 233984
rect 370968 233536 371064 234528
rect 370436 233440 371064 233536
rect 311942 232896 312200 232992
rect 311942 231904 312038 232896
rect 370968 232448 371064 233440
rect 370436 232352 371064 232448
rect 311942 231808 312200 231904
rect 311942 230816 312038 231808
rect 370968 231360 371064 232352
rect 370436 231264 371064 231360
rect 311942 230720 312200 230816
rect 311942 229728 312038 230720
rect 370968 230272 371064 231264
rect 370436 230176 371064 230272
rect 311942 229632 312200 229728
rect 311942 228640 312038 229632
rect 370968 229184 371064 230176
rect 370436 229088 371064 229184
rect 311942 228544 312200 228640
rect 311942 227552 312038 228544
rect 370968 228096 371064 229088
rect 370436 228000 371064 228096
rect 311942 227456 312200 227552
rect 311942 226464 312038 227456
rect 370968 227008 371064 228000
rect 370436 226912 371064 227008
rect 311942 226368 312200 226464
rect 311942 225376 312038 226368
rect 370968 225920 371064 226912
rect 370436 225824 371064 225920
rect 311942 225280 312200 225376
rect 311942 224288 312038 225280
rect 370968 224832 371064 225824
rect 370436 224736 371064 224832
rect 311942 224192 312200 224288
rect 311942 223200 312038 224192
rect 370968 223744 371064 224736
rect 370436 223648 371064 223744
rect 311942 223104 312200 223200
rect 311942 222112 312038 223104
rect 370968 222656 371064 223648
rect 370436 222560 371064 222656
rect 311942 222016 312200 222112
rect 311942 221024 312038 222016
rect 370968 221568 371064 222560
rect 370436 221472 371064 221568
rect 311942 220928 312200 221024
rect 311942 219936 312038 220928
rect 370968 220480 371064 221472
rect 370436 220384 371064 220480
rect 311942 219840 312200 219936
rect 311942 218848 312038 219840
rect 370968 219392 371064 220384
rect 370436 219296 371064 219392
rect 311942 218752 312200 218848
rect 311942 217760 312038 218752
rect 370968 218304 371064 219296
rect 370436 218208 371064 218304
rect 311942 217677 312200 217760
rect 306149 217664 312200 217677
rect 370968 217677 371064 218208
rect 376448 247236 376544 248228
rect 437262 248224 437358 252367
rect 437262 248128 437520 248224
rect 435468 247780 435474 247783
rect 435216 247687 435474 247780
rect 435570 247687 435576 247783
rect 435216 247684 435570 247687
rect 376448 247140 377076 247236
rect 376448 246148 376544 247140
rect 435474 246692 435570 247684
rect 435216 246596 435570 246692
rect 376448 246052 377076 246148
rect 376448 245060 376544 246052
rect 435474 245604 435570 246596
rect 435312 245508 435570 245604
rect 376448 244964 377076 245060
rect 376448 243972 376544 244964
rect 435474 244516 435570 245508
rect 435312 244420 435570 244516
rect 376448 243876 377076 243972
rect 376448 242884 376544 243876
rect 435474 243428 435570 244420
rect 435312 243332 435570 243428
rect 376448 242788 377076 242884
rect 376448 241796 376544 242788
rect 435474 242340 435570 243332
rect 435312 242244 435570 242340
rect 376448 241700 377076 241796
rect 376448 240708 376544 241700
rect 435474 241252 435570 242244
rect 435312 241156 435570 241252
rect 376448 240612 377076 240708
rect 376448 239620 376544 240612
rect 435474 240164 435570 241156
rect 435312 240068 435570 240164
rect 376448 239524 377076 239620
rect 376448 238532 376544 239524
rect 435474 239076 435570 240068
rect 435312 238980 435570 239076
rect 376448 238436 377076 238532
rect 376448 237444 376544 238436
rect 435474 237988 435570 238980
rect 435312 237892 435570 237988
rect 376448 237348 377076 237444
rect 376448 236356 376544 237348
rect 435474 236900 435570 237892
rect 435312 236804 435570 236900
rect 376448 236260 377076 236356
rect 376448 235268 376544 236260
rect 435474 235812 435570 236804
rect 435312 235716 435570 235812
rect 376448 235172 377076 235268
rect 376448 234180 376544 235172
rect 435474 234724 435570 235716
rect 435312 234628 435570 234724
rect 376448 234084 377076 234180
rect 376448 233092 376544 234084
rect 435474 233636 435570 234628
rect 435312 233540 435570 233636
rect 376448 232996 377076 233092
rect 376448 232004 376544 232996
rect 435474 232548 435570 233540
rect 435312 232452 435570 232548
rect 376448 231908 377076 232004
rect 376448 230916 376544 231908
rect 435474 231460 435570 232452
rect 435312 231364 435570 231460
rect 376448 230820 377076 230916
rect 376448 229828 376544 230820
rect 435474 230372 435570 231364
rect 435312 230276 435570 230372
rect 376448 229732 377076 229828
rect 376448 228740 376544 229732
rect 435474 229284 435570 230276
rect 435312 229188 435570 229284
rect 376448 228644 377076 228740
rect 376448 227652 376544 228644
rect 435474 228196 435570 229188
rect 435312 228100 435570 228196
rect 376448 227556 377076 227652
rect 376448 226564 376544 227556
rect 435474 227108 435570 228100
rect 435312 227012 435570 227108
rect 376448 226468 377076 226564
rect 376448 225476 376544 226468
rect 435474 226020 435570 227012
rect 435312 225924 435570 226020
rect 376448 225380 377076 225476
rect 376448 224388 376544 225380
rect 435474 224932 435570 225924
rect 435312 224836 435570 224932
rect 376448 224292 377076 224388
rect 376448 223300 376544 224292
rect 435474 223844 435570 224836
rect 435312 223748 435570 223844
rect 376448 223204 377076 223300
rect 376448 222212 376544 223204
rect 435474 222756 435570 223748
rect 435312 222660 435570 222756
rect 376448 222116 377076 222212
rect 376448 221124 376544 222116
rect 435474 221668 435570 222660
rect 435312 221572 435570 221668
rect 376448 221028 377076 221124
rect 376448 220036 376544 221028
rect 435474 220580 435570 221572
rect 435312 220484 435570 220580
rect 376448 219940 377076 220036
rect 376448 218948 376544 219940
rect 435474 219492 435570 220484
rect 435312 219396 435570 219492
rect 376448 218852 377076 218948
rect 376448 217860 376544 218852
rect 435474 218404 435570 219396
rect 435312 218308 435570 218404
rect 376448 217764 377076 217860
rect 376448 217677 376544 217764
rect 306149 217629 312038 217664
rect 306149 216701 307383 217629
rect 308407 216701 312038 217629
rect 370968 217629 376544 217677
rect 370968 217216 373176 217629
rect 370436 217120 373176 217216
rect 306149 216672 312038 216701
rect 370968 216701 373176 217120
rect 374200 216772 376544 217629
rect 435474 217316 435570 218308
rect 435312 217220 435570 217316
rect 374200 216701 377076 216772
rect 370968 216676 377076 216701
rect 306149 216653 312200 216672
rect 311942 216576 312200 216653
rect 370968 216653 376544 216676
rect 311942 215584 312038 216576
rect 370968 216128 371064 216653
rect 370436 216032 371064 216128
rect 311942 215488 312200 215584
rect 311942 214496 312038 215488
rect 370968 215040 371064 216032
rect 370436 214944 371064 215040
rect 311942 214400 312200 214496
rect 311942 213408 312038 214400
rect 370968 213952 371064 214944
rect 370436 213856 371064 213952
rect 311942 213312 312200 213408
rect 311942 212320 312038 213312
rect 370968 212864 371064 213856
rect 370436 212768 371064 212864
rect 311942 212224 312200 212320
rect 311942 211232 312038 212224
rect 370968 211776 371064 212768
rect 370436 211680 371064 211776
rect 311942 211136 312200 211232
rect 311942 210144 312038 211136
rect 370968 210688 371064 211680
rect 370436 210592 371064 210688
rect 311942 210048 312200 210144
rect 311942 209056 312038 210048
rect 370968 209600 371064 210592
rect 370436 209504 371064 209600
rect 311942 208960 312200 209056
rect 311942 207968 312038 208960
rect 370968 208512 371064 209504
rect 370436 208416 371064 208512
rect 311942 207872 312200 207968
rect 311942 206880 312038 207872
rect 370968 207424 371064 208416
rect 370436 207328 371064 207424
rect 311942 206784 312200 206880
rect 311942 205792 312038 206784
rect 370968 206336 371064 207328
rect 370436 206240 371064 206336
rect 311942 205696 312200 205792
rect 311942 204704 312038 205696
rect 370968 205248 371064 206240
rect 370436 205152 371064 205248
rect 311942 204608 312200 204704
rect 311942 203616 312038 204608
rect 370968 204160 371064 205152
rect 370436 204064 371064 204160
rect 311942 203520 312200 203616
rect 311942 202528 312038 203520
rect 370968 203072 371064 204064
rect 370436 202976 371064 203072
rect 311942 202432 312200 202528
rect 311942 201440 312038 202432
rect 370968 201984 371064 202976
rect 370436 201888 371064 201984
rect 311942 201344 312200 201440
rect 311942 200352 312038 201344
rect 370968 200896 371064 201888
rect 370436 200800 371064 200896
rect 311942 200256 312200 200352
rect 311942 199264 312038 200256
rect 370968 199808 371064 200800
rect 370436 199712 371064 199808
rect 311942 199168 312200 199264
rect 311942 198176 312038 199168
rect 370968 198720 371064 199712
rect 370436 198624 371064 198720
rect 311942 198080 312200 198176
rect 311942 197088 312038 198080
rect 370968 197632 371064 198624
rect 370436 197536 371064 197632
rect 311942 196992 312200 197088
rect 311942 196000 312038 196992
rect 370968 196544 371064 197536
rect 370436 196448 371064 196544
rect 311942 195904 312200 196000
rect 311942 194912 312038 195904
rect 370968 195456 371064 196448
rect 370436 195360 371064 195456
rect 311942 194816 312200 194912
rect 311942 193824 312038 194816
rect 370968 194368 371064 195360
rect 370436 194272 371064 194368
rect 311942 193728 312200 193824
rect 311942 192736 312038 193728
rect 370968 193280 371064 194272
rect 370436 193184 371064 193280
rect 311942 192640 312200 192736
rect 311942 191648 312038 192640
rect 370968 192192 371064 193184
rect 370436 192096 371064 192192
rect 311942 191552 312296 191648
rect 311942 190763 312038 191552
rect 370968 191104 371064 192096
rect 370436 191008 371064 191104
rect 309868 185579 309915 190663
rect 311944 190639 312038 190763
rect 311932 190543 311938 190639
rect 312046 190560 312052 190639
rect 312046 190543 312296 190560
rect 311944 190464 312296 190543
rect 311944 190124 312038 190152
rect 370968 190016 371064 191008
rect 376448 215684 376544 216653
rect 435474 216228 435570 217220
rect 435312 216132 435570 216228
rect 376448 215588 377076 215684
rect 376448 214596 376544 215588
rect 435474 215568 435570 216132
rect 437262 247136 437358 248128
rect 497104 247680 497200 252580
rect 500952 248324 501048 253224
rect 560794 252776 560890 253768
rect 560632 252680 560890 252776
rect 560794 248537 560890 252680
rect 560788 248441 560794 248537
rect 560890 248441 560896 248537
rect 500952 248228 502492 248324
rect 566745 248228 566821 253320
rect 495756 247584 497200 247680
rect 437262 247040 437520 247136
rect 437262 246048 437358 247040
rect 496288 246592 496384 247584
rect 495756 246496 496384 246592
rect 437262 245952 437520 246048
rect 437262 244960 437358 245952
rect 496288 245504 496384 246496
rect 495756 245408 496384 245504
rect 437262 244864 437520 244960
rect 437262 243872 437358 244864
rect 496288 244416 496384 245408
rect 495756 244320 496384 244416
rect 437262 243776 437520 243872
rect 437262 242784 437358 243776
rect 496288 243328 496384 244320
rect 495756 243232 496384 243328
rect 437262 242688 437520 242784
rect 437262 241696 437358 242688
rect 496288 242240 496384 243232
rect 495756 242144 496384 242240
rect 437262 241600 437520 241696
rect 437262 240608 437358 241600
rect 496288 241152 496384 242144
rect 495756 241056 496384 241152
rect 437262 240512 437520 240608
rect 437262 239520 437358 240512
rect 496288 240064 496384 241056
rect 495756 239968 496384 240064
rect 437262 239424 437520 239520
rect 437262 238432 437358 239424
rect 496288 238976 496384 239968
rect 495756 238880 496384 238976
rect 437262 238336 437520 238432
rect 437262 237344 437358 238336
rect 496288 237888 496384 238880
rect 495756 237792 496384 237888
rect 437262 237248 437520 237344
rect 437262 236256 437358 237248
rect 496288 236800 496384 237792
rect 495756 236704 496384 236800
rect 437262 236160 437520 236256
rect 437262 235168 437358 236160
rect 496288 235712 496384 236704
rect 495756 235616 496384 235712
rect 437262 235072 437520 235168
rect 437262 234080 437358 235072
rect 496288 234624 496384 235616
rect 495756 234528 496384 234624
rect 437262 233984 437520 234080
rect 437262 232992 437358 233984
rect 496288 233536 496384 234528
rect 495756 233440 496384 233536
rect 437262 232896 437520 232992
rect 437262 231904 437358 232896
rect 496288 232448 496384 233440
rect 495756 232352 496384 232448
rect 437262 231808 437520 231904
rect 437262 230816 437358 231808
rect 496288 231360 496384 232352
rect 495756 231264 496384 231360
rect 437262 230720 437520 230816
rect 437262 229728 437358 230720
rect 496288 230272 496384 231264
rect 495756 230176 496384 230272
rect 437262 229632 437520 229728
rect 437262 228640 437358 229632
rect 496288 229184 496384 230176
rect 495756 229088 496384 229184
rect 437262 228544 437520 228640
rect 437262 227552 437358 228544
rect 496288 228096 496384 229088
rect 495756 228000 496384 228096
rect 437262 227456 437520 227552
rect 437262 226464 437358 227456
rect 496288 227008 496384 228000
rect 495756 226912 496384 227008
rect 437262 226368 437520 226464
rect 437262 225376 437358 226368
rect 496288 225920 496384 226912
rect 495756 225824 496384 225920
rect 437262 225280 437520 225376
rect 437262 224288 437358 225280
rect 496288 224832 496384 225824
rect 495756 224736 496384 224832
rect 437262 224192 437520 224288
rect 437262 223200 437358 224192
rect 496288 223744 496384 224736
rect 495756 223648 496384 223744
rect 437262 223104 437520 223200
rect 437262 222112 437358 223104
rect 496288 222656 496384 223648
rect 495756 222560 496384 222656
rect 437262 222016 437520 222112
rect 437262 221024 437358 222016
rect 496288 221568 496384 222560
rect 495756 221472 496384 221568
rect 437262 220928 437520 221024
rect 437262 219936 437358 220928
rect 496288 220480 496384 221472
rect 495756 220384 496384 220480
rect 437262 219840 437520 219936
rect 437262 218848 437358 219840
rect 496288 219392 496384 220384
rect 495756 219296 496384 219392
rect 437262 218752 437520 218848
rect 437262 217760 437358 218752
rect 496288 218304 496384 219296
rect 495756 218208 496384 218304
rect 437262 217664 437520 217760
rect 496288 217677 496384 218208
rect 501768 247236 501864 248228
rect 560788 247780 560794 247783
rect 560536 247687 560794 247780
rect 560890 247687 560896 247783
rect 560536 247684 560890 247687
rect 501768 247140 502396 247236
rect 501768 246148 501864 247140
rect 560794 246692 560890 247684
rect 560536 246596 560890 246692
rect 501768 246052 502396 246148
rect 501768 245060 501864 246052
rect 560794 245604 560890 246596
rect 560632 245508 560890 245604
rect 501768 244964 502396 245060
rect 501768 243972 501864 244964
rect 560794 244516 560890 245508
rect 560632 244420 560890 244516
rect 501768 243876 502396 243972
rect 501768 242884 501864 243876
rect 560794 243428 560890 244420
rect 560632 243332 560890 243428
rect 501768 242788 502396 242884
rect 501768 241796 501864 242788
rect 560794 242340 560890 243332
rect 560632 242244 560890 242340
rect 501768 241700 502396 241796
rect 501768 240708 501864 241700
rect 560794 241252 560890 242244
rect 560632 241156 560890 241252
rect 501768 240612 502396 240708
rect 501768 239620 501864 240612
rect 560794 240164 560890 241156
rect 560632 240068 560890 240164
rect 501768 239524 502396 239620
rect 501768 238532 501864 239524
rect 560794 239076 560890 240068
rect 560632 238980 560890 239076
rect 501768 238436 502396 238532
rect 501768 237444 501864 238436
rect 560794 237988 560890 238980
rect 560632 237892 560890 237988
rect 501768 237348 502396 237444
rect 501768 236356 501864 237348
rect 560794 236900 560890 237892
rect 560632 236804 560890 236900
rect 501768 236260 502396 236356
rect 501768 235268 501864 236260
rect 560794 235812 560890 236804
rect 560632 235716 560890 235812
rect 501768 235172 502396 235268
rect 501768 234180 501864 235172
rect 560794 234724 560890 235716
rect 560632 234628 560890 234724
rect 501768 234084 502396 234180
rect 501768 233092 501864 234084
rect 560794 233636 560890 234628
rect 560632 233540 560890 233636
rect 501768 232996 502396 233092
rect 501768 232004 501864 232996
rect 560794 232548 560890 233540
rect 560632 232452 560890 232548
rect 501768 231908 502396 232004
rect 501768 230916 501864 231908
rect 560794 231460 560890 232452
rect 560632 231364 560890 231460
rect 501768 230820 502396 230916
rect 501768 229828 501864 230820
rect 560794 230372 560890 231364
rect 560632 230276 560890 230372
rect 501768 229732 502396 229828
rect 501768 228740 501864 229732
rect 560794 229284 560890 230276
rect 560632 229188 560890 229284
rect 501768 228644 502396 228740
rect 501768 227652 501864 228644
rect 560794 228196 560890 229188
rect 560632 228100 560890 228196
rect 501768 227556 502396 227652
rect 501768 226564 501864 227556
rect 560794 227108 560890 228100
rect 560632 227012 560890 227108
rect 501768 226468 502396 226564
rect 501768 225476 501864 226468
rect 560794 226020 560890 227012
rect 560632 225924 560890 226020
rect 501768 225380 502396 225476
rect 501768 224388 501864 225380
rect 560794 224932 560890 225924
rect 560632 224836 560890 224932
rect 501768 224292 502396 224388
rect 501768 223300 501864 224292
rect 560794 223844 560890 224836
rect 560632 223748 560890 223844
rect 501768 223204 502396 223300
rect 501768 222212 501864 223204
rect 560794 222756 560890 223748
rect 560632 222660 560890 222756
rect 501768 222116 502396 222212
rect 501768 221124 501864 222116
rect 560794 221668 560890 222660
rect 560632 221572 560890 221668
rect 501768 221028 502396 221124
rect 501768 220036 501864 221028
rect 560794 220580 560890 221572
rect 560632 220484 560890 220580
rect 501768 219940 502396 220036
rect 501768 218948 501864 219940
rect 560794 219492 560890 220484
rect 560632 219396 560890 219492
rect 501768 218852 502396 218948
rect 501768 217860 501864 218852
rect 560794 218404 560890 219396
rect 560632 218308 560890 218404
rect 501768 217764 502396 217860
rect 501768 217677 501864 217764
rect 437262 216672 437358 217664
rect 496288 217629 501864 217677
rect 496288 217216 498496 217629
rect 495756 217120 498496 217216
rect 496288 216701 498496 217120
rect 499520 216772 501864 217629
rect 560794 217677 560890 218308
rect 560794 217629 566821 217677
rect 560794 217316 564289 217629
rect 560632 217220 564289 217316
rect 499520 216701 502396 216772
rect 496288 216676 502396 216701
rect 560794 216701 564289 217220
rect 565313 216701 566821 217629
rect 437262 216576 437520 216672
rect 496288 216653 501864 216676
rect 437262 215584 437358 216576
rect 496288 216128 496384 216653
rect 495756 216032 496384 216128
rect 436432 215568 437075 215569
rect 435474 215563 437075 215568
rect 437262 215563 437520 215584
rect 435474 215515 437520 215563
rect 435474 215140 436583 215515
rect 435312 215044 436583 215140
rect 435474 214843 436583 215044
rect 437273 215488 437520 215515
rect 437273 214843 437358 215488
rect 496288 215040 496384 216032
rect 495756 214944 496384 215040
rect 435474 214771 437358 214843
rect 435474 214760 437075 214771
rect 376448 214500 377076 214596
rect 376448 213508 376544 214500
rect 435474 214052 435570 214760
rect 436432 214758 437075 214760
rect 435312 213956 435570 214052
rect 376448 213412 377076 213508
rect 376448 212420 376544 213412
rect 435474 212964 435570 213956
rect 435312 212868 435570 212964
rect 376448 212324 377076 212420
rect 376448 211332 376544 212324
rect 435474 211876 435570 212868
rect 435312 211780 435570 211876
rect 376448 211236 377076 211332
rect 376448 210244 376544 211236
rect 435474 210788 435570 211780
rect 435312 210692 435570 210788
rect 376448 210148 377076 210244
rect 376448 209156 376544 210148
rect 435474 209700 435570 210692
rect 435312 209604 435570 209700
rect 376448 209060 377076 209156
rect 376448 208068 376544 209060
rect 435474 208612 435570 209604
rect 435312 208516 435570 208612
rect 376448 207972 377076 208068
rect 376448 206980 376544 207972
rect 435474 207524 435570 208516
rect 435312 207428 435570 207524
rect 376448 206884 377076 206980
rect 376448 205892 376544 206884
rect 435474 206436 435570 207428
rect 435312 206340 435570 206436
rect 376448 205796 377076 205892
rect 376448 204804 376544 205796
rect 435474 205348 435570 206340
rect 435312 205252 435570 205348
rect 376448 204708 377076 204804
rect 376448 203716 376544 204708
rect 435474 204260 435570 205252
rect 435312 204164 435570 204260
rect 376448 203620 377076 203716
rect 376448 202628 376544 203620
rect 435474 203172 435570 204164
rect 435312 203076 435570 203172
rect 376448 202532 377076 202628
rect 376448 201540 376544 202532
rect 435474 202084 435570 203076
rect 435312 201988 435570 202084
rect 376448 201444 377076 201540
rect 376448 200452 376544 201444
rect 435474 200996 435570 201988
rect 435312 200900 435570 200996
rect 376448 200356 377076 200452
rect 376448 199364 376544 200356
rect 435474 199908 435570 200900
rect 435312 199812 435570 199908
rect 376448 199268 377076 199364
rect 376448 198276 376544 199268
rect 435474 198820 435570 199812
rect 435312 198724 435570 198820
rect 376448 198180 377076 198276
rect 376448 197188 376544 198180
rect 435474 197732 435570 198724
rect 435312 197636 435570 197732
rect 376448 197092 377076 197188
rect 376448 196100 376544 197092
rect 435474 196644 435570 197636
rect 435312 196548 435570 196644
rect 376448 196004 377076 196100
rect 376448 195012 376544 196004
rect 435474 195556 435570 196548
rect 435312 195460 435570 195556
rect 376448 194916 377076 195012
rect 376448 193924 376544 194916
rect 435474 194468 435570 195460
rect 435312 194372 435570 194468
rect 376448 193828 377076 193924
rect 376448 192836 376544 193828
rect 435474 193380 435570 194372
rect 435312 193284 435570 193380
rect 376448 192740 377076 192836
rect 376448 191748 376544 192740
rect 435474 192292 435570 193284
rect 435312 192196 435570 192292
rect 376448 191652 377076 191748
rect 376448 190663 376544 191652
rect 435474 191204 435570 192196
rect 435312 191108 435570 191204
rect 375661 190660 376544 190663
rect 435474 190974 435570 191108
rect 437262 214496 437358 214771
rect 437262 214400 437520 214496
rect 437262 213408 437358 214400
rect 496288 213952 496384 214944
rect 495756 213856 496384 213952
rect 437262 213312 437520 213408
rect 437262 212320 437358 213312
rect 496288 212864 496384 213856
rect 495756 212768 496384 212864
rect 437262 212224 437520 212320
rect 437262 211232 437358 212224
rect 496288 211776 496384 212768
rect 495756 211680 496384 211776
rect 437262 211136 437520 211232
rect 437262 210144 437358 211136
rect 496288 210688 496384 211680
rect 495756 210592 496384 210688
rect 437262 210048 437520 210144
rect 437262 209056 437358 210048
rect 496288 209600 496384 210592
rect 495756 209504 496384 209600
rect 437262 208960 437520 209056
rect 437262 207968 437358 208960
rect 496288 208512 496384 209504
rect 495756 208416 496384 208512
rect 437262 207872 437520 207968
rect 437262 206880 437358 207872
rect 496288 207424 496384 208416
rect 495756 207328 496384 207424
rect 437262 206784 437520 206880
rect 437262 205792 437358 206784
rect 496288 206336 496384 207328
rect 495756 206240 496384 206336
rect 437262 205696 437520 205792
rect 437262 204704 437358 205696
rect 496288 205248 496384 206240
rect 495756 205152 496384 205248
rect 437262 204608 437520 204704
rect 437262 203616 437358 204608
rect 496288 204160 496384 205152
rect 495756 204064 496384 204160
rect 437262 203520 437520 203616
rect 437262 202528 437358 203520
rect 496288 203072 496384 204064
rect 495756 202976 496384 203072
rect 437262 202432 437520 202528
rect 437262 201440 437358 202432
rect 496288 201984 496384 202976
rect 495756 201888 496384 201984
rect 437262 201344 437520 201440
rect 437262 200352 437358 201344
rect 496288 200896 496384 201888
rect 495756 200800 496384 200896
rect 437262 200256 437520 200352
rect 437262 199264 437358 200256
rect 496288 199808 496384 200800
rect 495756 199712 496384 199808
rect 437262 199168 437520 199264
rect 437262 198176 437358 199168
rect 496288 198720 496384 199712
rect 495756 198624 496384 198720
rect 437262 198080 437520 198176
rect 437262 197088 437358 198080
rect 496288 197632 496384 198624
rect 495756 197536 496384 197632
rect 437262 196992 437520 197088
rect 437262 196000 437358 196992
rect 496288 196544 496384 197536
rect 495756 196448 496384 196544
rect 437262 195904 437520 196000
rect 437262 194912 437358 195904
rect 496288 195456 496384 196448
rect 495756 195360 496384 195456
rect 437262 194816 437520 194912
rect 437262 193824 437358 194816
rect 496288 194368 496384 195360
rect 495756 194272 496384 194368
rect 437262 193728 437520 193824
rect 437262 192736 437358 193728
rect 496288 193280 496384 194272
rect 495756 193184 496384 193280
rect 437262 192640 437520 192736
rect 437262 191648 437358 192640
rect 496288 192192 496384 193184
rect 495756 192096 496384 192192
rect 437262 191552 437616 191648
rect 375661 190567 377076 190660
rect 370340 190005 371850 190016
rect 370340 189920 371851 190005
rect 309869 185568 309915 185579
rect 311944 189715 312040 189727
rect 311944 185564 312040 189619
rect 311944 185468 312200 185564
rect 311944 184610 312038 185468
rect 370436 185017 371064 185020
rect 371755 185017 371851 189920
rect 375661 185664 375757 190567
rect 376448 190564 377076 190567
rect 435474 190116 435568 190974
rect 437262 190763 437358 191552
rect 496288 191104 496384 192096
rect 495756 191008 496384 191104
rect 437264 190639 437358 190763
rect 437252 190543 437258 190639
rect 437366 190560 437372 190639
rect 437366 190543 437616 190560
rect 437264 190464 437616 190543
rect 437264 190124 437358 190152
rect 435312 190020 435568 190116
rect 435472 185965 435568 190020
rect 496288 190016 496384 191008
rect 501768 215684 501864 216653
rect 560794 216653 566821 216701
rect 560794 216228 560890 216653
rect 560632 216132 560890 216228
rect 501768 215588 502396 215684
rect 501768 214596 501864 215588
rect 560794 215140 560890 216132
rect 560632 215044 560890 215140
rect 501768 214500 502396 214596
rect 501768 213508 501864 214500
rect 560794 214052 560890 215044
rect 560632 213956 560890 214052
rect 501768 213412 502396 213508
rect 501768 212420 501864 213412
rect 560794 212964 560890 213956
rect 560632 212868 560890 212964
rect 501768 212324 502396 212420
rect 501768 211332 501864 212324
rect 560794 211876 560890 212868
rect 560632 211780 560890 211876
rect 501768 211236 502396 211332
rect 501768 210244 501864 211236
rect 560794 210788 560890 211780
rect 560632 210692 560890 210788
rect 501768 210148 502396 210244
rect 501768 209156 501864 210148
rect 560794 209700 560890 210692
rect 560632 209604 560890 209700
rect 501768 209060 502396 209156
rect 501768 208068 501864 209060
rect 560794 208612 560890 209604
rect 560632 208516 560890 208612
rect 501768 207972 502396 208068
rect 501768 206980 501864 207972
rect 560794 207524 560890 208516
rect 560632 207428 560890 207524
rect 501768 206884 502396 206980
rect 501768 205892 501864 206884
rect 560794 206436 560890 207428
rect 560632 206340 560890 206436
rect 501768 205796 502396 205892
rect 501768 204804 501864 205796
rect 560794 205348 560890 206340
rect 560632 205252 560890 205348
rect 501768 204708 502396 204804
rect 501768 203716 501864 204708
rect 560794 204260 560890 205252
rect 560632 204164 560890 204260
rect 501768 203620 502396 203716
rect 501768 202628 501864 203620
rect 560794 203172 560890 204164
rect 560632 203076 560890 203172
rect 501768 202532 502396 202628
rect 501768 201540 501864 202532
rect 560794 202084 560890 203076
rect 560632 201988 560890 202084
rect 501768 201444 502396 201540
rect 501768 200452 501864 201444
rect 560794 200996 560890 201988
rect 560632 200900 560890 200996
rect 501768 200356 502396 200452
rect 501768 199364 501864 200356
rect 560794 199908 560890 200900
rect 560632 199812 560890 199908
rect 501768 199268 502396 199364
rect 501768 198276 501864 199268
rect 560794 198820 560890 199812
rect 560632 198724 560890 198820
rect 501768 198180 502396 198276
rect 501768 197188 501864 198180
rect 560794 197732 560890 198724
rect 560632 197636 560890 197732
rect 501768 197092 502396 197188
rect 501768 196100 501864 197092
rect 560794 196644 560890 197636
rect 560632 196548 560890 196644
rect 501768 196004 502396 196100
rect 501768 195012 501864 196004
rect 560794 195556 560890 196548
rect 560632 195460 560890 195556
rect 501768 194916 502396 195012
rect 501768 193924 501864 194916
rect 560794 194468 560890 195460
rect 560632 194372 560890 194468
rect 501768 193828 502396 193924
rect 501768 192836 501864 193828
rect 560794 193380 560890 194372
rect 560632 193284 560890 193380
rect 501768 192740 502396 192836
rect 501768 191748 501864 192740
rect 560794 192292 560890 193284
rect 560632 192196 560890 192292
rect 501768 191652 502396 191748
rect 501768 190663 501864 191652
rect 560794 191204 560890 192196
rect 560632 191108 560890 191204
rect 500981 190660 501864 190663
rect 560794 190974 560890 191108
rect 500981 190567 502396 190660
rect 495660 190005 497170 190016
rect 495660 189920 497171 190005
rect 435472 185857 435568 185869
rect 437264 189715 437360 189727
rect 375661 185579 377172 185664
rect 375662 185568 377172 185579
rect 370436 184924 371851 185017
rect 311942 184476 312038 184610
rect 370968 184921 371851 184924
rect 311942 184380 312200 184476
rect 311942 183388 312038 184380
rect 370968 183932 371064 184921
rect 370436 183836 371064 183932
rect 311942 183292 312200 183388
rect 311942 182300 312038 183292
rect 370968 182844 371064 183836
rect 370436 182748 371064 182844
rect 311942 182204 312200 182300
rect 311942 181212 312038 182204
rect 370968 181756 371064 182748
rect 370436 181660 371064 181756
rect 311942 181116 312200 181212
rect 311942 180124 312038 181116
rect 370968 180668 371064 181660
rect 370436 180572 371064 180668
rect 311942 180028 312200 180124
rect 311942 179036 312038 180028
rect 370968 179580 371064 180572
rect 370436 179484 371064 179580
rect 311942 178940 312200 179036
rect 311942 177948 312038 178940
rect 370968 178492 371064 179484
rect 370436 178396 371064 178492
rect 311942 177852 312200 177948
rect 311942 176860 312038 177852
rect 370968 177404 371064 178396
rect 370436 177308 371064 177404
rect 311942 176764 312200 176860
rect 311942 175772 312038 176764
rect 370968 176316 371064 177308
rect 370436 176220 371064 176316
rect 311942 175676 312200 175772
rect 311942 174684 312038 175676
rect 370968 175228 371064 176220
rect 370436 175132 371064 175228
rect 311942 174588 312200 174684
rect 311942 173596 312038 174588
rect 370968 174140 371064 175132
rect 370436 174044 371064 174140
rect 311942 173500 312200 173596
rect 311942 172508 312038 173500
rect 370968 173052 371064 174044
rect 370436 172956 371064 173052
rect 311942 172412 312200 172508
rect 311942 171420 312038 172412
rect 370968 171964 371064 172956
rect 370436 171868 371064 171964
rect 311942 171324 312200 171420
rect 311942 170332 312038 171324
rect 370968 170876 371064 171868
rect 370436 170780 371064 170876
rect 311942 170236 312200 170332
rect 311942 169244 312038 170236
rect 370968 169788 371064 170780
rect 370436 169692 371064 169788
rect 311942 169148 312200 169244
rect 311942 168156 312038 169148
rect 370968 168700 371064 169692
rect 370436 168604 371064 168700
rect 311942 168060 312200 168156
rect 311942 167068 312038 168060
rect 370968 167612 371064 168604
rect 370436 167516 371064 167612
rect 311942 166972 312200 167068
rect 311942 165980 312038 166972
rect 370968 166524 371064 167516
rect 370436 166428 371064 166524
rect 311942 165884 312200 165980
rect 311942 164892 312038 165884
rect 370968 165436 371064 166428
rect 370436 165340 371064 165436
rect 311942 164796 312200 164892
rect 311942 163804 312038 164796
rect 370968 164348 371064 165340
rect 370436 164252 371064 164348
rect 311942 163708 312200 163804
rect 311942 162716 312038 163708
rect 370968 163260 371064 164252
rect 370436 163164 371064 163260
rect 311942 162620 312200 162716
rect 311942 161628 312038 162620
rect 370968 162172 371064 163164
rect 370436 162076 371064 162172
rect 311942 161532 312200 161628
rect 311942 160540 312038 161532
rect 370968 161084 371064 162076
rect 370436 160988 371064 161084
rect 311942 160444 312200 160540
rect 311942 159452 312038 160444
rect 370968 159996 371064 160988
rect 370436 159900 371064 159996
rect 311942 159356 312200 159452
rect 311942 158364 312038 159356
rect 370968 158908 371064 159900
rect 370436 158812 371064 158908
rect 311942 158268 312200 158364
rect 311942 157276 312038 158268
rect 370968 157820 371064 158812
rect 370436 157724 371064 157820
rect 311942 157180 312200 157276
rect 311942 156188 312038 157180
rect 370968 156732 371064 157724
rect 370436 156636 371064 156732
rect 311942 156092 312200 156188
rect 311942 155100 312038 156092
rect 370968 155644 371064 156636
rect 370436 155548 371064 155644
rect 311942 155017 312200 155100
rect 306149 155004 312200 155017
rect 370968 155017 371064 155548
rect 376448 184576 376544 185568
rect 437264 185564 437360 189619
rect 437264 185468 437520 185564
rect 435474 185432 435568 185460
rect 435216 185041 435568 185120
rect 435216 185024 435466 185041
rect 435460 184945 435466 185024
rect 435574 184945 435580 185041
rect 435474 184821 435568 184945
rect 376448 184480 377076 184576
rect 376448 183488 376544 184480
rect 435474 184032 435570 184821
rect 437264 184610 437358 185468
rect 495756 185017 496384 185020
rect 497075 185017 497171 189920
rect 500981 185664 501077 190567
rect 501768 190564 502396 190567
rect 560794 190116 560888 190974
rect 560632 190020 560888 190116
rect 560792 185965 560888 190020
rect 560792 185857 560888 185869
rect 500981 185579 502492 185664
rect 566774 185579 566821 190663
rect 500982 185568 502492 185579
rect 566775 185568 566821 185579
rect 495756 184924 497171 185017
rect 435216 183936 435570 184032
rect 376448 183392 377076 183488
rect 376448 182400 376544 183392
rect 435474 182944 435570 183936
rect 435312 182848 435570 182944
rect 376448 182304 377076 182400
rect 376448 181312 376544 182304
rect 435474 181856 435570 182848
rect 435312 181760 435570 181856
rect 376448 181216 377076 181312
rect 376448 180224 376544 181216
rect 435474 180768 435570 181760
rect 435312 180672 435570 180768
rect 376448 180128 377076 180224
rect 376448 179136 376544 180128
rect 435474 179680 435570 180672
rect 435312 179584 435570 179680
rect 376448 179040 377076 179136
rect 376448 178048 376544 179040
rect 435474 178592 435570 179584
rect 435312 178496 435570 178592
rect 376448 177952 377076 178048
rect 376448 176960 376544 177952
rect 435474 177504 435570 178496
rect 435312 177408 435570 177504
rect 376448 176864 377076 176960
rect 376448 175872 376544 176864
rect 435474 176416 435570 177408
rect 435312 176320 435570 176416
rect 376448 175776 377076 175872
rect 376448 174784 376544 175776
rect 435474 175328 435570 176320
rect 435312 175232 435570 175328
rect 376448 174688 377076 174784
rect 376448 173696 376544 174688
rect 435474 174240 435570 175232
rect 435312 174144 435570 174240
rect 376448 173600 377076 173696
rect 376448 172608 376544 173600
rect 435474 173152 435570 174144
rect 435312 173056 435570 173152
rect 376448 172512 377076 172608
rect 376448 171520 376544 172512
rect 435474 172064 435570 173056
rect 435312 171968 435570 172064
rect 376448 171424 377076 171520
rect 376448 170432 376544 171424
rect 435474 170976 435570 171968
rect 435312 170880 435570 170976
rect 376448 170336 377076 170432
rect 376448 169344 376544 170336
rect 435474 169888 435570 170880
rect 435312 169792 435570 169888
rect 376448 169248 377076 169344
rect 376448 168256 376544 169248
rect 435474 168800 435570 169792
rect 435312 168704 435570 168800
rect 376448 168160 377076 168256
rect 376448 167168 376544 168160
rect 435474 167712 435570 168704
rect 435312 167616 435570 167712
rect 376448 167072 377076 167168
rect 376448 166080 376544 167072
rect 435474 166624 435570 167616
rect 435312 166528 435570 166624
rect 376448 165984 377076 166080
rect 376448 164992 376544 165984
rect 435474 165536 435570 166528
rect 435312 165440 435570 165536
rect 376448 164896 377076 164992
rect 376448 163904 376544 164896
rect 435474 164448 435570 165440
rect 435312 164352 435570 164448
rect 376448 163808 377076 163904
rect 376448 162816 376544 163808
rect 435474 163360 435570 164352
rect 435312 163264 435570 163360
rect 376448 162720 377076 162816
rect 376448 161728 376544 162720
rect 435474 162272 435570 163264
rect 435312 162176 435570 162272
rect 376448 161632 377076 161728
rect 376448 160640 376544 161632
rect 435474 161184 435570 162176
rect 435312 161088 435570 161184
rect 376448 160544 377076 160640
rect 376448 159552 376544 160544
rect 435474 160096 435570 161088
rect 435312 160000 435570 160096
rect 376448 159456 377076 159552
rect 376448 158464 376544 159456
rect 435474 159008 435570 160000
rect 435312 158912 435570 159008
rect 376448 158368 377076 158464
rect 376448 157376 376544 158368
rect 435474 157920 435570 158912
rect 435312 157824 435570 157920
rect 376448 157280 377076 157376
rect 376448 156288 376544 157280
rect 435474 156832 435570 157824
rect 435312 156736 435570 156832
rect 376448 156192 377076 156288
rect 376448 155200 376544 156192
rect 435474 155744 435570 156736
rect 435312 155648 435570 155744
rect 376448 155104 377076 155200
rect 376448 155017 376544 155104
rect 306149 154969 312038 155004
rect 306149 154041 307383 154969
rect 308407 154041 312038 154969
rect 370968 154969 376544 155017
rect 370968 154556 373176 154969
rect 370436 154460 373176 154556
rect 306149 154012 312038 154041
rect 370968 154041 373176 154460
rect 374200 154112 376544 154969
rect 435474 154656 435570 155648
rect 435312 154560 435570 154656
rect 374200 154041 377076 154112
rect 370968 154016 377076 154041
rect 306149 153993 312200 154012
rect 311942 153916 312200 153993
rect 370968 153993 376544 154016
rect 311942 152924 312038 153916
rect 370968 153468 371064 153993
rect 370436 153372 371064 153468
rect 311942 152828 312200 152924
rect 311942 151836 312038 152828
rect 370968 152380 371064 153372
rect 370436 152284 371064 152380
rect 311942 151740 312200 151836
rect 311942 150748 312038 151740
rect 370968 151292 371064 152284
rect 370436 151196 371064 151292
rect 311942 150652 312200 150748
rect 311942 149660 312038 150652
rect 370968 150204 371064 151196
rect 370436 150108 371064 150204
rect 311942 149564 312200 149660
rect 311942 148572 312038 149564
rect 370968 149116 371064 150108
rect 370436 149020 371064 149116
rect 311942 148476 312200 148572
rect 311942 147484 312038 148476
rect 370968 148028 371064 149020
rect 370436 147932 371064 148028
rect 311942 147388 312200 147484
rect 311942 146396 312038 147388
rect 370968 146940 371064 147932
rect 370436 146844 371064 146940
rect 311942 146300 312200 146396
rect 311942 145308 312038 146300
rect 370968 145852 371064 146844
rect 370436 145756 371064 145852
rect 311942 145212 312200 145308
rect 311942 144220 312038 145212
rect 370968 144764 371064 145756
rect 370436 144668 371064 144764
rect 311942 144124 312200 144220
rect 311942 143132 312038 144124
rect 370968 143676 371064 144668
rect 370436 143580 371064 143676
rect 311942 143036 312200 143132
rect 311942 142044 312038 143036
rect 370968 142588 371064 143580
rect 370436 142492 371064 142588
rect 311942 141948 312200 142044
rect 311942 140956 312038 141948
rect 370968 141500 371064 142492
rect 370436 141404 371064 141500
rect 311942 140860 312200 140956
rect 311942 139868 312038 140860
rect 370968 140412 371064 141404
rect 370436 140316 371064 140412
rect 311942 139772 312200 139868
rect 311942 138780 312038 139772
rect 370968 139324 371064 140316
rect 370436 139228 371064 139324
rect 311942 138684 312200 138780
rect 311942 137692 312038 138684
rect 370968 138236 371064 139228
rect 370436 138140 371064 138236
rect 311942 137596 312200 137692
rect 311942 136604 312038 137596
rect 370968 137148 371064 138140
rect 370436 137052 371064 137148
rect 311942 136508 312200 136604
rect 311942 135516 312038 136508
rect 370968 136060 371064 137052
rect 370436 135964 371064 136060
rect 311942 135420 312200 135516
rect 311942 134428 312038 135420
rect 370968 134972 371064 135964
rect 370436 134876 371064 134972
rect 311942 134332 312200 134428
rect 311942 133340 312038 134332
rect 370968 133884 371064 134876
rect 370436 133788 371064 133884
rect 311942 133244 312200 133340
rect 311942 132252 312038 133244
rect 370968 132796 371064 133788
rect 370436 132700 371064 132796
rect 311942 132156 312200 132252
rect 311942 131164 312038 132156
rect 370968 131708 371064 132700
rect 370436 131612 371064 131708
rect 311942 131068 312200 131164
rect 311942 130076 312038 131068
rect 370968 130620 371064 131612
rect 370436 130524 371064 130620
rect 311942 129980 312200 130076
rect 311942 128988 312038 129980
rect 370968 129532 371064 130524
rect 370436 129436 371064 129532
rect 311942 128892 312296 128988
rect 309839 122908 309915 128000
rect 311942 127900 312038 128892
rect 370968 128444 371064 129436
rect 370436 128348 371064 128444
rect 311942 127897 312296 127900
rect 311936 127801 311942 127897
rect 312038 127804 312296 127897
rect 312038 127801 312044 127804
rect 370968 127356 371064 128348
rect 376448 153024 376544 153993
rect 435474 153568 435570 154560
rect 435312 153472 435570 153568
rect 376448 152928 377076 153024
rect 376448 151936 376544 152928
rect 435474 152908 435570 153472
rect 437262 184476 437358 184610
rect 496288 184921 497171 184924
rect 437262 184380 437520 184476
rect 437262 183388 437358 184380
rect 496288 183932 496384 184921
rect 495756 183836 496384 183932
rect 437262 183292 437520 183388
rect 437262 182300 437358 183292
rect 496288 182844 496384 183836
rect 495756 182748 496384 182844
rect 437262 182204 437520 182300
rect 437262 181212 437358 182204
rect 496288 181756 496384 182748
rect 495756 181660 496384 181756
rect 437262 181116 437520 181212
rect 437262 180124 437358 181116
rect 496288 180668 496384 181660
rect 495756 180572 496384 180668
rect 437262 180028 437520 180124
rect 437262 179036 437358 180028
rect 496288 179580 496384 180572
rect 495756 179484 496384 179580
rect 437262 178940 437520 179036
rect 437262 177948 437358 178940
rect 496288 178492 496384 179484
rect 495756 178396 496384 178492
rect 437262 177852 437520 177948
rect 437262 176860 437358 177852
rect 496288 177404 496384 178396
rect 495756 177308 496384 177404
rect 437262 176764 437520 176860
rect 437262 175772 437358 176764
rect 496288 176316 496384 177308
rect 495756 176220 496384 176316
rect 437262 175676 437520 175772
rect 437262 174684 437358 175676
rect 496288 175228 496384 176220
rect 495756 175132 496384 175228
rect 437262 174588 437520 174684
rect 437262 173596 437358 174588
rect 496288 174140 496384 175132
rect 495756 174044 496384 174140
rect 437262 173500 437520 173596
rect 437262 172508 437358 173500
rect 496288 173052 496384 174044
rect 495756 172956 496384 173052
rect 437262 172412 437520 172508
rect 437262 171420 437358 172412
rect 496288 171964 496384 172956
rect 495756 171868 496384 171964
rect 437262 171324 437520 171420
rect 437262 170332 437358 171324
rect 496288 170876 496384 171868
rect 495756 170780 496384 170876
rect 437262 170236 437520 170332
rect 437262 169244 437358 170236
rect 496288 169788 496384 170780
rect 495756 169692 496384 169788
rect 437262 169148 437520 169244
rect 437262 168156 437358 169148
rect 496288 168700 496384 169692
rect 495756 168604 496384 168700
rect 437262 168060 437520 168156
rect 437262 167068 437358 168060
rect 496288 167612 496384 168604
rect 495756 167516 496384 167612
rect 437262 166972 437520 167068
rect 437262 165980 437358 166972
rect 496288 166524 496384 167516
rect 495756 166428 496384 166524
rect 437262 165884 437520 165980
rect 437262 164892 437358 165884
rect 496288 165436 496384 166428
rect 495756 165340 496384 165436
rect 437262 164796 437520 164892
rect 437262 163804 437358 164796
rect 496288 164348 496384 165340
rect 495756 164252 496384 164348
rect 437262 163708 437520 163804
rect 437262 162716 437358 163708
rect 496288 163260 496384 164252
rect 495756 163164 496384 163260
rect 437262 162620 437520 162716
rect 437262 161628 437358 162620
rect 496288 162172 496384 163164
rect 495756 162076 496384 162172
rect 437262 161532 437520 161628
rect 437262 160540 437358 161532
rect 496288 161084 496384 162076
rect 495756 160988 496384 161084
rect 437262 160444 437520 160540
rect 437262 159452 437358 160444
rect 496288 159996 496384 160988
rect 495756 159900 496384 159996
rect 437262 159356 437520 159452
rect 437262 158364 437358 159356
rect 496288 158908 496384 159900
rect 495756 158812 496384 158908
rect 437262 158268 437520 158364
rect 437262 157276 437358 158268
rect 496288 157820 496384 158812
rect 495756 157724 496384 157820
rect 437262 157180 437520 157276
rect 437262 156188 437358 157180
rect 496288 156732 496384 157724
rect 495756 156636 496384 156732
rect 437262 156092 437520 156188
rect 437262 155100 437358 156092
rect 496288 155644 496384 156636
rect 495756 155548 496384 155644
rect 437262 155004 437520 155100
rect 496288 155017 496384 155548
rect 501768 184576 501864 185568
rect 560794 185432 560888 185460
rect 560536 185041 560888 185120
rect 560536 185024 560786 185041
rect 560780 184945 560786 185024
rect 560894 184945 560900 185041
rect 560794 184821 560888 184945
rect 501768 184480 502396 184576
rect 501768 183488 501864 184480
rect 560794 184032 560890 184821
rect 560536 183936 560890 184032
rect 501768 183392 502396 183488
rect 501768 182400 501864 183392
rect 560794 182944 560890 183936
rect 560632 182848 560890 182944
rect 501768 182304 502396 182400
rect 501768 181312 501864 182304
rect 560794 181856 560890 182848
rect 560632 181760 560890 181856
rect 501768 181216 502396 181312
rect 501768 180224 501864 181216
rect 560794 180768 560890 181760
rect 560632 180672 560890 180768
rect 501768 180128 502396 180224
rect 501768 179136 501864 180128
rect 560794 179680 560890 180672
rect 560632 179584 560890 179680
rect 501768 179040 502396 179136
rect 501768 178048 501864 179040
rect 560794 178592 560890 179584
rect 560632 178496 560890 178592
rect 501768 177952 502396 178048
rect 501768 176960 501864 177952
rect 560794 177504 560890 178496
rect 560632 177408 560890 177504
rect 501768 176864 502396 176960
rect 501768 175872 501864 176864
rect 560794 176416 560890 177408
rect 560632 176320 560890 176416
rect 501768 175776 502396 175872
rect 501768 174784 501864 175776
rect 560794 175328 560890 176320
rect 560632 175232 560890 175328
rect 501768 174688 502396 174784
rect 501768 173696 501864 174688
rect 560794 174240 560890 175232
rect 560632 174144 560890 174240
rect 501768 173600 502396 173696
rect 501768 172608 501864 173600
rect 560794 173152 560890 174144
rect 560632 173056 560890 173152
rect 501768 172512 502396 172608
rect 501768 171520 501864 172512
rect 560794 172064 560890 173056
rect 560632 171968 560890 172064
rect 501768 171424 502396 171520
rect 501768 170432 501864 171424
rect 560794 170976 560890 171968
rect 560632 170880 560890 170976
rect 501768 170336 502396 170432
rect 501768 169344 501864 170336
rect 560794 169888 560890 170880
rect 560632 169792 560890 169888
rect 501768 169248 502396 169344
rect 501768 168256 501864 169248
rect 560794 168800 560890 169792
rect 560632 168704 560890 168800
rect 501768 168160 502396 168256
rect 501768 167168 501864 168160
rect 560794 167712 560890 168704
rect 560632 167616 560890 167712
rect 501768 167072 502396 167168
rect 501768 166080 501864 167072
rect 560794 166624 560890 167616
rect 560632 166528 560890 166624
rect 501768 165984 502396 166080
rect 501768 164992 501864 165984
rect 560794 165536 560890 166528
rect 560632 165440 560890 165536
rect 501768 164896 502396 164992
rect 501768 163904 501864 164896
rect 560794 164448 560890 165440
rect 560632 164352 560890 164448
rect 501768 163808 502396 163904
rect 501768 162816 501864 163808
rect 560794 163360 560890 164352
rect 560632 163264 560890 163360
rect 501768 162720 502396 162816
rect 501768 161728 501864 162720
rect 560794 162272 560890 163264
rect 560632 162176 560890 162272
rect 501768 161632 502396 161728
rect 501768 160640 501864 161632
rect 560794 161184 560890 162176
rect 560632 161088 560890 161184
rect 501768 160544 502396 160640
rect 501768 159552 501864 160544
rect 560794 160096 560890 161088
rect 560632 160000 560890 160096
rect 501768 159456 502396 159552
rect 501768 158464 501864 159456
rect 560794 159008 560890 160000
rect 560632 158912 560890 159008
rect 501768 158368 502396 158464
rect 501768 157376 501864 158368
rect 560794 157920 560890 158912
rect 560632 157824 560890 157920
rect 501768 157280 502396 157376
rect 501768 156288 501864 157280
rect 560794 156832 560890 157824
rect 560632 156736 560890 156832
rect 501768 156192 502396 156288
rect 501768 155200 501864 156192
rect 560794 155744 560890 156736
rect 560632 155648 560890 155744
rect 501768 155104 502396 155200
rect 501768 155017 501864 155104
rect 437262 154012 437358 155004
rect 496288 154969 501864 155017
rect 496288 154556 498496 154969
rect 495756 154460 498496 154556
rect 496288 154041 498496 154460
rect 499520 154112 501864 154969
rect 560794 155017 560890 155648
rect 560794 154969 566821 155017
rect 560794 154656 564289 154969
rect 560632 154560 564289 154656
rect 499520 154041 502396 154112
rect 496288 154016 502396 154041
rect 560794 154041 564289 154560
rect 565313 154041 566821 154969
rect 437262 153916 437520 154012
rect 496288 153993 501864 154016
rect 437262 152924 437358 153916
rect 496288 153468 496384 153993
rect 495756 153372 496384 153468
rect 436432 152908 437075 152909
rect 435474 152903 437075 152908
rect 437262 152903 437520 152924
rect 435474 152855 437520 152903
rect 435474 152480 436583 152855
rect 435312 152384 436583 152480
rect 435474 152183 436583 152384
rect 437273 152828 437520 152855
rect 437273 152183 437358 152828
rect 496288 152380 496384 153372
rect 495756 152284 496384 152380
rect 435474 152111 437358 152183
rect 435474 152100 437075 152111
rect 376448 151840 377076 151936
rect 376448 150848 376544 151840
rect 435474 151392 435570 152100
rect 436432 152098 437075 152100
rect 435312 151296 435570 151392
rect 376448 150752 377076 150848
rect 376448 149760 376544 150752
rect 435474 150304 435570 151296
rect 435312 150208 435570 150304
rect 376448 149664 377076 149760
rect 376448 148672 376544 149664
rect 435474 149216 435570 150208
rect 435312 149120 435570 149216
rect 376448 148576 377076 148672
rect 376448 147584 376544 148576
rect 435474 148128 435570 149120
rect 435312 148032 435570 148128
rect 376448 147488 377076 147584
rect 376448 146496 376544 147488
rect 435474 147040 435570 148032
rect 435312 146944 435570 147040
rect 376448 146400 377076 146496
rect 376448 145408 376544 146400
rect 435474 145952 435570 146944
rect 435312 145856 435570 145952
rect 376448 145312 377076 145408
rect 376448 144320 376544 145312
rect 435474 144864 435570 145856
rect 435312 144768 435570 144864
rect 376448 144224 377076 144320
rect 376448 143232 376544 144224
rect 435474 143776 435570 144768
rect 435312 143680 435570 143776
rect 376448 143136 377076 143232
rect 376448 142144 376544 143136
rect 435474 142688 435570 143680
rect 435312 142592 435570 142688
rect 376448 142048 377076 142144
rect 376448 141056 376544 142048
rect 435474 141600 435570 142592
rect 435312 141504 435570 141600
rect 376448 140960 377076 141056
rect 376448 139968 376544 140960
rect 435474 140512 435570 141504
rect 435312 140416 435570 140512
rect 376448 139872 377076 139968
rect 376448 138880 376544 139872
rect 435474 139424 435570 140416
rect 435312 139328 435570 139424
rect 376448 138784 377076 138880
rect 376448 137792 376544 138784
rect 435474 138336 435570 139328
rect 435312 138240 435570 138336
rect 376448 137696 377076 137792
rect 376448 136704 376544 137696
rect 435474 137248 435570 138240
rect 435312 137152 435570 137248
rect 376448 136608 377076 136704
rect 376448 135616 376544 136608
rect 435474 136160 435570 137152
rect 435312 136064 435570 136160
rect 376448 135520 377076 135616
rect 376448 134528 376544 135520
rect 435474 135072 435570 136064
rect 435312 134976 435570 135072
rect 376448 134432 377076 134528
rect 376448 133440 376544 134432
rect 435474 133984 435570 134976
rect 435312 133888 435570 133984
rect 376448 133344 377076 133440
rect 376448 132352 376544 133344
rect 435474 132896 435570 133888
rect 435312 132800 435570 132896
rect 376448 132256 377076 132352
rect 376448 131264 376544 132256
rect 435474 131808 435570 132800
rect 435312 131712 435570 131808
rect 376448 131168 377076 131264
rect 376448 130176 376544 131168
rect 435474 130720 435570 131712
rect 435312 130624 435570 130720
rect 376448 130080 377076 130176
rect 376448 129088 376544 130080
rect 435474 129632 435570 130624
rect 435312 129536 435570 129632
rect 376448 128992 377076 129088
rect 376448 128000 376544 128992
rect 435474 128544 435570 129536
rect 435312 128448 435570 128544
rect 375632 127904 377076 128000
rect 370340 127260 371880 127356
rect 311936 127047 311942 127143
rect 312038 127047 312044 127143
rect 311942 122904 312038 127047
rect 311942 122808 312200 122904
rect 311942 121816 312038 122808
rect 371784 122360 371880 127260
rect 375632 123004 375728 127904
rect 435474 127456 435570 128448
rect 437262 151836 437358 152111
rect 437262 151740 437520 151836
rect 437262 150748 437358 151740
rect 496288 151292 496384 152284
rect 495756 151196 496384 151292
rect 437262 150652 437520 150748
rect 437262 149660 437358 150652
rect 496288 150204 496384 151196
rect 495756 150108 496384 150204
rect 437262 149564 437520 149660
rect 437262 148572 437358 149564
rect 496288 149116 496384 150108
rect 495756 149020 496384 149116
rect 437262 148476 437520 148572
rect 437262 147484 437358 148476
rect 496288 148028 496384 149020
rect 495756 147932 496384 148028
rect 437262 147388 437520 147484
rect 437262 146396 437358 147388
rect 496288 146940 496384 147932
rect 495756 146844 496384 146940
rect 437262 146300 437520 146396
rect 437262 145308 437358 146300
rect 496288 145852 496384 146844
rect 495756 145756 496384 145852
rect 437262 145212 437520 145308
rect 437262 144220 437358 145212
rect 496288 144764 496384 145756
rect 495756 144668 496384 144764
rect 437262 144124 437520 144220
rect 437262 143132 437358 144124
rect 496288 143676 496384 144668
rect 495756 143580 496384 143676
rect 437262 143036 437520 143132
rect 437262 142044 437358 143036
rect 496288 142588 496384 143580
rect 495756 142492 496384 142588
rect 437262 141948 437520 142044
rect 437262 140956 437358 141948
rect 496288 141500 496384 142492
rect 495756 141404 496384 141500
rect 437262 140860 437520 140956
rect 437262 139868 437358 140860
rect 496288 140412 496384 141404
rect 495756 140316 496384 140412
rect 437262 139772 437520 139868
rect 437262 138780 437358 139772
rect 496288 139324 496384 140316
rect 495756 139228 496384 139324
rect 437262 138684 437520 138780
rect 437262 137692 437358 138684
rect 496288 138236 496384 139228
rect 495756 138140 496384 138236
rect 437262 137596 437520 137692
rect 437262 136604 437358 137596
rect 496288 137148 496384 138140
rect 495756 137052 496384 137148
rect 437262 136508 437520 136604
rect 437262 135516 437358 136508
rect 496288 136060 496384 137052
rect 495756 135964 496384 136060
rect 437262 135420 437520 135516
rect 437262 134428 437358 135420
rect 496288 134972 496384 135964
rect 495756 134876 496384 134972
rect 437262 134332 437520 134428
rect 437262 133340 437358 134332
rect 496288 133884 496384 134876
rect 495756 133788 496384 133884
rect 437262 133244 437520 133340
rect 437262 132252 437358 133244
rect 496288 132796 496384 133788
rect 495756 132700 496384 132796
rect 437262 132156 437520 132252
rect 437262 131164 437358 132156
rect 496288 131708 496384 132700
rect 495756 131612 496384 131708
rect 437262 131068 437520 131164
rect 437262 130076 437358 131068
rect 496288 130620 496384 131612
rect 495756 130524 496384 130620
rect 437262 129980 437520 130076
rect 437262 128988 437358 129980
rect 496288 129532 496384 130524
rect 495756 129436 496384 129532
rect 437262 128892 437616 128988
rect 437262 127900 437358 128892
rect 496288 128444 496384 129436
rect 495756 128348 496384 128444
rect 437262 127897 437616 127900
rect 437256 127801 437262 127897
rect 437358 127804 437616 127897
rect 437358 127801 437364 127804
rect 435312 127360 435570 127456
rect 435474 123217 435570 127360
rect 496288 127356 496384 128348
rect 501768 153024 501864 153993
rect 560794 153993 566821 154041
rect 560794 153568 560890 153993
rect 560632 153472 560890 153568
rect 501768 152928 502396 153024
rect 501768 151936 501864 152928
rect 560794 152480 560890 153472
rect 560632 152384 560890 152480
rect 501768 151840 502396 151936
rect 501768 150848 501864 151840
rect 560794 151392 560890 152384
rect 560632 151296 560890 151392
rect 501768 150752 502396 150848
rect 501768 149760 501864 150752
rect 560794 150304 560890 151296
rect 560632 150208 560890 150304
rect 501768 149664 502396 149760
rect 501768 148672 501864 149664
rect 560794 149216 560890 150208
rect 560632 149120 560890 149216
rect 501768 148576 502396 148672
rect 501768 147584 501864 148576
rect 560794 148128 560890 149120
rect 560632 148032 560890 148128
rect 501768 147488 502396 147584
rect 501768 146496 501864 147488
rect 560794 147040 560890 148032
rect 560632 146944 560890 147040
rect 501768 146400 502396 146496
rect 501768 145408 501864 146400
rect 560794 145952 560890 146944
rect 560632 145856 560890 145952
rect 501768 145312 502396 145408
rect 501768 144320 501864 145312
rect 560794 144864 560890 145856
rect 560632 144768 560890 144864
rect 501768 144224 502396 144320
rect 501768 143232 501864 144224
rect 560794 143776 560890 144768
rect 560632 143680 560890 143776
rect 501768 143136 502396 143232
rect 501768 142144 501864 143136
rect 560794 142688 560890 143680
rect 560632 142592 560890 142688
rect 501768 142048 502396 142144
rect 501768 141056 501864 142048
rect 560794 141600 560890 142592
rect 560632 141504 560890 141600
rect 501768 140960 502396 141056
rect 501768 139968 501864 140960
rect 560794 140512 560890 141504
rect 560632 140416 560890 140512
rect 501768 139872 502396 139968
rect 501768 138880 501864 139872
rect 560794 139424 560890 140416
rect 560632 139328 560890 139424
rect 501768 138784 502396 138880
rect 501768 137792 501864 138784
rect 560794 138336 560890 139328
rect 560632 138240 560890 138336
rect 501768 137696 502396 137792
rect 501768 136704 501864 137696
rect 560794 137248 560890 138240
rect 560632 137152 560890 137248
rect 501768 136608 502396 136704
rect 501768 135616 501864 136608
rect 560794 136160 560890 137152
rect 560632 136064 560890 136160
rect 501768 135520 502396 135616
rect 501768 134528 501864 135520
rect 560794 135072 560890 136064
rect 560632 134976 560890 135072
rect 501768 134432 502396 134528
rect 501768 133440 501864 134432
rect 560794 133984 560890 134976
rect 560632 133888 560890 133984
rect 501768 133344 502396 133440
rect 501768 132352 501864 133344
rect 560794 132896 560890 133888
rect 560632 132800 560890 132896
rect 501768 132256 502396 132352
rect 501768 131264 501864 132256
rect 560794 131808 560890 132800
rect 560632 131712 560890 131808
rect 501768 131168 502396 131264
rect 501768 130176 501864 131168
rect 560794 130720 560890 131712
rect 560632 130624 560890 130720
rect 501768 130080 502396 130176
rect 501768 129088 501864 130080
rect 560794 129632 560890 130624
rect 560632 129536 560890 129632
rect 501768 128992 502396 129088
rect 501768 128000 501864 128992
rect 560794 128544 560890 129536
rect 560632 128448 560890 128544
rect 500952 127904 502396 128000
rect 495660 127260 497200 127356
rect 437256 127047 437262 127143
rect 437358 127047 437364 127143
rect 435468 123121 435474 123217
rect 435570 123121 435576 123217
rect 375632 122908 377172 123004
rect 370436 122264 371880 122360
rect 311942 121720 312200 121816
rect 311942 120728 312038 121720
rect 370968 121272 371064 122264
rect 370436 121176 371064 121272
rect 311942 120632 312200 120728
rect 311942 119640 312038 120632
rect 370968 120184 371064 121176
rect 370436 120088 371064 120184
rect 311942 119544 312200 119640
rect 311942 118552 312038 119544
rect 370968 119096 371064 120088
rect 370436 119000 371064 119096
rect 311942 118456 312200 118552
rect 311942 117464 312038 118456
rect 370968 118008 371064 119000
rect 370436 117912 371064 118008
rect 311942 117368 312200 117464
rect 311942 116376 312038 117368
rect 370968 116920 371064 117912
rect 370436 116824 371064 116920
rect 311942 116280 312200 116376
rect 311942 115288 312038 116280
rect 370968 115832 371064 116824
rect 370436 115736 371064 115832
rect 311942 115192 312200 115288
rect 311942 114200 312038 115192
rect 370968 114744 371064 115736
rect 370436 114648 371064 114744
rect 311942 114104 312200 114200
rect 311942 113112 312038 114104
rect 370968 113656 371064 114648
rect 370436 113560 371064 113656
rect 311942 113016 312200 113112
rect 311942 112024 312038 113016
rect 370968 112568 371064 113560
rect 370436 112472 371064 112568
rect 311942 111928 312200 112024
rect 311942 110936 312038 111928
rect 370968 111480 371064 112472
rect 370436 111384 371064 111480
rect 311942 110840 312200 110936
rect 311942 109848 312038 110840
rect 370968 110392 371064 111384
rect 370436 110296 371064 110392
rect 311942 109752 312200 109848
rect 311942 108760 312038 109752
rect 370968 109304 371064 110296
rect 370436 109208 371064 109304
rect 311942 108664 312200 108760
rect 311942 107672 312038 108664
rect 370968 108216 371064 109208
rect 370436 108120 371064 108216
rect 311942 107576 312200 107672
rect 311942 106584 312038 107576
rect 370968 107128 371064 108120
rect 370436 107032 371064 107128
rect 311942 106488 312200 106584
rect 311942 105496 312038 106488
rect 370968 106040 371064 107032
rect 370436 105944 371064 106040
rect 311942 105400 312200 105496
rect 311942 104408 312038 105400
rect 370968 104952 371064 105944
rect 370436 104856 371064 104952
rect 311942 104312 312200 104408
rect 311942 103320 312038 104312
rect 370968 103864 371064 104856
rect 370436 103768 371064 103864
rect 311942 103224 312200 103320
rect 311942 102232 312038 103224
rect 370968 102776 371064 103768
rect 370436 102680 371064 102776
rect 311942 102136 312200 102232
rect 311942 101144 312038 102136
rect 370968 101688 371064 102680
rect 370436 101592 371064 101688
rect 311942 101048 312200 101144
rect 311942 100056 312038 101048
rect 370968 100600 371064 101592
rect 370436 100504 371064 100600
rect 311942 99960 312200 100056
rect 311942 98968 312038 99960
rect 370968 99512 371064 100504
rect 370436 99416 371064 99512
rect 311942 98872 312200 98968
rect 311942 97880 312038 98872
rect 370968 98424 371064 99416
rect 370436 98328 371064 98424
rect 311942 97784 312200 97880
rect 311942 96792 312038 97784
rect 370968 97336 371064 98328
rect 370436 97240 371064 97336
rect 311942 96696 312200 96792
rect 311942 95704 312038 96696
rect 370968 96248 371064 97240
rect 370436 96152 371064 96248
rect 311942 95608 312200 95704
rect 311942 94616 312038 95608
rect 370968 95160 371064 96152
rect 370436 95064 371064 95160
rect 311942 94520 312200 94616
rect 311942 93528 312038 94520
rect 370968 94072 371064 95064
rect 370436 93976 371064 94072
rect 311942 93432 312200 93528
rect 311942 92440 312038 93432
rect 370968 92984 371064 93976
rect 370436 92888 371064 92984
rect 311942 92357 312200 92440
rect 306149 92344 312200 92357
rect 370968 92357 371064 92888
rect 376448 121916 376544 122908
rect 437262 122904 437358 127047
rect 437262 122808 437520 122904
rect 435468 122460 435474 122463
rect 435216 122367 435474 122460
rect 435570 122367 435576 122463
rect 435216 122364 435570 122367
rect 376448 121820 377076 121916
rect 376448 120828 376544 121820
rect 435474 121372 435570 122364
rect 435216 121276 435570 121372
rect 376448 120732 377076 120828
rect 376448 119740 376544 120732
rect 435474 120284 435570 121276
rect 435312 120188 435570 120284
rect 376448 119644 377076 119740
rect 376448 118652 376544 119644
rect 435474 119196 435570 120188
rect 435312 119100 435570 119196
rect 376448 118556 377076 118652
rect 376448 117564 376544 118556
rect 435474 118108 435570 119100
rect 435312 118012 435570 118108
rect 376448 117468 377076 117564
rect 376448 116476 376544 117468
rect 435474 117020 435570 118012
rect 435312 116924 435570 117020
rect 376448 116380 377076 116476
rect 376448 115388 376544 116380
rect 435474 115932 435570 116924
rect 435312 115836 435570 115932
rect 376448 115292 377076 115388
rect 376448 114300 376544 115292
rect 435474 114844 435570 115836
rect 435312 114748 435570 114844
rect 376448 114204 377076 114300
rect 376448 113212 376544 114204
rect 435474 113756 435570 114748
rect 435312 113660 435570 113756
rect 376448 113116 377076 113212
rect 376448 112124 376544 113116
rect 435474 112668 435570 113660
rect 435312 112572 435570 112668
rect 376448 112028 377076 112124
rect 376448 111036 376544 112028
rect 435474 111580 435570 112572
rect 435312 111484 435570 111580
rect 376448 110940 377076 111036
rect 376448 109948 376544 110940
rect 435474 110492 435570 111484
rect 435312 110396 435570 110492
rect 376448 109852 377076 109948
rect 376448 108860 376544 109852
rect 435474 109404 435570 110396
rect 435312 109308 435570 109404
rect 376448 108764 377076 108860
rect 376448 107772 376544 108764
rect 435474 108316 435570 109308
rect 435312 108220 435570 108316
rect 376448 107676 377076 107772
rect 376448 106684 376544 107676
rect 435474 107228 435570 108220
rect 435312 107132 435570 107228
rect 376448 106588 377076 106684
rect 376448 105596 376544 106588
rect 435474 106140 435570 107132
rect 435312 106044 435570 106140
rect 376448 105500 377076 105596
rect 376448 104508 376544 105500
rect 435474 105052 435570 106044
rect 435312 104956 435570 105052
rect 376448 104412 377076 104508
rect 376448 103420 376544 104412
rect 435474 103964 435570 104956
rect 435312 103868 435570 103964
rect 376448 103324 377076 103420
rect 376448 102332 376544 103324
rect 435474 102876 435570 103868
rect 435312 102780 435570 102876
rect 376448 102236 377076 102332
rect 376448 101244 376544 102236
rect 435474 101788 435570 102780
rect 435312 101692 435570 101788
rect 376448 101148 377076 101244
rect 376448 100156 376544 101148
rect 435474 100700 435570 101692
rect 435312 100604 435570 100700
rect 376448 100060 377076 100156
rect 376448 99068 376544 100060
rect 435474 99612 435570 100604
rect 435312 99516 435570 99612
rect 376448 98972 377076 99068
rect 376448 97980 376544 98972
rect 435474 98524 435570 99516
rect 435312 98428 435570 98524
rect 376448 97884 377076 97980
rect 376448 96892 376544 97884
rect 435474 97436 435570 98428
rect 435312 97340 435570 97436
rect 376448 96796 377076 96892
rect 376448 95804 376544 96796
rect 435474 96348 435570 97340
rect 435312 96252 435570 96348
rect 376448 95708 377076 95804
rect 376448 94716 376544 95708
rect 435474 95260 435570 96252
rect 435312 95164 435570 95260
rect 376448 94620 377076 94716
rect 376448 93628 376544 94620
rect 435474 94172 435570 95164
rect 435312 94076 435570 94172
rect 376448 93532 377076 93628
rect 376448 92540 376544 93532
rect 435474 93084 435570 94076
rect 435312 92988 435570 93084
rect 376448 92444 377076 92540
rect 376448 92357 376544 92444
rect 306149 92309 312038 92344
rect 306149 91381 307383 92309
rect 308407 91381 312038 92309
rect 370968 92309 376544 92357
rect 370968 91896 373176 92309
rect 370436 91800 373176 91896
rect 306149 91352 312038 91381
rect 370968 91381 373176 91800
rect 374200 91452 376544 92309
rect 435474 91996 435570 92988
rect 435312 91900 435570 91996
rect 374200 91381 377076 91452
rect 370968 91356 377076 91381
rect 306149 91333 312200 91352
rect 311942 91256 312200 91333
rect 370968 91333 376544 91356
rect 311942 90264 312038 91256
rect 370968 90808 371064 91333
rect 370436 90712 371064 90808
rect 311942 90168 312200 90264
rect 311942 89176 312038 90168
rect 370968 89720 371064 90712
rect 370436 89624 371064 89720
rect 311942 89080 312200 89176
rect 311942 88088 312038 89080
rect 370968 88632 371064 89624
rect 370436 88536 371064 88632
rect 311942 87992 312200 88088
rect 311942 87000 312038 87992
rect 370968 87544 371064 88536
rect 370436 87448 371064 87544
rect 311942 86904 312200 87000
rect 311942 85912 312038 86904
rect 370968 86456 371064 87448
rect 370436 86360 371064 86456
rect 311942 85816 312200 85912
rect 311942 84824 312038 85816
rect 370968 85368 371064 86360
rect 370436 85272 371064 85368
rect 311942 84728 312200 84824
rect 311942 83736 312038 84728
rect 370968 84280 371064 85272
rect 370436 84184 371064 84280
rect 311942 83640 312200 83736
rect 311942 82648 312038 83640
rect 370968 83192 371064 84184
rect 370436 83096 371064 83192
rect 311942 82552 312200 82648
rect 311942 81560 312038 82552
rect 370968 82104 371064 83096
rect 370436 82008 371064 82104
rect 311942 81464 312200 81560
rect 311942 80472 312038 81464
rect 370968 81016 371064 82008
rect 370436 80920 371064 81016
rect 311942 80376 312200 80472
rect 311942 79384 312038 80376
rect 370968 79928 371064 80920
rect 370436 79832 371064 79928
rect 311942 79288 312200 79384
rect 311942 78296 312038 79288
rect 370968 78840 371064 79832
rect 370436 78744 371064 78840
rect 311942 78200 312200 78296
rect 311942 77208 312038 78200
rect 370968 77752 371064 78744
rect 370436 77656 371064 77752
rect 311942 77112 312200 77208
rect 311942 76120 312038 77112
rect 370968 76664 371064 77656
rect 370436 76568 371064 76664
rect 311942 76024 312200 76120
rect 311942 75032 312038 76024
rect 370968 75576 371064 76568
rect 370436 75480 371064 75576
rect 311942 74936 312200 75032
rect 311942 73944 312038 74936
rect 370968 74488 371064 75480
rect 370436 74392 371064 74488
rect 311942 73848 312200 73944
rect 311942 72856 312038 73848
rect 370968 73400 371064 74392
rect 370436 73304 371064 73400
rect 311942 72760 312200 72856
rect 311942 71768 312038 72760
rect 370968 72312 371064 73304
rect 370436 72216 371064 72312
rect 311942 71672 312200 71768
rect 311942 70680 312038 71672
rect 370968 71224 371064 72216
rect 370436 71128 371064 71224
rect 311942 70584 312200 70680
rect 311942 69592 312038 70584
rect 370968 70136 371064 71128
rect 370436 70040 371064 70136
rect 311942 69496 312200 69592
rect 311942 68504 312038 69496
rect 370968 69048 371064 70040
rect 370436 68952 371064 69048
rect 311942 68408 312200 68504
rect 311942 67416 312038 68408
rect 370968 67960 371064 68952
rect 370436 67864 371064 67960
rect 311942 67320 312200 67416
rect 311942 66328 312038 67320
rect 370968 66872 371064 67864
rect 370436 66776 371064 66872
rect 311942 66232 312296 66328
rect 311942 65443 312038 66232
rect 370968 65784 371064 66776
rect 370436 65688 371064 65784
rect 311944 65319 312038 65443
rect 311932 65223 311938 65319
rect 312046 65240 312052 65319
rect 312046 65223 312296 65240
rect 311944 65144 312296 65223
rect 311944 64804 312038 64832
rect 370968 64696 371064 65688
rect 376448 90364 376544 91333
rect 435474 90908 435570 91900
rect 435312 90812 435570 90908
rect 376448 90268 377076 90364
rect 376448 89276 376544 90268
rect 435474 90249 435570 90812
rect 437262 121816 437358 122808
rect 497104 122360 497200 127260
rect 500952 123004 501048 127904
rect 560794 127456 560890 128448
rect 560632 127360 560890 127456
rect 560794 123217 560890 127360
rect 560788 123121 560794 123217
rect 560890 123121 560896 123217
rect 500952 122908 502492 123004
rect 495756 122264 497200 122360
rect 437262 121720 437520 121816
rect 437262 120728 437358 121720
rect 496288 121272 496384 122264
rect 495756 121176 496384 121272
rect 437262 120632 437520 120728
rect 437262 119640 437358 120632
rect 496288 120184 496384 121176
rect 495756 120088 496384 120184
rect 437262 119544 437520 119640
rect 437262 118552 437358 119544
rect 496288 119096 496384 120088
rect 495756 119000 496384 119096
rect 437262 118456 437520 118552
rect 437262 117464 437358 118456
rect 496288 118008 496384 119000
rect 495756 117912 496384 118008
rect 437262 117368 437520 117464
rect 437262 116376 437358 117368
rect 496288 116920 496384 117912
rect 495756 116824 496384 116920
rect 437262 116280 437520 116376
rect 437262 115288 437358 116280
rect 496288 115832 496384 116824
rect 495756 115736 496384 115832
rect 437262 115192 437520 115288
rect 437262 114200 437358 115192
rect 496288 114744 496384 115736
rect 495756 114648 496384 114744
rect 437262 114104 437520 114200
rect 437262 113112 437358 114104
rect 496288 113656 496384 114648
rect 495756 113560 496384 113656
rect 437262 113016 437520 113112
rect 437262 112024 437358 113016
rect 496288 112568 496384 113560
rect 495756 112472 496384 112568
rect 437262 111928 437520 112024
rect 437262 110936 437358 111928
rect 496288 111480 496384 112472
rect 495756 111384 496384 111480
rect 437262 110840 437520 110936
rect 437262 109848 437358 110840
rect 496288 110392 496384 111384
rect 495756 110296 496384 110392
rect 437262 109752 437520 109848
rect 437262 108760 437358 109752
rect 496288 109304 496384 110296
rect 495756 109208 496384 109304
rect 437262 108664 437520 108760
rect 437262 107672 437358 108664
rect 496288 108216 496384 109208
rect 495756 108120 496384 108216
rect 437262 107576 437520 107672
rect 437262 106584 437358 107576
rect 496288 107128 496384 108120
rect 495756 107032 496384 107128
rect 437262 106488 437520 106584
rect 437262 105496 437358 106488
rect 496288 106040 496384 107032
rect 495756 105944 496384 106040
rect 437262 105400 437520 105496
rect 437262 104408 437358 105400
rect 496288 104952 496384 105944
rect 495756 104856 496384 104952
rect 437262 104312 437520 104408
rect 437262 103320 437358 104312
rect 496288 103864 496384 104856
rect 495756 103768 496384 103864
rect 437262 103224 437520 103320
rect 437262 102232 437358 103224
rect 496288 102776 496384 103768
rect 495756 102680 496384 102776
rect 437262 102136 437520 102232
rect 437262 101144 437358 102136
rect 496288 101688 496384 102680
rect 495756 101592 496384 101688
rect 437262 101048 437520 101144
rect 437262 100056 437358 101048
rect 496288 100600 496384 101592
rect 495756 100504 496384 100600
rect 437262 99960 437520 100056
rect 437262 98968 437358 99960
rect 496288 99512 496384 100504
rect 495756 99416 496384 99512
rect 437262 98872 437520 98968
rect 437262 97880 437358 98872
rect 496288 98424 496384 99416
rect 495756 98328 496384 98424
rect 437262 97784 437520 97880
rect 437262 96792 437358 97784
rect 496288 97336 496384 98328
rect 495756 97240 496384 97336
rect 437262 96696 437520 96792
rect 437262 95704 437358 96696
rect 496288 96248 496384 97240
rect 495756 96152 496384 96248
rect 437262 95608 437520 95704
rect 437262 94616 437358 95608
rect 496288 95160 496384 96152
rect 495756 95064 496384 95160
rect 437262 94520 437520 94616
rect 437262 93528 437358 94520
rect 496288 94072 496384 95064
rect 495756 93976 496384 94072
rect 437262 93432 437520 93528
rect 437262 92440 437358 93432
rect 496288 92984 496384 93976
rect 495756 92888 496384 92984
rect 437262 92344 437520 92440
rect 496288 92357 496384 92888
rect 501768 121916 501864 122908
rect 560788 122460 560794 122463
rect 560536 122367 560794 122460
rect 560890 122367 560896 122463
rect 560536 122364 560890 122367
rect 501768 121820 502396 121916
rect 501768 120828 501864 121820
rect 560794 121372 560890 122364
rect 560536 121276 560890 121372
rect 501768 120732 502396 120828
rect 501768 119740 501864 120732
rect 560794 120284 560890 121276
rect 560632 120188 560890 120284
rect 501768 119644 502396 119740
rect 501768 118652 501864 119644
rect 560794 119196 560890 120188
rect 560632 119100 560890 119196
rect 501768 118556 502396 118652
rect 501768 117564 501864 118556
rect 560794 118108 560890 119100
rect 560632 118012 560890 118108
rect 501768 117468 502396 117564
rect 501768 116476 501864 117468
rect 560794 117020 560890 118012
rect 560632 116924 560890 117020
rect 501768 116380 502396 116476
rect 501768 115388 501864 116380
rect 560794 115932 560890 116924
rect 560632 115836 560890 115932
rect 501768 115292 502396 115388
rect 501768 114300 501864 115292
rect 560794 114844 560890 115836
rect 560632 114748 560890 114844
rect 501768 114204 502396 114300
rect 501768 113212 501864 114204
rect 560794 113756 560890 114748
rect 560632 113660 560890 113756
rect 501768 113116 502396 113212
rect 501768 112124 501864 113116
rect 560794 112668 560890 113660
rect 560632 112572 560890 112668
rect 501768 112028 502396 112124
rect 501768 111036 501864 112028
rect 560794 111580 560890 112572
rect 560632 111484 560890 111580
rect 501768 110940 502396 111036
rect 501768 109948 501864 110940
rect 560794 110492 560890 111484
rect 560632 110396 560890 110492
rect 501768 109852 502396 109948
rect 501768 108860 501864 109852
rect 560794 109404 560890 110396
rect 560632 109308 560890 109404
rect 501768 108764 502396 108860
rect 501768 107772 501864 108764
rect 560794 108316 560890 109308
rect 560632 108220 560890 108316
rect 501768 107676 502396 107772
rect 501768 106684 501864 107676
rect 560794 107228 560890 108220
rect 560632 107132 560890 107228
rect 501768 106588 502396 106684
rect 501768 105596 501864 106588
rect 560794 106140 560890 107132
rect 560632 106044 560890 106140
rect 501768 105500 502396 105596
rect 501768 104508 501864 105500
rect 560794 105052 560890 106044
rect 560632 104956 560890 105052
rect 501768 104412 502396 104508
rect 501768 103420 501864 104412
rect 560794 103964 560890 104956
rect 560632 103868 560890 103964
rect 501768 103324 502396 103420
rect 501768 102332 501864 103324
rect 560794 102876 560890 103868
rect 560632 102780 560890 102876
rect 501768 102236 502396 102332
rect 501768 101244 501864 102236
rect 560794 101788 560890 102780
rect 560632 101692 560890 101788
rect 501768 101148 502396 101244
rect 501768 100156 501864 101148
rect 560794 100700 560890 101692
rect 560632 100604 560890 100700
rect 501768 100060 502396 100156
rect 501768 99068 501864 100060
rect 560794 99612 560890 100604
rect 560632 99516 560890 99612
rect 501768 98972 502396 99068
rect 501768 97980 501864 98972
rect 560794 98524 560890 99516
rect 560632 98428 560890 98524
rect 501768 97884 502396 97980
rect 501768 96892 501864 97884
rect 560794 97436 560890 98428
rect 560632 97340 560890 97436
rect 501768 96796 502396 96892
rect 501768 95804 501864 96796
rect 560794 96348 560890 97340
rect 560632 96252 560890 96348
rect 501768 95708 502396 95804
rect 501768 94716 501864 95708
rect 560794 95260 560890 96252
rect 560632 95164 560890 95260
rect 501768 94620 502396 94716
rect 501768 93628 501864 94620
rect 560794 94172 560890 95164
rect 560632 94076 560890 94172
rect 501768 93532 502396 93628
rect 501768 92540 501864 93532
rect 560794 93084 560890 94076
rect 560632 92988 560890 93084
rect 501768 92444 502396 92540
rect 501768 92357 501864 92444
rect 437262 91352 437358 92344
rect 496288 92309 501864 92357
rect 496288 91896 498496 92309
rect 495756 91800 498496 91896
rect 496288 91381 498496 91800
rect 499520 91452 501864 92309
rect 560794 92357 560890 92988
rect 560794 92309 566198 92357
rect 560794 91996 564289 92309
rect 560632 91900 564289 91996
rect 499520 91381 502396 91452
rect 496288 91356 502396 91381
rect 560794 91381 564289 91900
rect 565313 91381 566198 92309
rect 437262 91256 437520 91352
rect 496288 91333 501864 91356
rect 437262 90264 437358 91256
rect 496288 90808 496384 91333
rect 495756 90712 496384 90808
rect 435474 90243 437075 90249
rect 437262 90243 437520 90264
rect 435474 90195 437520 90243
rect 435474 89820 436583 90195
rect 435312 89724 436583 89820
rect 435474 89523 436583 89724
rect 437273 90168 437520 90195
rect 437273 89523 437358 90168
rect 496288 89720 496384 90712
rect 495756 89624 496384 89720
rect 435474 89451 437358 89523
rect 435474 89438 437075 89451
rect 376448 89180 377076 89276
rect 376448 88188 376544 89180
rect 435474 88732 435570 89438
rect 435312 88636 435570 88732
rect 376448 88092 377076 88188
rect 376448 87100 376544 88092
rect 435474 87644 435570 88636
rect 435312 87548 435570 87644
rect 376448 87004 377076 87100
rect 376448 86012 376544 87004
rect 435474 86556 435570 87548
rect 435312 86460 435570 86556
rect 376448 85916 377076 86012
rect 376448 84924 376544 85916
rect 435474 85468 435570 86460
rect 435312 85372 435570 85468
rect 376448 84828 377076 84924
rect 376448 83836 376544 84828
rect 435474 84380 435570 85372
rect 435312 84284 435570 84380
rect 376448 83740 377076 83836
rect 376448 82748 376544 83740
rect 435474 83292 435570 84284
rect 435312 83196 435570 83292
rect 376448 82652 377076 82748
rect 376448 81660 376544 82652
rect 435474 82204 435570 83196
rect 435312 82108 435570 82204
rect 376448 81564 377076 81660
rect 376448 80572 376544 81564
rect 435474 81116 435570 82108
rect 435312 81020 435570 81116
rect 376448 80476 377076 80572
rect 376448 79484 376544 80476
rect 435474 80028 435570 81020
rect 435312 79932 435570 80028
rect 376448 79388 377076 79484
rect 376448 78396 376544 79388
rect 435474 78940 435570 79932
rect 435312 78844 435570 78940
rect 376448 78300 377076 78396
rect 376448 77308 376544 78300
rect 435474 77852 435570 78844
rect 435312 77756 435570 77852
rect 376448 77212 377076 77308
rect 376448 76220 376544 77212
rect 435474 76764 435570 77756
rect 435312 76668 435570 76764
rect 376448 76124 377076 76220
rect 376448 75132 376544 76124
rect 435474 75676 435570 76668
rect 435312 75580 435570 75676
rect 376448 75036 377076 75132
rect 376448 74044 376544 75036
rect 435474 74588 435570 75580
rect 435312 74492 435570 74588
rect 376448 73948 377076 74044
rect 376448 72956 376544 73948
rect 435474 73500 435570 74492
rect 435312 73404 435570 73500
rect 376448 72860 377076 72956
rect 376448 71868 376544 72860
rect 435474 72412 435570 73404
rect 435312 72316 435570 72412
rect 376448 71772 377076 71868
rect 376448 70780 376544 71772
rect 435474 71324 435570 72316
rect 435312 71228 435570 71324
rect 376448 70684 377076 70780
rect 376448 69692 376544 70684
rect 435474 70236 435570 71228
rect 435312 70140 435570 70236
rect 376448 69596 377076 69692
rect 376448 68604 376544 69596
rect 435474 69148 435570 70140
rect 435312 69052 435570 69148
rect 376448 68508 377076 68604
rect 376448 67516 376544 68508
rect 435474 68060 435570 69052
rect 435312 67964 435570 68060
rect 376448 67420 377076 67516
rect 376448 66428 376544 67420
rect 435474 66972 435570 67964
rect 435312 66876 435570 66972
rect 376448 66332 377076 66428
rect 376448 65343 376544 66332
rect 435474 65884 435570 66876
rect 435312 65788 435570 65884
rect 375661 65340 376544 65343
rect 435474 65654 435570 65788
rect 437262 89176 437358 89451
rect 437262 89080 437520 89176
rect 437262 88088 437358 89080
rect 496288 88632 496384 89624
rect 495756 88536 496384 88632
rect 437262 87992 437520 88088
rect 437262 87000 437358 87992
rect 496288 87544 496384 88536
rect 495756 87448 496384 87544
rect 437262 86904 437520 87000
rect 437262 85912 437358 86904
rect 496288 86456 496384 87448
rect 495756 86360 496384 86456
rect 437262 85816 437520 85912
rect 437262 84824 437358 85816
rect 496288 85368 496384 86360
rect 495756 85272 496384 85368
rect 437262 84728 437520 84824
rect 437262 83736 437358 84728
rect 496288 84280 496384 85272
rect 495756 84184 496384 84280
rect 437262 83640 437520 83736
rect 437262 82648 437358 83640
rect 496288 83192 496384 84184
rect 495756 83096 496384 83192
rect 437262 82552 437520 82648
rect 437262 81560 437358 82552
rect 496288 82104 496384 83096
rect 495756 82008 496384 82104
rect 437262 81464 437520 81560
rect 437262 80472 437358 81464
rect 496288 81016 496384 82008
rect 495756 80920 496384 81016
rect 437262 80376 437520 80472
rect 437262 79384 437358 80376
rect 496288 79928 496384 80920
rect 495756 79832 496384 79928
rect 437262 79288 437520 79384
rect 437262 78296 437358 79288
rect 496288 78840 496384 79832
rect 495756 78744 496384 78840
rect 437262 78200 437520 78296
rect 437262 77208 437358 78200
rect 496288 77752 496384 78744
rect 495756 77656 496384 77752
rect 437262 77112 437520 77208
rect 437262 76120 437358 77112
rect 496288 76664 496384 77656
rect 495756 76568 496384 76664
rect 437262 76024 437520 76120
rect 437262 75032 437358 76024
rect 496288 75576 496384 76568
rect 495756 75480 496384 75576
rect 437262 74936 437520 75032
rect 437262 73944 437358 74936
rect 496288 74488 496384 75480
rect 495756 74392 496384 74488
rect 437262 73848 437520 73944
rect 437262 72856 437358 73848
rect 496288 73400 496384 74392
rect 495756 73304 496384 73400
rect 437262 72760 437520 72856
rect 437262 71768 437358 72760
rect 496288 72312 496384 73304
rect 495756 72216 496384 72312
rect 437262 71672 437520 71768
rect 437262 70680 437358 71672
rect 496288 71224 496384 72216
rect 495756 71128 496384 71224
rect 437262 70584 437520 70680
rect 437262 69592 437358 70584
rect 496288 70136 496384 71128
rect 495756 70040 496384 70136
rect 437262 69496 437520 69592
rect 437262 68504 437358 69496
rect 496288 69048 496384 70040
rect 495756 68952 496384 69048
rect 437262 68408 437520 68504
rect 437262 67416 437358 68408
rect 496288 67960 496384 68952
rect 495756 67864 496384 67960
rect 437262 67320 437520 67416
rect 437262 66328 437358 67320
rect 496288 66872 496384 67864
rect 495756 66776 496384 66872
rect 437262 66232 437616 66328
rect 375661 65247 377076 65340
rect 370340 64685 371850 64696
rect 370340 64600 371851 64685
rect 311944 64395 312040 64407
rect 311944 62472 312040 64299
rect 371755 62472 371851 64600
rect 375661 62472 375757 65247
rect 376448 65244 377076 65247
rect 435474 64796 435568 65654
rect 437262 65443 437358 66232
rect 496288 65784 496384 66776
rect 495756 65688 496384 65784
rect 437264 65319 437358 65443
rect 437252 65240 437372 65319
rect 437252 65223 437616 65240
rect 437264 65144 437616 65223
rect 435312 64700 435568 64796
rect 435472 64243 435568 64700
rect 496288 64696 496384 65688
rect 501768 90364 501864 91333
rect 560794 91333 566198 91381
rect 560794 90908 560890 91333
rect 560632 90812 560890 90908
rect 501768 90268 502396 90364
rect 501768 89276 501864 90268
rect 560794 89820 560890 90812
rect 560632 89724 560890 89820
rect 501768 89180 502396 89276
rect 501768 88188 501864 89180
rect 560794 88732 560890 89724
rect 560632 88636 560890 88732
rect 501768 88092 502396 88188
rect 501768 87100 501864 88092
rect 560794 87644 560890 88636
rect 560632 87548 560890 87644
rect 501768 87004 502396 87100
rect 501768 86012 501864 87004
rect 560794 86556 560890 87548
rect 560632 86460 560890 86556
rect 501768 85916 502396 86012
rect 501768 84924 501864 85916
rect 560794 85468 560890 86460
rect 560632 85372 560890 85468
rect 501768 84828 502396 84924
rect 501768 83836 501864 84828
rect 560794 84380 560890 85372
rect 560632 84284 560890 84380
rect 501768 83740 502396 83836
rect 501768 82748 501864 83740
rect 560794 83292 560890 84284
rect 560632 83196 560890 83292
rect 501768 82652 502396 82748
rect 501768 81660 501864 82652
rect 560794 82204 560890 83196
rect 560632 82108 560890 82204
rect 501768 81564 502396 81660
rect 501768 80572 501864 81564
rect 560794 81116 560890 82108
rect 560632 81020 560890 81116
rect 501768 80476 502396 80572
rect 501768 79484 501864 80476
rect 560794 80028 560890 81020
rect 560632 79932 560890 80028
rect 501768 79388 502396 79484
rect 501768 78396 501864 79388
rect 560794 78940 560890 79932
rect 560632 78844 560890 78940
rect 501768 78300 502396 78396
rect 501768 77308 501864 78300
rect 560794 77852 560890 78844
rect 560632 77756 560890 77852
rect 501768 77212 502396 77308
rect 501768 76220 501864 77212
rect 560794 76764 560890 77756
rect 560632 76668 560890 76764
rect 501768 76124 502396 76220
rect 501768 75132 501864 76124
rect 560794 75676 560890 76668
rect 560632 75580 560890 75676
rect 501768 75036 502396 75132
rect 501768 74044 501864 75036
rect 560794 74588 560890 75580
rect 560632 74492 560890 74588
rect 501768 73948 502396 74044
rect 501768 72956 501864 73948
rect 560794 73500 560890 74492
rect 560632 73404 560890 73500
rect 501768 72860 502396 72956
rect 501768 71868 501864 72860
rect 560794 72412 560890 73404
rect 560632 72316 560890 72412
rect 501768 71772 502396 71868
rect 501768 70780 501864 71772
rect 560794 71324 560890 72316
rect 560632 71228 560890 71324
rect 501768 70684 502396 70780
rect 501768 69692 501864 70684
rect 560794 70236 560890 71228
rect 560632 70140 560890 70236
rect 501768 69596 502396 69692
rect 501768 68604 501864 69596
rect 560794 69148 560890 70140
rect 560632 69052 560890 69148
rect 501768 68508 502396 68604
rect 501768 67516 501864 68508
rect 560794 68060 560890 69052
rect 560632 67964 560890 68060
rect 501768 67420 502396 67516
rect 501768 66428 501864 67420
rect 560794 66972 560890 67964
rect 560632 66876 560890 66972
rect 501768 66332 502396 66428
rect 501768 65343 501864 66332
rect 560794 65884 560890 66876
rect 560632 65788 560890 65884
rect 500981 65340 501864 65343
rect 560794 65654 560890 65788
rect 500981 65247 502396 65340
rect 495660 64685 497170 64696
rect 495660 64600 497171 64685
rect 497075 62472 497171 64600
rect 500981 62472 501077 65247
rect 501768 65244 502396 65247
rect 560794 64796 560888 65654
rect 560632 64700 560888 64796
rect 560792 62472 560888 64700
<< via1 >>
rect 102332 651892 102424 651972
rect 95870 644429 96526 646722
rect 119296 646120 119388 646200
rect 119128 645916 119228 646006
rect 119968 645938 120060 646018
rect 127470 642700 128350 642780
rect 123830 642040 123960 642610
rect 131500 642060 131630 642630
rect 127460 641880 128340 641960
rect 119290 640060 119382 640140
rect 119128 639582 119228 639672
rect 120010 639576 120102 639656
rect 115455 637499 115663 638077
rect 126070 636580 126950 636660
rect 129100 635900 129230 636470
rect 126080 635680 126960 635760
rect 119292 633678 119384 633758
rect 119138 633304 119220 633388
rect 119936 633142 120028 633222
rect 126290 630500 127170 630580
rect 129170 629840 129300 630410
rect 126290 629690 127170 629770
rect 119308 627140 119400 627220
rect 119136 626806 119218 626890
rect 119918 626702 120010 626782
rect 126540 623980 127420 624060
rect 128820 623320 128950 623890
rect 126540 623170 127420 623250
rect 119296 620764 119388 620844
rect 119142 620400 119224 620484
rect 119950 620294 120042 620374
rect 128380 618620 128860 618680
rect 128380 618400 128860 618460
rect 131940 618240 132070 618810
rect 119304 614284 119396 614364
rect 119142 613974 119224 614058
rect 119978 613888 120070 613968
rect 128030 611170 128510 611230
rect 128030 610800 128510 610860
rect 131590 610790 131720 611360
rect 119308 607978 119400 608058
rect 119138 607592 119220 607676
rect 119914 607480 120006 607560
rect 128160 605120 128640 605180
rect 128160 604650 128640 604710
rect 131720 604640 131850 605310
rect 119296 601686 119388 601766
rect 119144 601222 119226 601306
rect 119958 601104 120050 601184
rect 127960 598860 128440 598920
rect 127960 598290 128440 598350
rect 131520 598280 131650 599050
rect 119336 594154 119428 594234
rect 119104 593672 119186 593756
rect 119926 593546 120018 593626
rect 119610 592870 119690 592880
rect 119610 592810 119620 592870
rect 119620 592810 119680 592870
rect 119680 592810 119690 592870
rect 119610 592800 119690 592810
rect 127920 591310 128400 591370
rect 127920 590640 128400 590700
rect 131480 590630 131610 591500
rect 119306 584602 119398 584682
rect 119144 584130 119226 584214
rect 120128 584028 120220 584108
rect 119650 583330 119730 583340
rect 119650 583270 119660 583330
rect 119660 583270 119720 583330
rect 119720 583270 119730 583330
rect 119650 583260 119730 583270
rect 128370 582330 128870 582390
rect 128370 582110 128870 582170
rect 132890 581950 133020 582520
rect 119318 575480 119410 575560
rect 119138 575094 119220 575178
rect 120036 575004 120128 575084
rect 119690 574310 119770 574320
rect 119690 574250 119700 574310
rect 119700 574250 119760 574310
rect 119760 574250 119770 574310
rect 119690 574240 119770 574250
rect 128410 573310 128910 573370
rect 128410 572990 128910 573050
rect 132930 572830 133060 573500
rect 119374 567962 119466 568042
rect 119134 567426 119216 567510
rect 119994 567302 120086 567382
rect 119640 566640 119720 566650
rect 119640 566580 119650 566640
rect 119650 566580 119710 566640
rect 119710 566580 119720 566640
rect 119640 566570 119720 566580
rect 128360 565640 128860 565700
rect 128360 565220 128860 565280
rect 132880 565060 133010 565830
rect 119314 561344 119406 561424
rect 119124 560864 119206 560948
rect 120034 560874 120126 560954
rect 435472 561829 435568 561925
rect 119640 560100 119720 560110
rect 119640 560040 119650 560100
rect 119650 560040 119710 560100
rect 119710 560040 119720 560100
rect 119640 560030 119720 560040
rect 128360 559100 128860 559160
rect 128360 558580 128860 558640
rect 132880 558420 133010 559290
rect 119350 554560 119442 554640
rect 119132 553978 119214 554062
rect 120078 553952 120170 554032
rect 119710 553270 119790 553280
rect 119710 553210 119720 553270
rect 119720 553210 119780 553270
rect 119780 553210 119790 553270
rect 119710 553200 119790 553210
rect 128830 552270 129380 552330
rect 128830 552050 129380 552110
rect 133900 551890 134030 552460
rect 119336 546942 119428 547022
rect 119128 546408 119210 546492
rect 120170 546368 120262 546448
rect 119710 545700 119790 545710
rect 119710 545640 119720 545700
rect 119720 545640 119780 545700
rect 119780 545640 119790 545700
rect 119710 545630 119790 545640
rect 128830 544700 129380 544760
rect 128830 544280 129380 544340
rect 133900 544120 134030 544890
rect 119318 538902 119410 538982
rect 119132 538390 119214 538474
rect 120046 538344 120138 538424
rect 119680 537640 119760 537650
rect 119680 537580 119690 537640
rect 119690 537580 119750 537640
rect 119750 537580 119760 537640
rect 119680 537570 119760 537580
rect 128800 536640 129350 536700
rect 128800 536020 129350 536080
rect 133870 535860 134000 536830
rect 435466 560905 435574 561001
rect 560792 561829 560888 561925
rect 307383 530001 308407 530929
rect 373176 530001 374200 530929
rect 311942 503761 312038 503857
rect 560786 560905 560894 561001
rect 498496 530001 499520 530929
rect 564289 530001 565313 530929
rect 436583 528143 437273 528815
rect 311942 503007 312038 503103
rect 437262 503761 437358 503857
rect 437262 503007 437358 503103
rect 435474 499081 435570 499177
rect 435474 498327 435570 498423
rect 307383 467341 308407 468269
rect 373176 467341 374200 468269
rect 311938 441183 312046 441279
rect 560794 499081 560890 499177
rect 560794 498327 560890 498423
rect 498496 467341 499520 468269
rect 564289 467341 565313 468269
rect 436583 465483 437273 466155
rect 311944 440259 312040 440355
rect 437258 441183 437366 441279
rect 435472 436509 435568 436605
rect 437264 440259 437360 440355
rect 435466 435585 435574 435681
rect 560792 436509 560888 436605
rect 307383 404681 308407 405609
rect 373176 404681 374200 405609
rect 311942 378441 312038 378537
rect 560786 435585 560894 435681
rect 498496 404681 499520 405609
rect 564289 404681 565313 405609
rect 436583 402823 437273 403495
rect 311942 377687 312038 377783
rect 437262 378441 437358 378537
rect 437262 377687 437358 377783
rect 435474 373761 435570 373857
rect 435474 373007 435570 373103
rect 307383 342021 308407 342949
rect 373176 342021 374200 342949
rect 311938 315863 312046 315959
rect 560794 373761 560890 373857
rect 560794 373007 560890 373103
rect 498496 342021 499520 342949
rect 564289 342021 565313 342949
rect 436583 340163 437273 340835
rect 311944 314939 312040 315035
rect 437258 315863 437366 315959
rect 435472 311189 435568 311285
rect 437264 314939 437360 315035
rect 435466 310265 435574 310361
rect 560792 311189 560888 311285
rect 307383 279361 308407 280289
rect 373176 279361 374200 280289
rect 311942 253121 312038 253217
rect 560786 310265 560894 310361
rect 498496 279361 499520 280289
rect 564289 279361 565313 280289
rect 436583 277503 437273 278175
rect 311942 252367 312038 252463
rect 437262 253121 437358 253217
rect 437262 252367 437358 252463
rect 435474 248441 435570 248537
rect 435474 247687 435570 247783
rect 307383 216701 308407 217629
rect 373176 216701 374200 217629
rect 311938 190543 312046 190639
rect 560794 248441 560890 248537
rect 560794 247687 560890 247783
rect 498496 216701 499520 217629
rect 564289 216701 565313 217629
rect 436583 214843 437273 215515
rect 311944 189619 312040 189715
rect 437258 190543 437366 190639
rect 435472 185869 435568 185965
rect 437264 189619 437360 189715
rect 435466 184945 435574 185041
rect 560792 185869 560888 185965
rect 307383 154041 308407 154969
rect 373176 154041 374200 154969
rect 311942 127801 312038 127897
rect 560786 184945 560894 185041
rect 498496 154041 499520 154969
rect 564289 154041 565313 154969
rect 436583 152183 437273 152855
rect 311942 127047 312038 127143
rect 437262 127801 437358 127897
rect 437262 127047 437358 127143
rect 435474 123121 435570 123217
rect 435474 122367 435570 122463
rect 307383 91381 308407 92309
rect 373176 91381 374200 92309
rect 311938 65223 312046 65319
rect 560794 123121 560890 123217
rect 560794 122367 560890 122463
rect 498496 91381 499520 92309
rect 564289 91381 565313 92309
rect 436583 89523 437273 90195
rect 311944 64299 312040 64395
<< metal2 >>
rect 110936 654114 117074 654170
rect 102943 654016 103167 654048
rect 102943 653874 102991 654016
rect 103145 653874 103167 654016
rect 102943 653840 103167 653874
rect 105519 654041 105743 654073
rect 105519 653899 105567 654041
rect 105721 653899 105743 654041
rect 105519 653865 105743 653899
rect 108275 654056 108499 654088
rect 108275 653914 108323 654056
rect 108477 653914 108499 654056
rect 110936 653914 110992 654114
rect 113619 653915 113843 653947
rect 108275 653880 108499 653914
rect 105600 653794 105656 653865
rect 108356 653809 108412 653880
rect 113619 653773 113667 653915
rect 113821 653773 113843 653915
rect 116272 653774 116874 653830
rect 113619 653739 113843 653773
rect 113700 653668 113756 653739
rect 102308 651972 102442 651990
rect 102308 651892 102332 651972
rect 102424 651892 102442 651972
rect 102308 651870 102442 651892
rect 95499 646722 96634 646815
rect 95499 644429 95870 646722
rect 96526 644429 96634 646722
rect 95499 644298 96634 644429
rect 103948 636952 104004 637032
rect 112040 636952 112096 637002
rect 101366 636922 101486 636952
rect 101366 636822 101376 636922
rect 101456 636822 101486 636922
rect 101366 636802 101486 636822
rect 103946 636922 104066 636952
rect 103946 636822 103956 636922
rect 104036 636822 104066 636922
rect 103946 636802 104066 636822
rect 96576 634523 96764 634558
rect 96576 634384 96598 634523
rect 96722 634474 96764 634523
rect 106704 634474 106760 636920
rect 109236 636902 109386 636942
rect 109236 636822 109266 636902
rect 109356 636822 109386 636902
rect 109236 636802 109386 636822
rect 111996 636912 112146 636952
rect 111996 636832 112026 636912
rect 112116 636832 112146 636912
rect 111996 636812 112146 636832
rect 114432 636150 114488 638270
rect 115410 638077 115696 638189
rect 115410 637499 115455 638077
rect 115663 637499 115696 638077
rect 115410 637416 115696 637499
rect 114620 636862 114676 636912
rect 114576 636822 114726 636862
rect 114576 636742 114606 636822
rect 114696 636742 114726 636822
rect 114576 636722 114726 636742
rect 107078 636094 114488 636150
rect 96722 634418 106760 634474
rect 96722 634384 96764 634418
rect 96576 634360 96764 634384
rect 96583 634245 96771 634280
rect 96583 634106 96605 634245
rect 96729 634185 96771 634245
rect 107079 634185 107134 636094
rect 116818 635930 116874 653774
rect 96729 634130 107134 634185
rect 96729 634106 96771 634130
rect 107079 634124 107134 634130
rect 107368 635874 116874 635930
rect 96583 634082 96771 634106
rect 96591 633985 96779 634020
rect 96591 633846 96613 633985
rect 96737 633955 96779 633985
rect 107368 633955 107424 635874
rect 117018 635600 117074 654114
rect 119272 646200 119406 646218
rect 119272 646120 119296 646200
rect 119388 646120 119406 646200
rect 119272 646098 119406 646120
rect 119112 646006 119242 646020
rect 119112 645916 119128 646006
rect 119228 645916 119242 646006
rect 119944 646018 120078 646036
rect 119944 645938 119968 646018
rect 120060 645938 120078 646018
rect 119944 645916 120078 645938
rect 119112 645902 119242 645916
rect 127460 642780 128360 642790
rect 127460 642700 127470 642780
rect 128350 642700 128360 642780
rect 127460 642690 128360 642700
rect 131470 642630 131660 642650
rect 123800 642610 123990 642630
rect 123800 642040 123830 642610
rect 123960 642040 123990 642610
rect 131470 642060 131500 642630
rect 131630 642060 131660 642630
rect 131470 642040 131660 642060
rect 123800 642020 123990 642040
rect 127450 641960 128350 641970
rect 127450 641880 127460 641960
rect 128340 641880 128350 641960
rect 127450 641870 128350 641880
rect 119266 640140 119400 640158
rect 119266 640060 119290 640140
rect 119382 640060 119400 640140
rect 119266 640038 119400 640060
rect 119112 639672 119242 639686
rect 119112 639582 119128 639672
rect 119228 639582 119242 639672
rect 119112 639568 119242 639582
rect 119986 639656 120120 639674
rect 119986 639576 120010 639656
rect 120102 639576 120120 639656
rect 119986 639554 120120 639576
rect 126060 636660 126960 636670
rect 126060 636580 126070 636660
rect 126950 636580 126960 636660
rect 126060 636570 126960 636580
rect 129070 636470 129260 636490
rect 129070 635900 129100 636470
rect 129230 635900 129260 636470
rect 129070 635880 129260 635900
rect 126070 635760 126970 635770
rect 126070 635680 126080 635760
rect 126960 635680 126970 635760
rect 126070 635670 126970 635680
rect 96737 633899 107424 633955
rect 96737 633846 96779 633899
rect 107368 633866 107424 633899
rect 107668 635544 117074 635600
rect 96591 633822 96779 633846
rect 107668 633766 107724 635544
rect 96634 633735 107724 633766
rect 96598 633710 107724 633735
rect 96598 633700 96786 633710
rect 107668 633708 107724 633710
rect 119268 633758 119402 633776
rect 96598 633561 96620 633700
rect 96744 633561 96786 633700
rect 119268 633678 119292 633758
rect 119384 633678 119402 633758
rect 119268 633656 119402 633678
rect 96598 633537 96786 633561
rect 119128 633388 119234 633400
rect 119128 633304 119138 633388
rect 119220 633304 119234 633388
rect 119128 633294 119234 633304
rect 119912 633222 120046 633240
rect 119912 633142 119936 633222
rect 120028 633142 120046 633222
rect 119912 633120 120046 633142
rect 126280 630580 127180 630590
rect 126280 630500 126290 630580
rect 127170 630500 127180 630580
rect 126280 630490 127180 630500
rect 129140 630410 129330 630430
rect 129140 629840 129170 630410
rect 129300 629840 129330 630410
rect 129140 629820 129330 629840
rect 126280 629770 127180 629780
rect 126280 629690 126290 629770
rect 127170 629690 127180 629770
rect 126280 629680 127180 629690
rect 119284 627220 119418 627238
rect 119284 627140 119308 627220
rect 119400 627140 119418 627220
rect 119284 627118 119418 627140
rect 119126 626890 119232 626902
rect 119126 626806 119136 626890
rect 119218 626806 119232 626890
rect 119126 626796 119232 626806
rect 119894 626782 120028 626800
rect 119894 626702 119918 626782
rect 120010 626702 120028 626782
rect 119894 626680 120028 626702
rect 126530 624060 127430 624070
rect 126530 623980 126540 624060
rect 127420 623980 127430 624060
rect 126530 623970 127430 623980
rect 128790 623890 128980 623910
rect 128790 623320 128820 623890
rect 128950 623320 128980 623890
rect 128790 623300 128980 623320
rect 126530 623250 127430 623260
rect 126530 623170 126540 623250
rect 127420 623170 127430 623250
rect 126530 623160 127430 623170
rect 119272 620844 119406 620862
rect 119272 620764 119296 620844
rect 119388 620764 119406 620844
rect 119272 620742 119406 620764
rect 119132 620484 119238 620496
rect 119132 620400 119142 620484
rect 119224 620400 119238 620484
rect 119132 620390 119238 620400
rect 119926 620374 120060 620392
rect 119926 620294 119950 620374
rect 120042 620294 120060 620374
rect 119926 620272 120060 620294
rect 128360 619460 128880 619480
rect 128360 619330 128380 619460
rect 128860 619330 128880 619460
rect 128360 618680 128880 619330
rect 128360 618620 128380 618680
rect 128860 618620 128880 618680
rect 128360 618610 128880 618620
rect 131910 618810 132100 618830
rect 128360 618460 128880 618470
rect 128360 618400 128380 618460
rect 128860 618400 128880 618460
rect 128360 617710 128880 618400
rect 131910 618240 131940 618810
rect 132070 618240 132100 618810
rect 131910 618220 132100 618240
rect 128360 617580 128380 617710
rect 128860 617580 128880 617710
rect 128360 617560 128880 617580
rect 119280 614364 119414 614382
rect 119280 614284 119304 614364
rect 119396 614284 119414 614364
rect 119280 614262 119414 614284
rect 119132 614058 119238 614070
rect 119132 613974 119142 614058
rect 119224 613974 119238 614058
rect 119132 613964 119238 613974
rect 119954 613968 120088 613986
rect 119954 613888 119978 613968
rect 120070 613888 120088 613968
rect 119954 613866 120088 613888
rect 128010 612010 128530 612030
rect 128010 611880 128030 612010
rect 128510 611880 128530 612010
rect 128010 611230 128530 611880
rect 128010 611170 128030 611230
rect 128510 611170 128530 611230
rect 128010 611160 128530 611170
rect 131560 611360 131750 611380
rect 128010 610860 128530 610870
rect 128010 610800 128030 610860
rect 128510 610800 128530 610860
rect 128010 610260 128530 610800
rect 131560 610790 131590 611360
rect 131720 610790 131750 611360
rect 131560 610770 131750 610790
rect 128010 610130 128030 610260
rect 128510 610130 128530 610260
rect 128010 610110 128530 610130
rect 119284 608058 119418 608076
rect 119284 607978 119308 608058
rect 119400 607978 119418 608058
rect 119284 607956 119418 607978
rect 119128 607676 119234 607688
rect 119128 607592 119138 607676
rect 119220 607592 119234 607676
rect 119128 607582 119234 607592
rect 119890 607560 120024 607578
rect 119890 607480 119914 607560
rect 120006 607480 120024 607560
rect 119890 607458 120024 607480
rect 128140 605960 128660 605980
rect 128140 605830 128160 605960
rect 128640 605830 128660 605960
rect 128140 605180 128660 605830
rect 128140 605120 128160 605180
rect 128640 605120 128660 605180
rect 128140 605110 128660 605120
rect 131690 605310 131880 605330
rect 128140 604710 128660 604720
rect 128140 604650 128160 604710
rect 128640 604650 128660 604710
rect 128140 604110 128660 604650
rect 131690 604640 131720 605310
rect 131850 604640 131880 605310
rect 131690 604620 131880 604640
rect 128140 603980 128160 604110
rect 128640 603980 128660 604110
rect 128140 603960 128660 603980
rect 119272 601766 119406 601784
rect 119272 601686 119296 601766
rect 119388 601686 119406 601766
rect 119272 601664 119406 601686
rect 119134 601306 119240 601318
rect 119134 601222 119144 601306
rect 119226 601222 119240 601306
rect 119134 601212 119240 601222
rect 119934 601184 120068 601202
rect 119934 601104 119958 601184
rect 120050 601104 120068 601184
rect 119934 601082 120068 601104
rect 127940 599700 128460 599720
rect 127940 599570 127960 599700
rect 128440 599570 128460 599700
rect 127940 598920 128460 599570
rect 127940 598860 127960 598920
rect 128440 598860 128460 598920
rect 127940 598850 128460 598860
rect 131490 599050 131680 599070
rect 127940 598350 128460 598360
rect 127940 598290 127960 598350
rect 128440 598290 128460 598350
rect 127940 597750 128460 598290
rect 131490 598280 131520 599050
rect 131650 598280 131680 599050
rect 131490 598260 131680 598280
rect 127940 597620 127960 597750
rect 128440 597620 128460 597750
rect 127940 597600 128460 597620
rect 119312 594234 119446 594252
rect 119312 594154 119336 594234
rect 119428 594154 119446 594234
rect 119312 594132 119446 594154
rect 119094 593756 119200 593768
rect 119094 593672 119104 593756
rect 119186 593672 119200 593756
rect 119094 593662 119200 593672
rect 119902 593626 120036 593644
rect 119902 593546 119926 593626
rect 120018 593546 120036 593626
rect 119902 593524 120036 593546
rect 118690 592880 119700 592890
rect 118690 592800 118700 592880
rect 118790 592800 119610 592880
rect 119690 592800 119700 592880
rect 118690 592790 119700 592800
rect 127900 592150 128420 592170
rect 127900 592020 127920 592150
rect 128400 592020 128420 592150
rect 127900 591370 128420 592020
rect 127900 591310 127920 591370
rect 128400 591310 128420 591370
rect 127900 591300 128420 591310
rect 131450 591500 131640 591520
rect 127900 590700 128420 590710
rect 127900 590640 127920 590700
rect 128400 590640 128420 590700
rect 127900 590100 128420 590640
rect 131450 590630 131480 591500
rect 131610 590630 131640 591500
rect 131450 590610 131640 590630
rect 127900 589970 127920 590100
rect 128400 589970 128420 590100
rect 127900 589950 128420 589970
rect 119282 584682 119416 584700
rect 119282 584602 119306 584682
rect 119398 584602 119416 584682
rect 119282 584580 119416 584602
rect 119134 584214 119240 584226
rect 119134 584130 119144 584214
rect 119226 584130 119240 584214
rect 119134 584120 119240 584130
rect 120104 584108 120238 584126
rect 120104 584028 120128 584108
rect 120220 584028 120238 584108
rect 120104 584006 120238 584028
rect 118730 583340 119740 583350
rect 118730 583260 118740 583340
rect 118830 583260 119650 583340
rect 119730 583260 119740 583340
rect 118730 583250 119740 583260
rect 128360 583170 128880 583200
rect 128360 583040 128380 583170
rect 128860 583040 128880 583170
rect 128360 582390 128880 583040
rect 128360 582330 128370 582390
rect 128870 582330 128880 582390
rect 132860 582520 133050 582540
rect 128360 582110 128370 582170
rect 128870 582110 128880 582170
rect 128360 581422 128880 582110
rect 132860 581950 132890 582520
rect 133020 581950 133050 582520
rect 132860 581930 133050 581950
rect 128360 581292 128376 581422
rect 128856 581292 128880 581422
rect 128360 581260 128880 581292
rect 119294 575560 119428 575578
rect 119294 575480 119318 575560
rect 119410 575480 119428 575560
rect 119294 575458 119428 575480
rect 119128 575178 119234 575190
rect 119128 575094 119138 575178
rect 119220 575094 119234 575178
rect 119128 575084 119234 575094
rect 120012 575084 120146 575102
rect 120012 575004 120036 575084
rect 120128 575004 120146 575084
rect 120012 574982 120146 575004
rect 118770 574320 119780 574330
rect 118770 574240 118780 574320
rect 118870 574240 119690 574320
rect 119770 574240 119780 574320
rect 118770 574230 119780 574240
rect 128400 574150 128920 574180
rect 128400 574020 128420 574150
rect 128900 574020 128920 574150
rect 128400 573370 128920 574020
rect 128400 573310 128410 573370
rect 128910 573310 128920 573370
rect 132900 573500 133090 573520
rect 128400 572990 128410 573050
rect 128910 572990 128920 573050
rect 128400 572302 128920 572990
rect 132900 572830 132930 573500
rect 133060 572830 133090 573500
rect 132900 572810 133090 572830
rect 128400 572172 128416 572302
rect 128896 572172 128920 572302
rect 128400 572140 128920 572172
rect 119350 568042 119484 568060
rect 119350 567962 119374 568042
rect 119466 567962 119484 568042
rect 119350 567940 119484 567962
rect 119124 567510 119230 567522
rect 119124 567426 119134 567510
rect 119216 567426 119230 567510
rect 119124 567416 119230 567426
rect 119970 567382 120104 567400
rect 119970 567302 119994 567382
rect 120086 567302 120104 567382
rect 119970 567280 120104 567302
rect 118720 566650 119730 566660
rect 118720 566570 118730 566650
rect 118820 566570 119640 566650
rect 119720 566570 119730 566650
rect 118720 566560 119730 566570
rect 128350 566480 128870 566510
rect 128350 566350 128370 566480
rect 128850 566350 128870 566480
rect 128350 565700 128870 566350
rect 128350 565640 128360 565700
rect 128860 565640 128870 565700
rect 132850 565830 133040 565850
rect 128350 565220 128360 565280
rect 128860 565220 128870 565280
rect 128350 564532 128870 565220
rect 132850 565060 132880 565830
rect 133010 565060 133040 565830
rect 132850 565040 133040 565060
rect 128350 564402 128376 564532
rect 128856 564402 128870 564532
rect 128350 564370 128870 564402
rect 337242 563696 402174 563752
rect 337242 562954 337298 563696
rect 402118 562952 402174 563696
rect 462562 563696 527494 563752
rect 462562 562954 462618 563696
rect 527438 562952 527494 563696
rect 435466 561829 435472 561925
rect 435568 561829 435574 561925
rect 119290 561424 119424 561442
rect 119290 561344 119314 561424
rect 119406 561344 119424 561424
rect 119290 561322 119424 561344
rect 435466 561001 435574 561829
rect 119114 560948 119220 560960
rect 119114 560864 119124 560948
rect 119206 560864 119220 560948
rect 119114 560854 119220 560864
rect 120010 560954 120144 560972
rect 120010 560874 120034 560954
rect 120126 560874 120144 560954
rect 435466 560899 435574 560905
rect 560786 561829 560792 561925
rect 560888 561829 560894 561925
rect 560786 561001 560894 561829
rect 560786 560899 560894 560905
rect 120010 560852 120144 560874
rect 118720 560110 119730 560120
rect 118720 560030 118730 560110
rect 118820 560030 119640 560110
rect 119720 560030 119730 560110
rect 118720 560020 119730 560030
rect 128350 559940 128870 559970
rect 128350 559810 128370 559940
rect 128850 559810 128870 559940
rect 128350 559160 128870 559810
rect 128350 559100 128360 559160
rect 128860 559100 128870 559160
rect 132850 559290 133040 559310
rect 128350 558580 128360 558640
rect 128860 558580 128870 558640
rect 128350 557892 128870 558580
rect 132850 558420 132880 559290
rect 133010 558420 133040 559290
rect 132850 558400 133040 558420
rect 128350 557762 128376 557892
rect 128856 557762 128870 557892
rect 128350 557730 128870 557762
rect 119326 554640 119460 554658
rect 119326 554560 119350 554640
rect 119442 554560 119460 554640
rect 119326 554538 119460 554560
rect 119122 554062 119228 554074
rect 119122 553978 119132 554062
rect 119214 553978 119228 554062
rect 119122 553968 119228 553978
rect 120054 554032 120188 554050
rect 120054 553952 120078 554032
rect 120170 553952 120188 554032
rect 120054 553930 120188 553952
rect 118790 553280 119800 553290
rect 118790 553200 118800 553280
rect 118890 553200 119710 553280
rect 119790 553200 119800 553280
rect 118790 553190 119800 553200
rect 128820 553110 129390 553140
rect 128820 552980 128840 553110
rect 129370 552980 129390 553110
rect 128820 552330 129390 552980
rect 128820 552270 128830 552330
rect 129380 552270 129390 552330
rect 133870 552460 134060 552480
rect 128820 552050 128830 552110
rect 129380 552050 129390 552110
rect 128820 551362 129390 552050
rect 133870 551890 133900 552460
rect 134030 551890 134060 552460
rect 133870 551870 134060 551890
rect 128820 551232 128846 551362
rect 129326 551232 129390 551362
rect 128820 551200 129390 551232
rect 119312 547022 119446 547040
rect 119312 546942 119336 547022
rect 119428 546942 119446 547022
rect 119312 546920 119446 546942
rect 119118 546492 119224 546504
rect 119118 546408 119128 546492
rect 119210 546408 119224 546492
rect 119118 546398 119224 546408
rect 120146 546448 120280 546466
rect 120146 546368 120170 546448
rect 120262 546368 120280 546448
rect 120146 546346 120280 546368
rect 118790 545710 119800 545720
rect 118790 545630 118800 545710
rect 118890 545630 119710 545710
rect 119790 545630 119800 545710
rect 118790 545620 119800 545630
rect 128820 545540 129390 545570
rect 128820 545410 128840 545540
rect 129370 545410 129390 545540
rect 128820 544760 129390 545410
rect 128820 544700 128830 544760
rect 129380 544700 129390 544760
rect 133870 544890 134060 544910
rect 128820 544280 128830 544340
rect 129380 544280 129390 544340
rect 128820 543592 129390 544280
rect 133870 544120 133900 544890
rect 134030 544120 134060 544890
rect 133870 544100 134060 544120
rect 128820 543462 128866 543592
rect 129346 543462 129390 543592
rect 128820 543430 129390 543462
rect 119294 538982 119428 539000
rect 119294 538902 119318 538982
rect 119410 538902 119428 538982
rect 119294 538880 119428 538902
rect 119122 538474 119228 538486
rect 119122 538390 119132 538474
rect 119214 538390 119228 538474
rect 119122 538380 119228 538390
rect 120022 538424 120156 538442
rect 120022 538344 120046 538424
rect 120138 538344 120156 538424
rect 120022 538322 120156 538344
rect 118760 537650 119770 537660
rect 118760 537570 118770 537650
rect 118860 537570 119680 537650
rect 119760 537570 119770 537650
rect 118760 537560 119770 537570
rect 128790 537480 129360 537510
rect 128790 537350 128810 537480
rect 129340 537350 129360 537480
rect 128790 536700 129360 537350
rect 128790 536640 128800 536700
rect 129350 536640 129360 536700
rect 133840 536830 134030 536850
rect 128790 536020 128800 536080
rect 129350 536020 129360 536080
rect 128790 535342 129360 536020
rect 133840 535860 133870 536830
rect 134000 535860 134030 536830
rect 133840 535840 134030 535860
rect 128790 535212 128826 535342
rect 129306 535212 129360 535342
rect 128790 535170 129360 535212
rect 307335 530929 308448 530969
rect 307335 530001 307383 530929
rect 308407 530001 308448 530929
rect 307335 529957 308448 530001
rect 373128 530929 374241 530969
rect 373128 530001 373176 530929
rect 374200 530001 374241 530929
rect 373128 529957 374241 530001
rect 498448 530929 499561 530969
rect 498448 530001 498496 530929
rect 499520 530001 499561 530929
rect 498448 529957 499561 530001
rect 564241 530929 565354 530969
rect 564241 530001 564289 530929
rect 565313 530001 565354 530929
rect 564241 529957 565354 530001
rect 436522 528815 437319 528863
rect 436522 528143 436583 528815
rect 437273 528143 437319 528815
rect 436522 528071 437319 528143
rect 311942 503857 312038 503863
rect 311942 503103 312038 503761
rect 311942 503001 312038 503007
rect 437262 503857 437358 503863
rect 437262 503103 437358 503761
rect 437262 503001 437358 503007
rect 345338 501092 345394 501892
rect 410214 501148 410270 501890
rect 337242 501036 345394 501092
rect 402118 501092 410270 501148
rect 470658 501092 470714 501892
rect 535534 501148 535590 501890
rect 337242 500294 337298 501036
rect 402118 500292 402174 501092
rect 462562 501036 470714 501092
rect 527438 501092 535590 501148
rect 462562 500294 462618 501036
rect 527438 500292 527494 501092
rect 435474 499177 435570 499183
rect 435474 498423 435570 499081
rect 435474 498321 435570 498327
rect 560794 499177 560890 499183
rect 560794 498423 560890 499081
rect 560794 498321 560890 498327
rect 307335 468269 308448 468309
rect 307335 467341 307383 468269
rect 308407 467341 308448 468269
rect 307335 467297 308448 467341
rect 373128 468269 374241 468309
rect 373128 467341 373176 468269
rect 374200 467341 374241 468269
rect 373128 467297 374241 467341
rect 498448 468269 499561 468309
rect 498448 467341 498496 468269
rect 499520 467341 499561 468269
rect 498448 467297 499561 467341
rect 564241 468269 565354 468309
rect 564241 467341 564289 468269
rect 565313 467341 565354 468269
rect 564241 467297 565354 467341
rect 436522 466155 437319 466203
rect 436522 465483 436583 466155
rect 437273 465483 437319 466155
rect 436522 465411 437319 465483
rect 311938 441279 312046 441285
rect 311938 440355 312046 441183
rect 311938 440259 311944 440355
rect 312040 440259 312046 440355
rect 437258 441279 437366 441285
rect 437258 440355 437366 441183
rect 437258 440259 437264 440355
rect 437360 440259 437366 440355
rect 345338 438432 345394 439232
rect 410214 438488 410270 439230
rect 337242 438376 345394 438432
rect 402118 438432 410270 438488
rect 470658 438432 470714 439232
rect 535534 438488 535590 439230
rect 337242 437634 337298 438376
rect 402118 437632 402174 438432
rect 462562 438376 470714 438432
rect 527438 438432 535590 438488
rect 462562 437634 462618 438376
rect 527438 437632 527494 438432
rect 435466 436509 435472 436605
rect 435568 436509 435574 436605
rect 435466 435681 435574 436509
rect 435466 435579 435574 435585
rect 560786 436509 560792 436605
rect 560888 436509 560894 436605
rect 560786 435681 560894 436509
rect 560786 435579 560894 435585
rect 307335 405609 308448 405649
rect 307335 404681 307383 405609
rect 308407 404681 308448 405609
rect 307335 404637 308448 404681
rect 373128 405609 374241 405649
rect 373128 404681 373176 405609
rect 374200 404681 374241 405609
rect 373128 404637 374241 404681
rect 498448 405609 499561 405649
rect 498448 404681 498496 405609
rect 499520 404681 499561 405609
rect 498448 404637 499561 404681
rect 564241 405609 565354 405649
rect 564241 404681 564289 405609
rect 565313 404681 565354 405609
rect 564241 404637 565354 404681
rect 436522 403495 437319 403543
rect 436522 402823 436583 403495
rect 437273 402823 437319 403495
rect 436522 402751 437319 402823
rect 311942 378537 312038 378543
rect 311942 377783 312038 378441
rect 311942 377681 312038 377687
rect 437262 378537 437358 378543
rect 437262 377783 437358 378441
rect 437262 377681 437358 377687
rect 345338 375772 345394 376572
rect 410214 375828 410270 376570
rect 337242 375716 345394 375772
rect 402118 375772 410270 375828
rect 470658 375772 470714 376572
rect 535534 375828 535590 376570
rect 337242 374974 337298 375716
rect 402118 374972 402174 375772
rect 462562 375716 470714 375772
rect 527438 375772 535590 375828
rect 462562 374974 462618 375716
rect 527438 374972 527494 375772
rect 435474 373857 435570 373863
rect 435474 373103 435570 373761
rect 435474 373001 435570 373007
rect 560794 373857 560890 373863
rect 560794 373103 560890 373761
rect 560794 373001 560890 373007
rect 307335 342949 308448 342989
rect 307335 342021 307383 342949
rect 308407 342021 308448 342949
rect 307335 341977 308448 342021
rect 373128 342949 374241 342989
rect 373128 342021 373176 342949
rect 374200 342021 374241 342949
rect 373128 341977 374241 342021
rect 498448 342949 499561 342989
rect 498448 342021 498496 342949
rect 499520 342021 499561 342949
rect 498448 341977 499561 342021
rect 564241 342949 565354 342989
rect 564241 342021 564289 342949
rect 565313 342021 565354 342949
rect 564241 341977 565354 342021
rect 436522 340835 437319 340883
rect 436522 340163 436583 340835
rect 437273 340163 437319 340835
rect 436522 340091 437319 340163
rect 311938 315959 312046 315965
rect 311938 315035 312046 315863
rect 311938 314939 311944 315035
rect 312040 314939 312046 315035
rect 437258 315959 437366 315965
rect 437258 315035 437366 315863
rect 437258 314939 437264 315035
rect 437360 314939 437366 315035
rect 345338 313112 345394 313912
rect 410214 313168 410270 313910
rect 337242 313056 345394 313112
rect 402118 313112 410270 313168
rect 470658 313112 470714 313912
rect 535534 313168 535590 313910
rect 337242 312314 337298 313056
rect 402118 312312 402174 313112
rect 462562 313056 470714 313112
rect 527438 313112 535590 313168
rect 462562 312314 462618 313056
rect 527438 312312 527494 313112
rect 435466 311189 435472 311285
rect 435568 311189 435574 311285
rect 435466 310361 435574 311189
rect 435466 310259 435574 310265
rect 560786 311189 560792 311285
rect 560888 311189 560894 311285
rect 560786 310361 560894 311189
rect 560786 310259 560894 310265
rect 307335 280289 308448 280329
rect 307335 279361 307383 280289
rect 308407 279361 308448 280289
rect 307335 279317 308448 279361
rect 373128 280289 374241 280329
rect 373128 279361 373176 280289
rect 374200 279361 374241 280289
rect 373128 279317 374241 279361
rect 498448 280289 499561 280329
rect 498448 279361 498496 280289
rect 499520 279361 499561 280289
rect 498448 279317 499561 279361
rect 564241 280289 565354 280329
rect 564241 279361 564289 280289
rect 565313 279361 565354 280289
rect 564241 279317 565354 279361
rect 436522 278175 437319 278223
rect 436522 277503 436583 278175
rect 437273 277503 437319 278175
rect 436522 277431 437319 277503
rect 311942 253217 312038 253223
rect 311942 252463 312038 253121
rect 311942 252361 312038 252367
rect 437262 253217 437358 253223
rect 437262 252463 437358 253121
rect 437262 252361 437358 252367
rect 345338 250452 345394 251252
rect 410214 250508 410270 251250
rect 337242 250396 345394 250452
rect 402118 250452 410270 250508
rect 470658 250452 470714 251252
rect 535534 250508 535590 251250
rect 337242 249654 337298 250396
rect 402118 249652 402174 250452
rect 462562 250396 470714 250452
rect 527438 250452 535590 250508
rect 462562 249654 462618 250396
rect 527438 249652 527494 250452
rect 435474 248537 435570 248543
rect 435474 247783 435570 248441
rect 435474 247681 435570 247687
rect 560794 248537 560890 248543
rect 560794 247783 560890 248441
rect 560794 247681 560890 247687
rect 307335 217629 308448 217669
rect 307335 216701 307383 217629
rect 308407 216701 308448 217629
rect 307335 216657 308448 216701
rect 373128 217629 374241 217669
rect 373128 216701 373176 217629
rect 374200 216701 374241 217629
rect 373128 216657 374241 216701
rect 498448 217629 499561 217669
rect 498448 216701 498496 217629
rect 499520 216701 499561 217629
rect 498448 216657 499561 216701
rect 564241 217629 565354 217669
rect 564241 216701 564289 217629
rect 565313 216701 565354 217629
rect 564241 216657 565354 216701
rect 436522 215515 437319 215563
rect 436522 214843 436583 215515
rect 437273 214843 437319 215515
rect 436522 214771 437319 214843
rect 311938 190639 312046 190645
rect 311938 189715 312046 190543
rect 311938 189619 311944 189715
rect 312040 189619 312046 189715
rect 437258 190639 437366 190645
rect 437258 189715 437366 190543
rect 437258 189619 437264 189715
rect 437360 189619 437366 189715
rect 345338 187792 345394 188592
rect 410214 187848 410270 188590
rect 337242 187736 345394 187792
rect 402118 187792 410270 187848
rect 470658 187792 470714 188592
rect 535534 187848 535590 188590
rect 337242 186994 337298 187736
rect 402118 186992 402174 187792
rect 462562 187736 470714 187792
rect 527438 187792 535590 187848
rect 462562 186994 462618 187736
rect 527438 186992 527494 187792
rect 435466 185869 435472 185965
rect 435568 185869 435574 185965
rect 435466 185041 435574 185869
rect 435466 184939 435574 184945
rect 560786 185869 560792 185965
rect 560888 185869 560894 185965
rect 560786 185041 560894 185869
rect 560786 184939 560894 184945
rect 307335 154969 308448 155009
rect 307335 154041 307383 154969
rect 308407 154041 308448 154969
rect 307335 153997 308448 154041
rect 373128 154969 374241 155009
rect 373128 154041 373176 154969
rect 374200 154041 374241 154969
rect 373128 153997 374241 154041
rect 498448 154969 499561 155009
rect 498448 154041 498496 154969
rect 499520 154041 499561 154969
rect 498448 153997 499561 154041
rect 564241 154969 565354 155009
rect 564241 154041 564289 154969
rect 565313 154041 565354 154969
rect 564241 153997 565354 154041
rect 436522 152855 437319 152903
rect 436522 152183 436583 152855
rect 437273 152183 437319 152855
rect 436522 152111 437319 152183
rect 311942 127897 312038 127903
rect 311942 127143 312038 127801
rect 311942 127041 312038 127047
rect 437262 127897 437358 127903
rect 437262 127143 437358 127801
rect 437262 127041 437358 127047
rect 345338 125132 345394 125932
rect 410214 125188 410270 125930
rect 337242 125076 345394 125132
rect 402118 125132 410270 125188
rect 470658 125132 470714 125932
rect 535534 125188 535590 125930
rect 337242 124334 337298 125076
rect 402118 124332 402174 125132
rect 462562 125076 470714 125132
rect 527438 125132 535590 125188
rect 462562 124334 462618 125076
rect 527438 124332 527494 125132
rect 561662 124574 561667 124630
rect 435474 123217 435570 123223
rect 435474 122463 435570 123121
rect 435474 122361 435570 122367
rect 560794 123217 560890 123223
rect 560794 122463 560890 123121
rect 561670 122766 561880 122821
rect 560794 122361 560890 122367
rect 307335 92309 308448 92349
rect 307335 91381 307383 92309
rect 308407 91381 308448 92309
rect 307335 91337 308448 91381
rect 373128 92309 374241 92349
rect 373128 91381 373176 92309
rect 374200 91381 374241 92309
rect 373128 91337 374241 91381
rect 498448 92309 499561 92349
rect 498448 91381 498496 92309
rect 499520 91381 499561 92309
rect 498448 91337 499561 91381
rect 436522 90195 437319 90243
rect 436522 89523 436583 90195
rect 437273 89523 437319 90195
rect 436522 89451 437319 89523
rect 311938 65319 312046 65325
rect 311938 64395 312046 65223
rect 311938 64299 311944 64395
rect 312040 64299 312046 64395
rect 561824 63757 561880 122766
rect 564241 92309 565354 92349
rect 564241 91381 564289 92309
rect 565313 91381 565354 92309
rect 564241 91337 565354 91381
rect 537485 63701 561880 63757
rect 345338 62180 345394 63272
rect 410214 62528 410270 63270
rect 470658 62528 470714 63272
rect 410214 62472 470714 62528
rect 501310 62223 501366 62541
rect 535534 62502 535590 63270
rect 535494 62483 535637 62502
rect 535494 62378 535511 62483
rect 535627 62378 535637 62483
rect 535494 62356 535637 62378
rect 345447 62194 345574 62202
rect 345447 62180 345461 62194
rect 345338 62124 345461 62180
rect 345447 62092 345461 62124
rect 345563 62092 345574 62194
rect 501310 62167 536675 62223
rect 345447 62080 345574 62092
rect 536619 61997 536675 62167
rect 537485 62046 537541 63701
rect 537443 62028 537586 62046
rect 536580 61973 536723 61997
rect 536580 61868 536597 61973
rect 536713 61868 536723 61973
rect 537443 61923 537460 62028
rect 537576 61923 537586 62028
rect 537443 61900 537586 61923
rect 536580 61851 536723 61868
<< via2 >>
rect 102991 653874 103145 654016
rect 105567 653899 105721 654041
rect 108323 653914 108477 654056
rect 113667 653773 113821 653915
rect 102332 651892 102424 651972
rect 95870 644429 96526 646722
rect 101376 636822 101456 636922
rect 103956 636822 104036 636922
rect 96598 634384 96722 634523
rect 109266 636822 109356 636902
rect 112026 636832 112116 636912
rect 115455 637499 115663 638077
rect 114606 636742 114696 636822
rect 96605 634106 96729 634245
rect 96613 633846 96737 633985
rect 119296 646120 119388 646200
rect 119128 645916 119228 646006
rect 119968 645938 120060 646018
rect 127470 642700 128350 642780
rect 123830 642040 123960 642610
rect 131500 642060 131630 642630
rect 127460 641880 128340 641960
rect 119290 640060 119382 640140
rect 119128 639582 119228 639672
rect 120010 639576 120102 639656
rect 126070 636580 126950 636660
rect 129100 635900 129230 636470
rect 126080 635680 126960 635760
rect 96620 633561 96744 633700
rect 119292 633678 119384 633758
rect 119138 633304 119220 633388
rect 119936 633142 120028 633222
rect 126290 630500 127170 630580
rect 129170 629840 129300 630410
rect 126290 629690 127170 629770
rect 119308 627140 119400 627220
rect 119136 626806 119218 626890
rect 119918 626702 120010 626782
rect 126540 623980 127420 624060
rect 128820 623320 128950 623890
rect 126540 623170 127420 623250
rect 119296 620764 119388 620844
rect 119142 620400 119224 620484
rect 119950 620294 120042 620374
rect 128380 619330 128860 619460
rect 131940 618240 132070 618810
rect 128380 617580 128860 617710
rect 119304 614284 119396 614364
rect 119142 613974 119224 614058
rect 119978 613888 120070 613968
rect 128030 611880 128510 612010
rect 131590 610790 131720 611360
rect 128030 610130 128510 610260
rect 119308 607978 119400 608058
rect 119138 607592 119220 607676
rect 119914 607480 120006 607560
rect 128160 605830 128640 605960
rect 131720 604640 131850 605310
rect 128160 603980 128640 604110
rect 119296 601686 119388 601766
rect 119144 601222 119226 601306
rect 119958 601104 120050 601184
rect 127960 599570 128440 599700
rect 131520 598280 131650 599050
rect 127960 597620 128440 597750
rect 119336 594154 119428 594234
rect 119104 593672 119186 593756
rect 119926 593546 120018 593626
rect 118700 592800 118790 592880
rect 127920 592020 128400 592150
rect 131480 590630 131610 591500
rect 127920 589970 128400 590100
rect 119306 584602 119398 584682
rect 119144 584130 119226 584214
rect 120128 584028 120220 584108
rect 118740 583260 118830 583340
rect 128380 583040 128860 583170
rect 132890 581950 133020 582520
rect 128376 581292 128856 581422
rect 119318 575480 119410 575560
rect 119138 575094 119220 575178
rect 120036 575004 120128 575084
rect 118780 574240 118870 574320
rect 128420 574020 128900 574150
rect 132930 572830 133060 573500
rect 128416 572172 128896 572302
rect 119374 567962 119466 568042
rect 119134 567426 119216 567510
rect 119994 567302 120086 567382
rect 118730 566570 118820 566650
rect 128370 566350 128850 566480
rect 132880 565060 133010 565830
rect 128376 564402 128856 564532
rect 119314 561344 119406 561424
rect 119124 560864 119206 560948
rect 120034 560874 120126 560954
rect 118730 560030 118820 560110
rect 128370 559810 128850 559940
rect 132880 558420 133010 559290
rect 128376 557762 128856 557892
rect 119350 554560 119442 554640
rect 119132 553978 119214 554062
rect 120078 553952 120170 554032
rect 118800 553200 118890 553280
rect 128840 552980 129370 553110
rect 133900 551890 134030 552460
rect 128846 551232 129326 551362
rect 119336 546942 119428 547022
rect 119128 546408 119210 546492
rect 120170 546368 120262 546448
rect 118800 545630 118890 545710
rect 128840 545410 129370 545540
rect 133900 544120 134030 544890
rect 128866 543462 129346 543592
rect 119318 538902 119410 538982
rect 119132 538390 119214 538474
rect 120046 538344 120138 538424
rect 118770 537570 118860 537650
rect 128810 537350 129340 537480
rect 133870 535860 134000 536830
rect 128826 535212 129306 535342
rect 307383 530001 308407 530929
rect 373176 530001 374200 530929
rect 498496 530001 499520 530929
rect 564289 530001 565313 530929
rect 436583 528143 437273 528815
rect 307383 467341 308407 468269
rect 373176 467341 374200 468269
rect 498496 467341 499520 468269
rect 564289 467341 565313 468269
rect 436583 465483 437273 466155
rect 307383 404681 308407 405609
rect 373176 404681 374200 405609
rect 498496 404681 499520 405609
rect 564289 404681 565313 405609
rect 436583 402823 437273 403495
rect 307383 342021 308407 342949
rect 373176 342021 374200 342949
rect 498496 342021 499520 342949
rect 564289 342021 565313 342949
rect 436583 340163 437273 340835
rect 307383 279361 308407 280289
rect 373176 279361 374200 280289
rect 498496 279361 499520 280289
rect 564289 279361 565313 280289
rect 436583 277503 437273 278175
rect 307383 216701 308407 217629
rect 373176 216701 374200 217629
rect 498496 216701 499520 217629
rect 564289 216701 565313 217629
rect 436583 214843 437273 215515
rect 307383 154041 308407 154969
rect 373176 154041 374200 154969
rect 498496 154041 499520 154969
rect 564289 154041 565313 154969
rect 436583 152183 437273 152855
rect 307383 91381 308407 92309
rect 373176 91381 374200 92309
rect 498496 91381 499520 92309
rect 436583 89523 437273 90195
rect 564289 91381 565313 92309
rect 535511 62378 535627 62483
rect 345461 62092 345563 62194
rect 536597 61868 536713 61973
rect 537460 61923 537576 62028
<< metal3 >>
rect 102943 655665 119850 655888
rect 102943 654048 103166 655665
rect 105519 655069 118084 655292
rect 105519 654073 105742 655069
rect 108275 654751 108498 654762
rect 108275 654528 117621 654751
rect 108275 654088 108498 654528
rect 102943 654016 103167 654048
rect 102943 653874 102991 654016
rect 103145 653874 103167 654016
rect 102943 653840 103167 653874
rect 105519 654041 105743 654073
rect 105519 653899 105567 654041
rect 105721 653899 105743 654041
rect 105519 653865 105743 653899
rect 108275 654056 108499 654088
rect 108275 653914 108323 654056
rect 108477 653914 108499 654056
rect 108275 653880 108499 653914
rect 113619 654082 117223 654305
rect 113619 653947 113842 654082
rect 113619 653915 113843 653947
rect 113619 653773 113667 653915
rect 113821 653773 113843 653915
rect 113619 653739 113843 653773
rect 98156 652322 101536 652442
rect 91826 646722 96646 646822
rect 91826 644429 95870 646722
rect 96526 644429 96646 646722
rect 91826 644292 96646 644429
rect 80486 638952 96096 639623
rect 80486 636805 94762 638952
rect 95963 636805 96096 638952
rect 80486 636526 96096 636805
rect 80486 561767 83583 636526
rect 96238 634901 96419 634924
rect 96238 634789 96262 634901
rect 96392 634789 96419 634901
rect 95614 634577 95795 634600
rect 95614 634561 95638 634577
rect 95604 634465 95638 634561
rect 95768 634465 95795 634577
rect 95604 634427 95795 634465
rect 96238 634541 96419 634789
rect 96578 634541 96766 634556
rect 96238 634523 96766 634541
rect 95604 634263 95785 634427
rect 96238 634384 96598 634523
rect 96722 634384 96766 634523
rect 96238 634360 96766 634384
rect 96578 634358 96766 634360
rect 96585 634263 96771 634278
rect 95604 634245 96771 634263
rect 95604 634106 96605 634245
rect 96729 634106 96771 634245
rect 95604 634082 96771 634106
rect 96593 634014 96779 634018
rect 95307 633985 96779 634014
rect 95307 633846 96613 633985
rect 96737 633846 96779 633985
rect 95307 633833 96779 633846
rect 95307 633710 95488 633833
rect 96593 633822 96779 633833
rect 96600 633718 96786 633733
rect 95307 633687 95504 633710
rect 95307 633575 95347 633687
rect 95477 633575 95504 633687
rect 95307 633537 95504 633575
rect 96024 633700 96786 633718
rect 96024 633561 96620 633700
rect 96744 633561 96786 633700
rect 96024 633537 96786 633561
rect 95307 633536 95488 633537
rect 96024 633370 96205 633537
rect 96024 633347 96222 633370
rect 96024 633235 96065 633347
rect 96195 633235 96222 633347
rect 96024 633197 96222 633235
rect 98156 568192 98276 652322
rect 102308 651972 102442 651990
rect 102308 651892 102332 651972
rect 102424 651892 102442 651972
rect 102308 651870 102442 651892
rect 116169 649874 116863 649994
rect 98496 648514 101676 648634
rect 98496 568832 98616 648514
rect 116218 646066 116588 646186
rect 98946 644434 101736 644554
rect 98946 569482 99066 644434
rect 99526 640626 101596 640746
rect 99526 570122 99646 640626
rect 115410 638077 115696 638189
rect 115410 637499 115455 638077
rect 115663 637499 115696 638077
rect 115410 637416 115696 637499
rect 101366 636922 101486 636942
rect 101366 636822 101376 636922
rect 101456 636822 101486 636922
rect 101366 636762 101486 636822
rect 103946 636922 104066 636942
rect 103946 636822 103956 636922
rect 104036 636822 104066 636922
rect 103946 636762 104066 636822
rect 99996 636642 101486 636762
rect 103826 636642 104066 636762
rect 109226 636902 109386 636942
rect 109226 636822 109266 636902
rect 109356 636822 109386 636902
rect 99996 571082 100116 636642
rect 103826 636372 103946 636642
rect 100516 636252 103946 636372
rect 100516 575172 100636 636252
rect 109226 584513 109386 636822
rect 111986 636912 112146 636952
rect 111986 636832 112026 636912
rect 112116 636832 112146 636912
rect 111986 593467 112146 636832
rect 114566 636822 114726 636862
rect 114566 636742 114606 636822
rect 114696 636742 114726 636822
rect 114566 600951 114726 636742
rect 116035 611288 116155 642106
rect 116468 618099 116588 646066
rect 116743 623455 116863 649874
rect 117000 631630 117223 654082
rect 117398 638053 117621 654528
rect 117861 644410 118084 655069
rect 119627 646971 119850 655665
rect 118893 646748 119850 646971
rect 118893 646024 119116 646748
rect 119272 646200 119406 646218
rect 119272 646120 119296 646200
rect 119388 646120 119406 646200
rect 119272 646098 119406 646120
rect 118893 646006 119261 646024
rect 118893 645916 119128 646006
rect 119228 645916 119261 646006
rect 119944 646018 120078 646036
rect 119944 645938 119968 646018
rect 120060 645938 120078 646018
rect 119944 645916 120078 645938
rect 118893 645801 119261 645916
rect 117861 644187 119894 644410
rect 119266 640140 119400 640158
rect 119266 640060 119290 640140
rect 119382 640060 119400 640140
rect 119266 640038 119400 640060
rect 119671 639854 119894 644187
rect 127460 642780 128360 642790
rect 127460 642700 127470 642780
rect 128350 642700 128360 642780
rect 127460 642690 128360 642700
rect 131470 642630 131660 642650
rect 123800 642610 123990 642630
rect 123800 642040 123830 642610
rect 123960 642040 123990 642610
rect 131470 642060 131500 642630
rect 131630 642060 131660 642630
rect 131470 642040 131660 642060
rect 123800 642020 123990 642040
rect 127450 641960 128350 641970
rect 127450 641880 127460 641960
rect 128340 641880 128350 641960
rect 127450 641870 128350 641880
rect 119106 639690 119898 639854
rect 119106 639672 119246 639690
rect 119106 639582 119128 639672
rect 119228 639582 119246 639672
rect 119106 639562 119246 639582
rect 119986 639656 120120 639674
rect 119986 639576 120010 639656
rect 120102 639576 120120 639656
rect 119986 639554 120120 639576
rect 117398 637830 119850 638053
rect 119268 633758 119402 633776
rect 119268 633678 119292 633758
rect 119384 633678 119402 633758
rect 119268 633656 119402 633678
rect 119627 633510 119850 637830
rect 126060 636660 126960 636670
rect 126060 636580 126070 636660
rect 126950 636580 126960 636660
rect 126060 636570 126960 636580
rect 129070 636470 129260 636490
rect 129070 635900 129100 636470
rect 129230 635900 129260 636470
rect 129070 635880 129260 635900
rect 126070 635760 126970 635770
rect 126070 635680 126080 635760
rect 126960 635680 126970 635760
rect 126070 635670 126970 635680
rect 576114 634523 580914 644396
rect 119061 633388 119850 633510
rect 119061 633304 119138 633388
rect 119220 633304 119850 633388
rect 119061 633287 119850 633304
rect 564550 634247 580914 634523
rect 119912 633222 120046 633240
rect 119912 633142 119936 633222
rect 120028 633142 120046 633222
rect 119912 633120 120046 633142
rect 117000 631407 120093 631630
rect 119284 627220 119418 627238
rect 119284 627140 119308 627220
rect 119400 627140 119418 627220
rect 119284 627118 119418 627140
rect 119870 627010 120093 631407
rect 126280 630580 127180 630590
rect 126280 630500 126290 630580
rect 127170 630500 127180 630580
rect 126280 630490 127180 630500
rect 129140 630410 129330 630430
rect 129140 629840 129170 630410
rect 129300 629840 129330 630410
rect 129140 629820 129330 629840
rect 564550 630082 564780 634247
rect 569092 630082 580914 634247
rect 126280 629770 127180 629780
rect 126280 629690 126290 629770
rect 127170 629690 127180 629770
rect 564550 629723 580914 630082
rect 126280 629680 127180 629690
rect 119124 626906 120093 627010
rect 119122 626905 120093 626906
rect 119122 626902 120058 626905
rect 119122 626890 119236 626902
rect 119122 626806 119136 626890
rect 119218 626806 119236 626890
rect 119122 626792 119236 626806
rect 119894 626782 120028 626800
rect 119894 626702 119918 626782
rect 120010 626702 120028 626782
rect 119894 626680 120028 626702
rect 126530 624060 127430 624070
rect 126530 623980 126540 624060
rect 127420 623980 127430 624060
rect 126530 623970 127430 623980
rect 128790 623890 128980 623910
rect 116743 623335 119799 623455
rect 119272 620844 119406 620862
rect 119272 620764 119296 620844
rect 119388 620764 119406 620844
rect 119272 620742 119406 620764
rect 119679 620522 119799 623335
rect 128790 623320 128820 623890
rect 128950 623320 128980 623890
rect 128790 623300 128980 623320
rect 126530 623250 127430 623260
rect 126530 623170 126540 623250
rect 127420 623170 127430 623250
rect 126530 623160 127430 623170
rect 119130 620500 119799 620522
rect 119128 620484 119799 620500
rect 119128 620400 119142 620484
rect 119224 620402 119799 620484
rect 119224 620400 119242 620402
rect 119128 620386 119242 620400
rect 119926 620374 120060 620392
rect 119926 620294 119950 620374
rect 120042 620294 120060 620374
rect 119926 620272 120060 620294
rect 128360 619460 128880 619480
rect 128360 619330 128380 619460
rect 128860 619330 128880 619460
rect 128360 619310 128880 619330
rect 131910 618810 132100 618830
rect 131910 618240 131940 618810
rect 132070 618240 132100 618810
rect 131910 618220 132100 618240
rect 116468 617979 119800 618099
rect 119280 614364 119414 614382
rect 119280 614284 119304 614364
rect 119396 614284 119414 614364
rect 119280 614262 119414 614284
rect 119680 614108 119800 617979
rect 128360 617710 128880 617730
rect 128360 617580 128380 617710
rect 128860 617580 128880 617710
rect 128360 617560 128880 617580
rect 119134 614074 119800 614108
rect 119128 614058 119800 614074
rect 119128 613974 119142 614058
rect 119224 613988 119800 614058
rect 119224 613974 119242 613988
rect 119128 613960 119242 613974
rect 119954 613968 120088 613986
rect 119954 613888 119978 613968
rect 120070 613888 120088 613968
rect 119954 613866 120088 613888
rect 128010 612010 128530 612030
rect 128010 611880 128030 612010
rect 128510 611880 128530 612010
rect 128010 611860 128530 611880
rect 131560 611360 131750 611380
rect 116035 611168 120051 611288
rect 119284 608058 119418 608076
rect 119284 607978 119308 608058
rect 119400 607978 119418 608058
rect 119284 607956 119418 607978
rect 119931 607792 120051 611168
rect 131560 610790 131590 611360
rect 131720 610790 131750 611360
rect 131560 610770 131750 610790
rect 128010 610260 128530 610280
rect 128010 610130 128030 610260
rect 128510 610130 128530 610260
rect 128010 610110 128530 610130
rect 119138 607692 120051 607792
rect 119124 607676 120051 607692
rect 119124 607592 119138 607676
rect 119220 607672 120051 607676
rect 119220 607592 119238 607672
rect 119124 607578 119238 607592
rect 119890 607560 120024 607578
rect 119890 607480 119914 607560
rect 120006 607480 120024 607560
rect 119890 607458 120024 607480
rect 128140 605960 128660 605980
rect 128140 605830 128160 605960
rect 128640 605830 128660 605960
rect 128140 605810 128660 605830
rect 131690 605310 131880 605330
rect 131690 604640 131720 605310
rect 131850 604640 131880 605310
rect 131690 604620 131880 604640
rect 128140 604110 128660 604130
rect 128140 603980 128160 604110
rect 128640 603980 128660 604110
rect 128140 603960 128660 603980
rect 119272 601766 119406 601784
rect 119272 601686 119296 601766
rect 119388 601686 119406 601766
rect 119272 601664 119406 601686
rect 117544 601322 119234 601324
rect 117544 601306 119244 601322
rect 117544 601222 119144 601306
rect 119226 601222 119244 601306
rect 117544 601208 119244 601222
rect 117544 601164 119234 601208
rect 119934 601184 120068 601202
rect 117544 600951 117704 601164
rect 119934 601104 119958 601184
rect 120050 601104 120068 601184
rect 119934 601082 120068 601104
rect 114566 600791 117704 600951
rect 127940 599700 128460 599720
rect 127940 599570 127960 599700
rect 128440 599570 128460 599700
rect 127940 599550 128460 599570
rect 131490 599050 131680 599070
rect 131490 598280 131520 599050
rect 131650 598280 131680 599050
rect 131490 598260 131680 598280
rect 127940 597750 128460 597770
rect 127940 597620 127960 597750
rect 128440 597620 128460 597750
rect 127940 597600 128460 597620
rect 119312 594234 119446 594252
rect 119312 594154 119336 594234
rect 119428 594154 119446 594234
rect 119312 594132 119446 594154
rect 117155 593756 119204 593794
rect 117155 593672 119104 593756
rect 119186 593672 119204 593756
rect 117155 593634 119204 593672
rect 117155 593467 117315 593634
rect 119902 593626 120036 593644
rect 119902 593546 119926 593626
rect 120018 593546 120036 593626
rect 119902 593524 120036 593546
rect 111986 593307 117315 593467
rect 118690 592880 118800 592890
rect 118690 592800 118700 592880
rect 118790 592800 118800 592880
rect 118690 592790 118800 592800
rect 127900 592150 128420 592170
rect 127900 592020 127920 592150
rect 128400 592020 128420 592150
rect 127900 592000 128420 592020
rect 131450 591500 131640 591520
rect 131450 590630 131480 591500
rect 131610 590630 131640 591500
rect 131450 590610 131640 590630
rect 127900 590100 128420 590120
rect 127900 589970 127920 590100
rect 128400 589970 128420 590100
rect 127900 589950 128420 589970
rect 561623 587024 581434 587032
rect 561616 586920 581434 587024
rect 119282 584682 119416 584700
rect 119282 584602 119306 584682
rect 119398 584602 119416 584682
rect 119282 584580 119416 584602
rect 109226 584353 119248 584513
rect 119088 584214 119248 584353
rect 119088 584146 119144 584214
rect 119130 584130 119144 584146
rect 119226 584146 119248 584214
rect 119226 584130 119244 584146
rect 119130 584116 119244 584130
rect 120104 584108 120238 584126
rect 120104 584028 120128 584108
rect 120220 584028 120238 584108
rect 120104 584006 120238 584028
rect 118730 583340 118840 583350
rect 118730 583260 118740 583340
rect 118830 583260 118840 583340
rect 118730 583250 118840 583260
rect 128360 583170 128880 583190
rect 128360 583040 128380 583170
rect 128860 583040 128880 583170
rect 128360 583020 128880 583040
rect 132860 582520 133050 582540
rect 132860 581950 132890 582520
rect 133020 581950 133050 582520
rect 132860 581930 133050 581950
rect 128360 581422 128880 581440
rect 128360 581292 128376 581422
rect 128856 581420 128880 581422
rect 128360 581290 128380 581292
rect 128860 581290 128880 581420
rect 128360 581270 128880 581290
rect 119294 575560 119428 575578
rect 119294 575480 119318 575560
rect 119410 575480 119428 575560
rect 119294 575458 119428 575480
rect 119124 575178 119238 575194
rect 119124 575172 119138 575178
rect 100516 575094 119138 575172
rect 119220 575094 119238 575178
rect 100516 575080 119238 575094
rect 120012 575084 120146 575102
rect 100516 575052 119228 575080
rect 120012 575004 120036 575084
rect 120128 575004 120146 575084
rect 120012 574982 120146 575004
rect 118770 574320 118880 574330
rect 118770 574240 118780 574320
rect 118870 574240 118880 574320
rect 118770 574230 118880 574240
rect 128400 574150 128920 574170
rect 128400 574020 128420 574150
rect 128900 574020 128920 574150
rect 128400 574000 128920 574020
rect 132900 573500 133090 573520
rect 132900 572830 132930 573500
rect 133060 572830 133090 573500
rect 132900 572810 133090 572830
rect 128400 572302 128920 572320
rect 128400 572172 128416 572302
rect 128896 572300 128920 572302
rect 128400 572170 128420 572172
rect 128900 572170 128920 572300
rect 128400 572150 128920 572170
rect 99996 570962 101556 571082
rect 99526 570002 100726 570122
rect 98946 569362 100096 569482
rect 98496 568712 99576 568832
rect 98156 568072 99156 568192
rect 68295 558670 83583 561767
rect 99036 539312 99156 568072
rect 99456 547822 99576 568712
rect 99976 555492 100096 569362
rect 100606 561722 100726 570002
rect 101436 567832 101556 570962
rect 119350 568042 119484 568060
rect 119350 567962 119374 568042
rect 119466 567962 119484 568042
rect 119350 567940 119484 567962
rect 101436 567712 119242 567832
rect 119122 567526 119242 567712
rect 119120 567510 119242 567526
rect 119120 567426 119134 567510
rect 119216 567426 119242 567510
rect 119120 567412 119242 567426
rect 119122 567386 119242 567412
rect 119970 567382 120104 567400
rect 119970 567302 119994 567382
rect 120086 567302 120104 567382
rect 119970 567280 120104 567302
rect 118720 566650 118830 566660
rect 118720 566570 118730 566650
rect 118820 566570 118830 566650
rect 118720 566560 118830 566570
rect 128350 566480 128870 566500
rect 128350 566350 128370 566480
rect 128850 566350 128870 566480
rect 128350 566330 128870 566350
rect 132850 565830 133040 565850
rect 132850 565060 132880 565830
rect 133010 565060 133040 565830
rect 132850 565040 133040 565060
rect 561616 565026 561736 586920
rect 311096 564906 561736 565026
rect 128350 564532 128870 564550
rect 128350 564530 128376 564532
rect 128350 564400 128370 564530
rect 128856 564402 128870 564532
rect 128850 564400 128870 564402
rect 128350 564380 128870 564400
rect 100606 561602 117532 561722
rect 117412 560966 117532 561602
rect 119290 561424 119424 561442
rect 119290 561344 119314 561424
rect 119406 561344 119424 561424
rect 119290 561322 119424 561344
rect 117412 560948 119232 560966
rect 117412 560864 119124 560948
rect 119206 560864 119232 560948
rect 117412 560846 119232 560864
rect 120010 560954 120144 560972
rect 120010 560874 120034 560954
rect 120126 560874 120144 560954
rect 120010 560852 120144 560874
rect 118720 560110 118830 560120
rect 118720 560030 118730 560110
rect 118820 560030 118830 560110
rect 118720 560020 118830 560030
rect 128350 559940 128870 559960
rect 128350 559810 128370 559940
rect 128850 559810 128870 559940
rect 128350 559790 128870 559810
rect 132850 559290 133040 559310
rect 132850 558420 132880 559290
rect 133010 558420 133040 559290
rect 132850 558400 133040 558420
rect 128350 557892 128870 557910
rect 128350 557890 128376 557892
rect 128350 557760 128370 557890
rect 128856 557762 128870 557892
rect 128850 557760 128870 557762
rect 128350 557740 128870 557760
rect 99976 555372 117718 555492
rect 117598 554060 117718 555372
rect 119326 554640 119460 554658
rect 119326 554560 119350 554640
rect 119442 554560 119460 554640
rect 119326 554538 119460 554560
rect 119118 554062 119232 554078
rect 119118 554060 119132 554062
rect 117598 553978 119132 554060
rect 119214 553978 119232 554062
rect 117598 553964 119232 553978
rect 120054 554032 120188 554050
rect 117598 553940 119218 553964
rect 120054 553952 120078 554032
rect 120170 553952 120188 554032
rect 120054 553930 120188 553952
rect 118790 553280 118900 553290
rect 118790 553200 118800 553280
rect 118890 553200 118900 553280
rect 118790 553190 118900 553200
rect 128820 553110 129390 553130
rect 128820 552980 128840 553110
rect 129370 552980 129390 553110
rect 128820 552960 129390 552980
rect 133870 552460 134060 552480
rect 133870 551890 133900 552460
rect 134030 551890 134060 552460
rect 133870 551870 134060 551890
rect 311096 551812 311216 564906
rect 436296 551812 436416 564906
rect 311096 551692 311896 551812
rect 436296 551692 437216 551812
rect 128820 551362 129390 551380
rect 128820 551360 128846 551362
rect 129326 551360 129390 551362
rect 128820 551230 128840 551360
rect 129370 551230 129390 551360
rect 128820 551210 129390 551230
rect 99456 547702 117660 547822
rect 117540 546462 117660 547702
rect 119312 547022 119446 547040
rect 119312 546942 119336 547022
rect 119428 546942 119446 547022
rect 119312 546920 119446 546942
rect 119114 546492 119228 546508
rect 119114 546462 119128 546492
rect 117540 546408 119128 546462
rect 119210 546408 119228 546492
rect 117540 546394 119228 546408
rect 120146 546448 120280 546466
rect 117540 546342 119222 546394
rect 120146 546368 120170 546448
rect 120262 546368 120280 546448
rect 120146 546346 120280 546368
rect 118790 545710 118900 545720
rect 118790 545630 118800 545710
rect 118890 545630 118900 545710
rect 118790 545620 118900 545630
rect 128820 545540 129390 545560
rect 128820 545410 128840 545540
rect 129370 545410 129390 545540
rect 128820 545390 129390 545410
rect 133870 544890 134060 544910
rect 133870 544120 133900 544890
rect 134030 544120 134060 544890
rect 133870 544100 134060 544120
rect 128820 543592 129390 543610
rect 128820 543590 128866 543592
rect 129346 543590 129390 543592
rect 128820 543460 128840 543590
rect 129370 543460 129390 543590
rect 128820 543440 129390 543460
rect 99036 539192 117740 539312
rect 117620 538462 117740 539192
rect 119294 538982 119428 539000
rect 119294 538902 119318 538982
rect 119410 538902 119428 538982
rect 119294 538880 119428 538902
rect 119118 538474 119232 538490
rect 119118 538462 119132 538474
rect 117620 538390 119132 538462
rect 119214 538462 119232 538474
rect 119214 538390 119238 538462
rect 117620 538342 119238 538390
rect 120022 538424 120156 538442
rect 120022 538344 120046 538424
rect 120138 538344 120156 538424
rect 120022 538322 120156 538344
rect 118760 537650 118870 537660
rect 118760 537570 118770 537650
rect 118860 537570 118870 537650
rect 118760 537560 118870 537570
rect 128790 537480 129360 537500
rect 128790 537350 128810 537480
rect 129340 537350 129360 537480
rect 128790 537330 129360 537350
rect 133840 536830 134030 536850
rect 133840 535860 133870 536830
rect 134000 535860 134030 536830
rect 133840 535840 134030 535860
rect 128790 535342 129360 535350
rect 128790 535330 128826 535342
rect 129306 535330 129360 535342
rect 128790 535200 128810 535330
rect 129340 535200 129360 535330
rect 128790 535180 129360 535200
rect 307335 530929 308448 530969
rect 307335 530001 307383 530929
rect 308407 530001 308448 530929
rect 307335 529957 308448 530001
rect 8842 512111 9055 512117
rect 8842 511892 9055 511898
rect 8892 507908 9004 511892
rect -1910 507796 9004 507908
rect 311096 489152 311216 551692
rect 373128 530929 374241 530969
rect 373128 530001 373176 530929
rect 374200 530001 374241 530929
rect 373128 529957 374241 530001
rect 436296 513152 436416 551692
rect 498448 530929 499561 530969
rect 498448 530001 498496 530929
rect 499520 530001 499561 530929
rect 498448 529957 499561 530001
rect 436522 528815 437319 528863
rect 436522 528143 436583 528815
rect 437273 528143 437319 528815
rect 436522 528071 437319 528143
rect 561616 513152 561736 564906
rect 564241 530929 565354 530969
rect 564241 530001 564289 530929
rect 565313 530001 565354 530929
rect 564241 529957 565354 530001
rect 435616 513032 436416 513152
rect 560936 513032 561736 513152
rect 436296 489152 436416 513032
rect 311096 489032 311896 489152
rect 436296 489032 437216 489152
rect 307335 468269 308448 468309
rect 307335 467341 307383 468269
rect 308407 467341 308448 468269
rect 307335 467297 308448 467341
rect 14566 466634 14770 466640
rect 14566 466424 14770 466430
rect 14612 464686 14724 466424
rect -1896 464574 14724 464686
rect 311096 426492 311216 489032
rect 373128 468269 374241 468309
rect 373128 467341 373176 468269
rect 374200 467341 374241 468269
rect 373128 467297 374241 467341
rect 436296 450492 436416 489032
rect 498448 468269 499561 468309
rect 498448 467341 498496 468269
rect 499520 467341 499561 468269
rect 498448 467297 499561 467341
rect 436522 466155 437319 466203
rect 436522 465483 436583 466155
rect 437273 465483 437319 466155
rect 436522 465411 437319 465483
rect 561616 450492 561736 513032
rect 564241 468269 565354 468309
rect 564241 467341 564289 468269
rect 565313 467341 565354 468269
rect 564241 467297 565354 467341
rect 435616 450372 436416 450492
rect 560936 450372 561736 450492
rect 436296 426492 436416 450372
rect 311096 426372 311896 426492
rect 436296 426372 437216 426492
rect 9274 422112 9478 422118
rect 9274 421902 9478 421908
rect 9320 421464 9432 421902
rect -1836 421352 9432 421464
rect 307335 405609 308448 405649
rect 307335 404681 307383 405609
rect 308407 404681 308448 405609
rect 307335 404637 308448 404681
rect 9254 380928 9458 380934
rect 9254 380718 9458 380724
rect 9300 378242 9412 380718
rect -1850 378130 9412 378242
rect 311096 363832 311216 426372
rect 373128 405609 374241 405649
rect 373128 404681 373176 405609
rect 374200 404681 374241 405609
rect 373128 404637 374241 404681
rect 436296 387832 436416 426372
rect 498448 405609 499561 405649
rect 498448 404681 498496 405609
rect 499520 404681 499561 405609
rect 498448 404637 499561 404681
rect 436522 403495 437319 403543
rect 436522 402823 436583 403495
rect 437273 402823 437319 403495
rect 436522 402751 437319 402823
rect 561616 387832 561736 450372
rect 564241 405609 565354 405649
rect 564241 404681 564289 405609
rect 565313 404681 565354 405609
rect 564241 404637 565354 404681
rect 435616 387712 436416 387832
rect 560936 387712 561736 387832
rect 436296 363832 436416 387712
rect 311096 363712 311896 363832
rect 436296 363712 437216 363832
rect 307335 342949 308448 342989
rect 307335 342021 307383 342949
rect 308407 342021 308448 342949
rect 307335 341977 308448 342021
rect 311096 301172 311216 363712
rect 373128 342949 374241 342989
rect 373128 342021 373176 342949
rect 374200 342021 374241 342949
rect 373128 341977 374241 342021
rect 436296 325172 436416 363712
rect 498448 342949 499561 342989
rect 498448 342021 498496 342949
rect 499520 342021 499561 342949
rect 498448 341977 499561 342021
rect 436522 340835 437319 340883
rect 436522 340163 436583 340835
rect 437273 340163 437319 340835
rect 436522 340091 437319 340163
rect 561616 325172 561736 387712
rect 564241 342949 565354 342989
rect 564241 342021 564289 342949
rect 565313 342021 565354 342949
rect 564241 341977 565354 342021
rect 435616 325052 436416 325172
rect 560936 325052 561736 325172
rect 436296 301172 436416 325052
rect 311096 301052 311896 301172
rect 436296 301052 437216 301172
rect 307335 280289 308448 280329
rect 307335 279361 307383 280289
rect 308407 279361 308448 280289
rect 307335 279317 308448 279361
rect 311096 238512 311216 301052
rect 373128 280289 374241 280329
rect 373128 279361 373176 280289
rect 374200 279361 374241 280289
rect 373128 279317 374241 279361
rect 436296 262512 436416 301052
rect 498448 280289 499561 280329
rect 498448 279361 498496 280289
rect 499520 279361 499561 280289
rect 498448 279317 499561 279361
rect 436522 278175 437319 278223
rect 436522 277503 436583 278175
rect 437273 277503 437319 278175
rect 436522 277431 437319 277503
rect 561616 262512 561736 325052
rect 564241 280289 565354 280329
rect 564241 279361 564289 280289
rect 565313 279361 565354 280289
rect 564241 279317 565354 279361
rect 435616 262392 436416 262512
rect 560936 262392 561736 262512
rect 436296 238512 436416 262392
rect 311096 238392 311896 238512
rect 436296 238392 437216 238512
rect 307335 217629 308448 217669
rect 307335 216701 307383 217629
rect 308407 216701 308448 217629
rect 307335 216657 308448 216701
rect 311096 175852 311216 238392
rect 373128 217629 374241 217669
rect 373128 216701 373176 217629
rect 374200 216701 374241 217629
rect 373128 216657 374241 216701
rect 436296 199852 436416 238392
rect 498448 217629 499561 217669
rect 498448 216701 498496 217629
rect 499520 216701 499561 217629
rect 498448 216657 499561 216701
rect 436522 215515 437319 215563
rect 436522 214843 436583 215515
rect 437273 214843 437319 215515
rect 436522 214771 437319 214843
rect 561616 199852 561736 262392
rect 564241 217629 565354 217669
rect 564241 216701 564289 217629
rect 565313 216701 565354 217629
rect 564241 216657 565354 216701
rect 435616 199732 436416 199852
rect 560936 199732 561736 199852
rect 436296 175852 436416 199732
rect 311096 175732 311896 175852
rect 436296 175732 437216 175852
rect 307335 154969 308448 155009
rect 307335 154041 307383 154969
rect 308407 154041 308448 154969
rect 307335 153997 308448 154041
rect 311096 113192 311216 175732
rect 373128 154969 374241 155009
rect 373128 154041 373176 154969
rect 374200 154041 374241 154969
rect 373128 153997 374241 154041
rect 436296 137192 436416 175732
rect 498448 154969 499561 155009
rect 498448 154041 498496 154969
rect 499520 154041 499561 154969
rect 498448 153997 499561 154041
rect 436522 152855 437319 152903
rect 436522 152183 436583 152855
rect 437273 152183 437319 152855
rect 436522 152111 437319 152183
rect 561616 137192 561736 199732
rect 564241 154969 565354 155009
rect 564241 154041 564289 154969
rect 565313 154041 565354 154969
rect 564241 153997 565354 154041
rect 576240 141435 581039 151446
rect 435616 137072 436416 137192
rect 560936 137072 561736 137192
rect 436296 113192 436416 137072
rect 311096 113072 311896 113192
rect 436296 113072 437216 113192
rect 307335 92309 308448 92349
rect 307335 91381 307383 92309
rect 308407 91381 308448 92309
rect 307335 91337 308448 91381
rect 373128 92309 374241 92349
rect 373128 91381 373176 92309
rect 374200 91381 374241 92309
rect 373128 91337 374241 91381
rect 436296 74532 436416 113072
rect 498448 92309 499561 92349
rect 498448 91381 498496 92309
rect 499520 91381 499561 92309
rect 498448 91337 499561 91381
rect 436522 90195 437319 90243
rect 436522 89523 436583 90195
rect 437273 89523 437319 90195
rect 436522 89451 437319 89523
rect 435616 74412 436416 74532
rect 501220 63674 501340 113428
rect 561616 74532 561736 137072
rect 566043 136613 566198 141435
rect 571009 139966 581039 141435
rect 571009 137124 572037 139966
rect 574879 137124 581039 139966
rect 571009 136636 581039 137124
rect 564241 92309 565354 92349
rect 564241 91381 564289 92309
rect 565313 91381 565354 92309
rect 564241 91337 565354 91381
rect 560936 74412 561736 74532
rect 501220 63554 538189 63674
rect 535494 62483 535637 62502
rect 535494 62378 535511 62483
rect 535627 62462 535637 62483
rect 535627 62378 535641 62462
rect 535494 62356 535641 62378
rect 345447 62194 345574 62202
rect 345447 62092 345461 62194
rect 345563 62092 345574 62194
rect 345447 62080 345574 62092
rect 345456 52428 345568 62080
rect 535496 53488 535641 62356
rect 537443 62028 537586 62046
rect 536580 61990 536723 61997
rect 536578 61973 536726 61990
rect 536578 61868 536597 61973
rect 536713 61868 536726 61973
rect 536578 54440 536726 61868
rect 537443 61923 537460 62028
rect 537576 62023 537586 62028
rect 537576 61923 537591 62023
rect 537443 55177 537591 61923
rect 538069 55592 538189 63554
rect 538069 55472 565388 55592
rect 537443 55166 563469 55177
rect 537443 55029 563567 55166
rect 536578 54434 561813 54440
rect 536578 54292 561829 54434
rect 535496 53409 560031 53488
rect 535496 53343 560035 53409
rect 345456 52316 556937 52428
rect 556825 2650 556937 52316
rect 559923 8560 560035 53343
rect 561717 13288 561829 54292
rect 563455 18016 563567 55029
rect 565193 22744 565305 55472
rect 565193 22632 581478 22744
rect 563455 17904 581485 18016
rect 561717 13176 581428 13288
rect 559923 8448 581552 8560
rect 556825 2538 581505 2650
<< via3 >>
rect 94762 636805 95963 638952
rect 96262 634789 96392 634901
rect 95638 634465 95768 634577
rect 95347 633575 95477 633687
rect 96065 633235 96195 633347
rect 102332 651892 102424 651972
rect 115455 637499 115663 638077
rect 119296 646120 119388 646200
rect 119968 645938 120060 646018
rect 119290 640060 119382 640140
rect 127470 642700 128350 642780
rect 131500 642060 131630 642630
rect 127460 641880 128340 641960
rect 120010 639576 120102 639656
rect 119292 633678 119384 633758
rect 126070 636580 126950 636660
rect 129100 635900 129230 636470
rect 126080 635680 126960 635760
rect 119936 633142 120028 633222
rect 119308 627140 119400 627220
rect 126290 630500 127170 630580
rect 129170 629840 129300 630410
rect 564780 630082 569092 634247
rect 126290 629690 127170 629770
rect 119918 626702 120010 626782
rect 126540 623980 127420 624060
rect 119296 620764 119388 620844
rect 128820 623320 128950 623890
rect 126540 623170 127420 623250
rect 119950 620294 120042 620374
rect 128380 619330 128860 619460
rect 131940 618240 132070 618810
rect 119304 614284 119396 614364
rect 128380 617580 128860 617710
rect 119978 613888 120070 613968
rect 128030 611880 128510 612010
rect 119308 607978 119400 608058
rect 131590 610790 131720 611360
rect 128030 610130 128510 610260
rect 119914 607480 120006 607560
rect 128160 605830 128640 605960
rect 131720 604640 131850 605310
rect 128160 603980 128640 604110
rect 119296 601686 119388 601766
rect 119958 601104 120050 601184
rect 127960 599570 128440 599700
rect 131520 598280 131650 599050
rect 127960 597620 128440 597750
rect 119336 594154 119428 594234
rect 119926 593546 120018 593626
rect 118700 592800 118790 592880
rect 127920 592020 128400 592150
rect 131480 590630 131610 591500
rect 127920 589970 128400 590100
rect 119306 584602 119398 584682
rect 120128 584028 120220 584108
rect 118740 583260 118830 583340
rect 128380 583040 128860 583170
rect 132890 581950 133020 582520
rect 128376 581292 128856 581422
rect 128856 581292 128860 581420
rect 128380 581290 128860 581292
rect 119318 575480 119410 575560
rect 120036 575004 120128 575084
rect 118780 574240 118870 574320
rect 128420 574020 128900 574150
rect 132930 572830 133060 573500
rect 128420 572172 128896 572300
rect 128896 572172 128900 572300
rect 128420 572170 128900 572172
rect 119374 567962 119466 568042
rect 119994 567302 120086 567382
rect 118730 566570 118820 566650
rect 128370 566350 128850 566480
rect 132880 565060 133010 565830
rect 128370 564402 128376 564530
rect 128376 564402 128850 564530
rect 128370 564400 128850 564402
rect 119314 561344 119406 561424
rect 120034 560874 120126 560954
rect 118730 560030 118820 560110
rect 128370 559810 128850 559940
rect 132880 558420 133010 559290
rect 128370 557762 128376 557890
rect 128376 557762 128850 557890
rect 128370 557760 128850 557762
rect 119350 554560 119442 554640
rect 120078 553952 120170 554032
rect 118800 553200 118890 553280
rect 128840 552980 129370 553110
rect 133900 551890 134030 552460
rect 128840 551232 128846 551360
rect 128846 551232 129326 551360
rect 129326 551232 129370 551360
rect 128840 551230 129370 551232
rect 119336 546942 119428 547022
rect 120170 546368 120262 546448
rect 118800 545630 118890 545710
rect 128840 545410 129370 545540
rect 133900 544120 134030 544890
rect 128840 543462 128866 543590
rect 128866 543462 129346 543590
rect 129346 543462 129370 543590
rect 128840 543460 129370 543462
rect 119318 538902 119410 538982
rect 120046 538344 120138 538424
rect 118770 537570 118860 537650
rect 128810 537350 129340 537480
rect 133870 535860 134000 536830
rect 128810 535212 128826 535330
rect 128826 535212 129306 535330
rect 129306 535212 129340 535330
rect 128810 535200 129340 535212
rect 307383 530001 308407 530929
rect 8842 511898 9055 512111
rect 373176 530001 374200 530929
rect 498496 530001 499520 530929
rect 436583 528143 437273 528815
rect 564289 530001 565313 530929
rect 307383 467341 308407 468269
rect 14566 466430 14770 466634
rect 373176 467341 374200 468269
rect 498496 467341 499520 468269
rect 436583 465483 437273 466155
rect 564289 467341 565313 468269
rect 9274 421908 9478 422112
rect 307383 404681 308407 405609
rect 9254 380724 9458 380928
rect 373176 404681 374200 405609
rect 498496 404681 499520 405609
rect 436583 402823 437273 403495
rect 564289 404681 565313 405609
rect 307383 342021 308407 342949
rect 373176 342021 374200 342949
rect 498496 342021 499520 342949
rect 436583 340163 437273 340835
rect 564289 342021 565313 342949
rect 307383 279361 308407 280289
rect 373176 279361 374200 280289
rect 498496 279361 499520 280289
rect 436583 277503 437273 278175
rect 564289 279361 565313 280289
rect 307383 216701 308407 217629
rect 373176 216701 374200 217629
rect 498496 216701 499520 217629
rect 436583 214843 437273 215515
rect 564289 216701 565313 217629
rect 307383 154041 308407 154969
rect 373176 154041 374200 154969
rect 498496 154041 499520 154969
rect 436583 152183 437273 152855
rect 564289 154041 565313 154969
rect 307383 91381 308407 92309
rect 373176 91381 374200 92309
rect 498496 91381 499520 92309
rect 436583 89523 437273 90195
rect 572037 137124 574879 139966
rect 564289 91381 565313 92309
<< metal4 >>
rect 102298 652002 102454 652004
rect 102298 651972 120893 652002
rect 102298 651892 102332 651972
rect 102424 651892 120893 651972
rect 102298 651856 120893 651892
rect 117846 646342 118109 646345
rect 117846 646200 119418 646342
rect 117846 646120 119296 646200
rect 119388 646120 119418 646200
rect 117846 646088 119418 646120
rect 117844 646082 119418 646088
rect 117844 640237 118110 646082
rect 119934 646018 120090 646050
rect 119934 646017 119968 646018
rect 119917 645938 119968 646017
rect 120060 646017 120090 646018
rect 120747 646017 120893 651856
rect 120060 645938 120893 646017
rect 119917 645871 120893 645938
rect 117844 640140 119447 640237
rect 117844 640060 119290 640140
rect 119382 640060 119447 640140
rect 117844 639971 119447 640060
rect 94565 638952 96078 639083
rect 94565 636805 94762 638952
rect 95963 638211 96078 638952
rect 117844 638211 118110 639971
rect 119976 639697 120132 639716
rect 120747 639697 120893 645871
rect 127390 643550 141652 644590
rect 127390 642780 128430 643550
rect 127390 642700 127470 642780
rect 128350 642700 128430 642780
rect 127390 642620 128430 642700
rect 131470 642630 146061 642650
rect 131470 642060 131500 642630
rect 131630 642060 146061 642630
rect 131470 642040 146061 642060
rect 127380 641960 128420 642040
rect 127380 641880 127460 641960
rect 128340 641880 128420 641960
rect 127380 641190 128420 641880
rect 127380 640150 150501 641190
rect 119976 639656 120893 639697
rect 119976 639576 120010 639656
rect 120102 639576 120893 639656
rect 119976 639551 120893 639576
rect 119976 639538 120132 639551
rect 95963 638077 118110 638211
rect 95963 637499 115455 638077
rect 115663 637499 118110 638077
rect 95963 637386 118110 637499
rect 95963 637364 118109 637386
rect 95963 636805 96078 637364
rect 94565 636665 96078 636805
rect 93849 634943 96423 634950
rect 93849 634901 96427 634943
rect 93849 634789 96262 634901
rect 96392 634789 96427 634901
rect 93849 634751 96427 634789
rect 93849 634737 96423 634751
rect 93849 512114 94062 634737
rect 8755 512111 94062 512114
rect 8755 511901 8842 512111
rect 8841 511898 8842 511901
rect 9055 511901 94062 512111
rect 94214 634577 95809 634625
rect 94214 634465 95638 634577
rect 95768 634465 95809 634577
rect 94214 634421 95809 634465
rect 9055 511898 9056 511901
rect 8841 511897 9056 511898
rect 94214 466641 94418 634421
rect 117846 633874 118109 637364
rect 117846 633758 119429 633874
rect 14509 466634 94418 466641
rect 14509 466437 14566 466634
rect 14565 466430 14566 466437
rect 14770 466437 94418 466634
rect 94620 633687 95512 633743
rect 94620 633575 95347 633687
rect 95477 633575 95512 633687
rect 94620 633539 95512 633575
rect 14770 466430 14771 466437
rect 14565 466429 14771 466430
rect 94620 422139 94824 633539
rect 95314 633537 95512 633539
rect 117846 633678 119292 633758
rect 119384 633678 119429 633758
rect 117846 633611 119429 633678
rect 9229 422112 94824 422139
rect 9229 421935 9274 422112
rect 9273 421908 9274 421935
rect 9478 421935 94824 422112
rect 95025 633347 96233 633396
rect 95025 633235 96065 633347
rect 96195 633235 96233 633347
rect 95025 633192 96233 633235
rect 9478 421908 9479 421935
rect 9273 421907 9479 421908
rect 9253 380928 9459 380929
rect 9253 380916 9254 380928
rect 9207 380724 9254 380916
rect 9458 380916 9459 380928
rect 95025 380916 95229 633192
rect 117846 627322 118109 633611
rect 119902 633235 120058 633282
rect 120747 633235 120893 639551
rect 125990 637800 141492 638840
rect 125990 636660 127030 637800
rect 125990 636580 126070 636660
rect 126950 636580 127030 636660
rect 125990 636500 127030 636580
rect 129640 636490 145501 636500
rect 129070 636470 145501 636490
rect 129070 635900 129100 636470
rect 129230 635900 145501 636470
rect 129070 635880 145501 635900
rect 126000 635760 127040 635840
rect 126000 635680 126080 635760
rect 126960 635680 127040 635760
rect 126000 634770 127040 635680
rect 126000 633730 150401 634770
rect 126000 633720 128140 633730
rect 553830 634247 569349 634522
rect 119902 633222 120893 633235
rect 119902 633142 119936 633222
rect 120028 633142 120893 633222
rect 119902 633104 120893 633142
rect 119955 633089 120893 633104
rect 117846 627280 119429 627322
rect 117846 627220 119430 627280
rect 117846 627140 119308 627220
rect 119400 627140 119430 627220
rect 117846 627102 119430 627140
rect 117846 627059 119429 627102
rect 117846 620952 118109 627059
rect 119884 626813 120040 626842
rect 120747 626813 120893 633089
rect 126206 631972 127246 632072
rect 126206 630932 141512 631972
rect 126210 630580 127250 630932
rect 126210 630500 126290 630580
rect 127170 630500 127250 630580
rect 126210 630420 127250 630500
rect 129496 630430 145621 630432
rect 129140 630410 145621 630430
rect 129140 629840 129170 630410
rect 129300 629840 145621 630410
rect 126210 629770 127250 629840
rect 129140 629822 145621 629840
rect 129140 629820 129530 629822
rect 126210 629690 126290 629770
rect 127170 629690 127250 629770
rect 126210 629442 127250 629690
rect 126206 629432 127250 629442
rect 126206 629352 127256 629432
rect 553830 630082 564780 634247
rect 569092 630082 569349 634247
rect 553830 629723 569349 630082
rect 126206 628312 139586 629352
rect 126206 628302 127246 628312
rect 138546 628302 139586 628312
rect 138546 627262 150261 628302
rect 119884 626782 120893 626813
rect 119884 626702 119918 626782
rect 120010 626702 120893 626782
rect 119884 626667 120893 626702
rect 119884 626664 120040 626667
rect 117846 620904 119417 620952
rect 117846 620844 119418 620904
rect 117846 620764 119296 620844
rect 119388 620764 119418 620844
rect 117846 620726 119418 620764
rect 117846 620689 119417 620726
rect 117846 614472 118109 620689
rect 119916 620403 120072 620434
rect 120747 620403 120893 626667
rect 126466 624512 141752 625552
rect 126466 624420 127506 624512
rect 126460 624242 127506 624420
rect 126460 624060 127500 624242
rect 126460 623980 126540 624060
rect 127420 623980 127500 624060
rect 126460 623930 127500 623980
rect 129076 623910 145841 623912
rect 128790 623890 145841 623910
rect 128790 623320 128820 623890
rect 128950 623320 145841 623890
rect 128790 623302 145841 623320
rect 128790 623300 129180 623302
rect 126460 623250 127500 623270
rect 126460 623170 126540 623250
rect 127420 623170 127500 623250
rect 126460 622932 127500 623170
rect 126456 622910 127500 622932
rect 126456 622662 127496 622910
rect 147251 623302 147266 623912
rect 126456 621622 150351 622662
rect 151541 621622 151596 622662
rect 119916 620374 120893 620403
rect 119916 620294 119950 620374
rect 120042 620294 120893 620374
rect 119916 620257 120893 620294
rect 119916 620256 120072 620257
rect 117846 614364 119435 614472
rect 117846 614284 119304 614364
rect 119396 614284 119435 614364
rect 117846 614209 119435 614284
rect 117846 608153 118109 614209
rect 119944 614015 120100 614028
rect 120747 614015 120893 620257
rect 128360 620200 141532 620720
rect 128360 619460 128880 620200
rect 128360 619330 128380 619460
rect 128860 619330 128880 619460
rect 128360 619310 128880 619330
rect 131910 618810 146031 618830
rect 131910 618680 131940 618810
rect 131900 618400 131940 618680
rect 131910 618240 131940 618400
rect 132070 618240 146031 618810
rect 131910 618220 146031 618240
rect 147441 618220 151341 618830
rect 128360 617710 128880 617730
rect 128360 617580 128380 617710
rect 128860 617580 128880 617710
rect 128360 616910 128880 617580
rect 128360 616390 150297 616910
rect 119944 613968 120893 614015
rect 119944 613888 119978 613968
rect 120070 613888 120893 613968
rect 119944 613869 120893 613888
rect 119944 613850 120100 613869
rect 117846 608058 119435 608153
rect 117846 607978 119308 608058
rect 119400 607978 119435 608058
rect 117846 607890 119435 607978
rect 117846 601857 118109 607890
rect 119880 607585 120036 607620
rect 120747 607585 120893 613869
rect 128010 612750 141662 613270
rect 128010 612010 128530 612750
rect 128010 611880 128030 612010
rect 128510 611880 128530 612010
rect 128010 611860 128530 611880
rect 131560 611360 145711 611380
rect 131560 611230 131590 611360
rect 131550 610950 131590 611230
rect 131560 610790 131590 610950
rect 131720 610790 145711 611360
rect 131560 610770 145711 610790
rect 128010 610260 128530 610280
rect 128010 610130 128030 610260
rect 128510 610130 128530 610260
rect 128010 609460 128530 610130
rect 128010 608940 150781 609460
rect 119880 607560 120893 607585
rect 119880 607480 119914 607560
rect 120006 607480 120893 607560
rect 119880 607442 120893 607480
rect 119885 607439 120893 607442
rect 117846 601766 119419 601857
rect 117846 601686 119296 601766
rect 119388 601686 119419 601766
rect 117846 601594 119419 601686
rect 117846 594396 118109 601594
rect 119924 601207 120080 601244
rect 120747 601207 120893 607439
rect 128140 606700 141692 607220
rect 128140 605960 128660 606700
rect 128140 605830 128160 605960
rect 128640 605830 128660 605960
rect 128140 605810 128660 605830
rect 131690 605310 145951 605330
rect 131690 605180 131720 605310
rect 131680 604800 131720 605180
rect 131690 604640 131720 604800
rect 131850 604640 145951 605310
rect 131690 604620 145951 604640
rect 128140 604110 128660 604130
rect 128140 603980 128160 604110
rect 128640 603980 128660 604110
rect 128140 603310 128660 603980
rect 128140 602790 150561 603310
rect 119924 601184 120893 601207
rect 119924 601104 119958 601184
rect 120050 601104 120893 601184
rect 119924 601066 120893 601104
rect 119945 601061 120893 601066
rect 117846 594234 119459 594396
rect 117846 594154 119336 594234
rect 119428 594154 119459 594234
rect 117846 594133 119459 594154
rect 117846 584823 118109 594133
rect 119302 594116 119458 594133
rect 119892 593627 120048 593686
rect 120747 593627 120893 601061
rect 127940 600440 141912 600960
rect 127940 599700 128460 600440
rect 127940 599570 127960 599700
rect 128440 599570 128460 599700
rect 127940 599550 128460 599570
rect 131490 599050 145831 599070
rect 131490 598920 131520 599050
rect 131480 598440 131520 598920
rect 131490 598280 131520 598440
rect 131650 598280 145831 599050
rect 131490 598260 145831 598280
rect 127940 597750 128460 597770
rect 127940 597620 127960 597750
rect 128440 597620 128460 597750
rect 127940 596950 128460 597620
rect 127940 596430 150541 596950
rect 119892 593626 120893 593627
rect 119892 593546 119926 593626
rect 120018 593546 120893 593626
rect 119892 593508 120893 593546
rect 119917 593481 120893 593508
rect 117846 584682 119433 584823
rect 117846 584602 119306 584682
rect 119398 584602 119433 584682
rect 117846 584560 119433 584602
rect 117846 575662 118109 584560
rect 120094 584121 120250 584168
rect 120747 584121 120893 593481
rect 127900 592890 141642 593410
rect 127900 592150 128420 592890
rect 127900 592020 127920 592150
rect 128400 592020 128420 592150
rect 127900 592000 128420 592020
rect 131450 591500 145491 591520
rect 131450 591370 131480 591500
rect 131440 590790 131480 591370
rect 131450 590630 131480 590790
rect 131610 590630 145491 591500
rect 131450 590610 145491 590630
rect 127900 590100 128420 590120
rect 127900 589970 127920 590100
rect 128400 589970 128420 590100
rect 127900 589300 128420 589970
rect 127900 588780 150591 589300
rect 120094 584108 120893 584121
rect 120094 584028 120128 584108
rect 120220 584028 120893 584108
rect 120094 583990 120893 584028
rect 120117 583975 120893 583990
rect 117846 575560 119463 575662
rect 117846 575480 119318 575560
rect 119410 575480 119463 575560
rect 117846 575399 119463 575480
rect 117846 568173 118109 575399
rect 120002 575111 120158 575144
rect 120747 575111 120893 583975
rect 128360 583910 141742 584430
rect 128360 583170 128880 583910
rect 128360 583040 128380 583170
rect 128860 583040 128880 583170
rect 128360 583020 128880 583040
rect 132860 582520 145731 582540
rect 132860 582390 132890 582520
rect 132850 582110 132890 582390
rect 132860 581950 132890 582110
rect 133020 581950 145731 582520
rect 132860 581930 145731 581950
rect 128360 581422 128880 581440
rect 128360 581292 128376 581422
rect 128856 581420 128880 581422
rect 128360 581290 128380 581292
rect 128860 581290 128880 581420
rect 128360 580620 128880 581290
rect 128360 580100 150461 580620
rect 120002 575084 120893 575111
rect 120002 575004 120036 575084
rect 120128 575004 120893 575084
rect 120002 574966 120893 575004
rect 120025 574965 120893 574966
rect 117846 568042 119511 568173
rect 117846 567962 119374 568042
rect 119466 567962 119511 568042
rect 117846 567910 119511 567962
rect 117846 561496 118109 567910
rect 119960 567431 120116 567442
rect 120747 567431 120893 574965
rect 128400 574890 141712 575410
rect 128400 574150 128920 574890
rect 128400 574020 128420 574150
rect 128900 574020 128920 574150
rect 128400 574000 128920 574020
rect 132900 573500 145541 573520
rect 132900 573370 132930 573500
rect 132890 572990 132930 573370
rect 132900 572830 132930 572990
rect 133060 572830 145541 573500
rect 132900 572810 145541 572830
rect 553830 572876 558629 629723
rect 128400 572300 128920 572320
rect 128400 572170 128420 572300
rect 128900 572170 128920 572300
rect 128400 571500 128920 572170
rect 128400 570980 150541 571500
rect 306139 570550 566055 572876
rect 119953 567382 120893 567431
rect 119953 567302 119994 567382
rect 120086 567302 120893 567382
rect 119953 567285 120893 567302
rect 119960 567264 120116 567285
rect 117846 561424 119469 561496
rect 117846 561344 119314 561424
rect 119406 561344 119469 561424
rect 117846 561233 119469 561344
rect 117846 554790 118109 561233
rect 120000 560975 120156 561014
rect 120747 560975 120893 567285
rect 128350 567220 141472 567740
rect 128350 566480 128870 567220
rect 306139 568077 566216 570550
rect 128350 566350 128370 566480
rect 128850 566350 128870 566480
rect 128350 566330 128870 566350
rect 132850 565830 145711 565850
rect 132850 565700 132880 565830
rect 132840 565220 132880 565700
rect 132850 565060 132880 565220
rect 133010 565060 145711 565830
rect 132850 565040 145711 565060
rect 128350 564530 128870 564550
rect 128350 564400 128370 564530
rect 128850 564400 128870 564530
rect 128350 563730 128870 564400
rect 128350 563210 150391 563730
rect 120000 560954 120893 560975
rect 120000 560874 120034 560954
rect 120126 560874 120893 560954
rect 120000 560836 120893 560874
rect 120011 560829 120893 560836
rect 117846 554640 119493 554790
rect 117846 554560 119350 554640
rect 119442 554560 119493 554640
rect 117846 554527 119493 554560
rect 117846 547122 118109 554527
rect 119316 554522 119472 554527
rect 120044 554039 120200 554092
rect 120747 554039 120893 560829
rect 128350 560680 141692 561200
rect 128350 559940 128870 560680
rect 128350 559810 128370 559940
rect 128850 559810 128870 559940
rect 128350 559790 128870 559810
rect 132850 559290 145561 559310
rect 132850 559160 132880 559290
rect 132840 558580 132880 559160
rect 132850 558420 132880 558580
rect 133010 558420 145561 559290
rect 132850 558400 145561 558420
rect 128350 557890 128870 557910
rect 128350 557760 128370 557890
rect 128850 557760 128870 557890
rect 128350 557090 128870 557760
rect 128350 556570 150491 557090
rect 120044 554032 120893 554039
rect 120044 553952 120078 554032
rect 120170 553952 120893 554032
rect 120044 553914 120893 553952
rect 120055 553893 120893 553914
rect 117846 547022 119483 547122
rect 117846 546942 119336 547022
rect 119428 546942 119483 547022
rect 117846 546859 119483 546942
rect 117846 539060 118109 546859
rect 120136 546448 120292 546508
rect 120136 546433 120170 546448
rect 120127 546368 120170 546433
rect 120262 546433 120292 546448
rect 120747 546433 120893 553893
rect 128820 553850 141832 554370
rect 128820 553110 129390 553850
rect 128820 552980 128840 553110
rect 129370 552980 129390 553110
rect 128820 552960 129390 552980
rect 133870 552460 145711 552480
rect 133870 552330 133900 552460
rect 133860 552050 133900 552330
rect 133870 551890 133900 552050
rect 134030 551890 145711 552460
rect 133870 551870 145711 551890
rect 128820 551360 129390 551380
rect 128820 551230 128840 551360
rect 129370 551230 129390 551360
rect 128820 550560 129390 551230
rect 128820 550040 150511 550560
rect 120262 546368 120893 546433
rect 120127 546287 120893 546368
rect 117846 538982 119497 539060
rect 117846 538902 119318 538982
rect 119410 538902 119497 538982
rect 117846 538797 119497 538902
rect 117846 538367 118109 538797
rect 120012 538437 120168 538484
rect 120747 538437 120893 546287
rect 128820 546280 141712 546800
rect 128820 545540 129390 546280
rect 128820 545410 128840 545540
rect 129370 545410 129390 545540
rect 128820 545390 129390 545410
rect 133870 544890 145591 544910
rect 133870 544760 133900 544890
rect 133860 544280 133900 544760
rect 133870 544120 133900 544280
rect 134030 544120 145591 544890
rect 133870 544100 145591 544120
rect 128820 543590 129390 543610
rect 128820 543460 128840 543590
rect 129370 543460 129390 543590
rect 128820 542790 129390 543460
rect 128820 542270 150391 542790
rect 119995 538424 120893 538437
rect 119995 538344 120046 538424
rect 120138 538344 120893 538424
rect 119995 538291 120893 538344
rect 128790 538220 141572 538740
rect 128790 537480 129360 538220
rect 128790 537350 128810 537480
rect 129340 537350 129360 537480
rect 128790 537330 129360 537350
rect 133840 536830 134920 536850
rect 133840 536700 133870 536830
rect 133830 536020 133870 536700
rect 133840 535860 133870 536020
rect 134000 536760 134920 536830
rect 134000 535860 145801 536760
rect 133840 535840 145801 535860
rect 128790 535330 129360 535350
rect 128790 535200 128810 535330
rect 129340 535200 129360 535330
rect 128790 534530 129360 535200
rect 128790 534010 150511 534530
rect 9458 380724 95229 380916
rect 9207 380712 95229 380724
rect 306543 530929 309310 568077
rect 306543 530001 307383 530929
rect 308407 530001 309310 530929
rect 306543 468269 309310 530001
rect 306543 467341 307383 468269
rect 308407 467341 309310 468269
rect 306543 405609 309310 467341
rect 306543 404681 307383 405609
rect 308407 404681 309310 405609
rect 306543 342949 309310 404681
rect 306543 342021 307383 342949
rect 308407 342021 309310 342949
rect 306543 280289 309310 342021
rect 306543 279361 307383 280289
rect 308407 279361 309310 280289
rect 306543 217629 309310 279361
rect 306543 216701 307383 217629
rect 308407 216701 309310 217629
rect 306543 154969 309310 216701
rect 306543 154041 307383 154969
rect 308407 154041 309310 154969
rect 306543 92309 309310 154041
rect 306543 91381 307383 92309
rect 308407 91381 309310 92309
rect 306543 88965 309310 91381
rect 372336 530929 375103 531840
rect 372336 530001 373176 530929
rect 374200 530001 375103 530929
rect 372336 468269 375103 530001
rect 372336 467341 373176 468269
rect 374200 467341 375103 468269
rect 372336 405609 375103 467341
rect 372336 404681 373176 405609
rect 374200 404681 375103 405609
rect 372336 342949 375103 404681
rect 372336 342021 373176 342949
rect 374200 342021 375103 342949
rect 372336 280289 375103 342021
rect 372336 279361 373176 280289
rect 374200 279361 375103 280289
rect 372336 217629 375103 279361
rect 372336 216701 373176 217629
rect 374200 216701 375103 217629
rect 372336 154969 375103 216701
rect 372336 154041 373176 154969
rect 374200 154041 375103 154969
rect 372336 92309 375103 154041
rect 372336 91381 373176 92309
rect 374200 91381 375103 92309
rect 372336 61795 375103 91381
rect 436473 528815 437380 568077
rect 436473 528143 436583 528815
rect 437273 528143 437380 528815
rect 436473 466155 437380 528143
rect 436473 465483 436583 466155
rect 437273 465483 437380 466155
rect 436473 403495 437380 465483
rect 436473 402823 436583 403495
rect 437273 402823 437380 403495
rect 436473 340835 437380 402823
rect 436473 340163 436583 340835
rect 437273 340163 437380 340835
rect 436473 278175 437380 340163
rect 436473 277503 436583 278175
rect 437273 277503 437380 278175
rect 436473 215515 437380 277503
rect 436473 214843 436583 215515
rect 437273 214843 437380 215515
rect 436473 152855 437380 214843
rect 436473 152183 436583 152855
rect 437273 152183 437380 152855
rect 436473 90195 437380 152183
rect 436473 89523 436583 90195
rect 437273 89523 437380 90195
rect 436473 89385 437380 89523
rect 497656 530929 500423 531840
rect 497656 530001 498496 530929
rect 499520 530001 500423 530929
rect 497656 468269 500423 530001
rect 497656 467341 498496 468269
rect 499520 467341 500423 468269
rect 497656 405609 500423 467341
rect 497656 404681 498496 405609
rect 499520 404681 500423 405609
rect 497656 342949 500423 404681
rect 497656 342021 498496 342949
rect 499520 342021 500423 342949
rect 497656 280289 500423 342021
rect 497656 279361 498496 280289
rect 499520 279361 500423 280289
rect 497656 217629 500423 279361
rect 497656 216701 498496 217629
rect 499520 216701 500423 217629
rect 497656 154969 500423 216701
rect 497656 154041 498496 154969
rect 499520 154041 500423 154969
rect 497656 92309 500423 154041
rect 497656 91381 498496 92309
rect 499520 91381 500423 92309
rect 497656 66275 500423 91381
rect 563449 530929 566216 568077
rect 563449 530001 564289 530929
rect 565313 530001 566216 530929
rect 563449 468269 566216 530001
rect 563449 467341 564289 468269
rect 565313 467341 566216 468269
rect 563449 405609 566216 467341
rect 563449 404681 564289 405609
rect 565313 404681 566216 405609
rect 563449 342949 566216 404681
rect 563449 342021 564289 342949
rect 565313 342021 566216 342949
rect 563449 280289 566216 342021
rect 563449 279361 564289 280289
rect 565313 279361 566216 280289
rect 563449 217629 566216 279361
rect 563449 216701 564289 217629
rect 565313 216701 566216 217629
rect 563449 154969 566216 216701
rect 563449 154041 564289 154969
rect 565313 154041 566216 154969
rect 563449 142311 566216 154041
rect 563449 92309 566198 142311
rect 563449 91381 564289 92309
rect 565313 91381 566198 92309
rect 563449 89001 566198 91381
rect 571860 139966 575029 140225
rect 571860 137124 572037 139966
rect 574879 137124 575029 139966
rect 563449 88965 564573 89001
rect 497656 61795 500428 66275
rect 371426 61781 564573 61795
rect 571860 61781 575029 137124
rect 371426 58612 575029 61781
<< via4 >>
rect 141652 643416 142960 644724
rect 146061 641640 147471 643050
rect 150501 640075 151691 641265
rect 141492 637666 142800 638974
rect 145501 635485 146911 636895
rect 150401 633655 151591 634845
rect 141512 630798 142820 632106
rect 145621 629422 147031 630832
rect 150261 627187 151451 628377
rect 141752 624378 143060 625686
rect 145841 622902 147251 624312
rect 150351 621547 151541 622737
rect 141532 619806 142840 621114
rect 146031 617820 147441 619230
rect 150297 616031 151535 617269
rect 141662 612356 142970 613664
rect 145711 610370 147121 611780
rect 150781 608605 151971 609795
rect 141692 606306 143000 607614
rect 145951 604270 147361 605680
rect 150561 602455 151751 603645
rect 141912 600046 143220 601354
rect 145831 597960 147241 599370
rect 150541 596095 151731 597285
rect 118620 592880 118860 592960
rect 118620 592800 118700 592880
rect 118700 592800 118790 592880
rect 118790 592800 118860 592880
rect 118620 592720 118860 592800
rect 141642 592496 142950 593804
rect 145491 590360 146901 591770
rect 150591 588445 151781 589635
rect 118660 583340 118900 583420
rect 118660 583260 118740 583340
rect 118740 583260 118830 583340
rect 118830 583260 118900 583340
rect 118660 583180 118900 583260
rect 141742 583516 143050 584824
rect 145731 581530 147141 582940
rect 150461 579765 151651 580955
rect 118700 574320 118940 574400
rect 118700 574240 118780 574320
rect 118780 574240 118870 574320
rect 118870 574240 118940 574320
rect 118700 574160 118940 574240
rect 141712 574496 143020 575804
rect 145541 572460 146951 573870
rect 150541 570645 151731 571835
rect 118650 566650 118890 566730
rect 118650 566570 118730 566650
rect 118730 566570 118820 566650
rect 118820 566570 118890 566650
rect 118650 566490 118890 566570
rect 141472 566826 142780 568134
rect 145711 564740 147121 566150
rect 150391 562875 151581 564065
rect 118650 560110 118890 560190
rect 118650 560030 118730 560110
rect 118730 560030 118820 560110
rect 118820 560030 118890 560110
rect 118650 559950 118890 560030
rect 141692 560286 143000 561594
rect 145561 558150 146971 559560
rect 150491 556235 151681 557425
rect 118720 553280 118960 553360
rect 118720 553200 118800 553280
rect 118800 553200 118890 553280
rect 118890 553200 118960 553280
rect 118720 553120 118960 553200
rect 141832 553456 143140 554764
rect 145711 551470 147121 552880
rect 150511 549705 151701 550895
rect 118720 545710 118960 545790
rect 118720 545630 118800 545710
rect 118800 545630 118890 545710
rect 118890 545630 118960 545710
rect 118720 545550 118960 545630
rect 141712 545886 143020 547194
rect 145591 543800 147001 545210
rect 150391 541935 151581 543125
rect 118690 537650 118930 537730
rect 118690 537570 118770 537650
rect 118770 537570 118860 537650
rect 118860 537570 118930 537650
rect 118690 537490 118930 537570
rect 141572 537826 142880 539134
rect 145801 535595 147211 537005
rect 150511 533675 151701 534865
<< metal5 >>
rect 118356 658802 119246 658822
rect 169886 658802 172386 665582
rect 118356 656302 172386 658802
rect 118356 592960 119246 656302
rect 221626 654062 224126 665802
rect 141816 651572 224126 654062
rect 141816 651562 143126 651572
rect 144346 651562 224126 651572
rect 141818 644748 143126 651562
rect 239546 646952 242046 666002
rect 141628 644724 143126 644748
rect 141628 643416 141652 644724
rect 142960 643416 143126 644724
rect 141628 643392 143126 643416
rect 141818 638998 143126 643392
rect 141468 638974 143126 638998
rect 141468 637666 141492 638974
rect 142800 637666 143126 638974
rect 141468 637642 143126 637666
rect 141818 632130 143126 637642
rect 145861 645542 242046 646952
rect 145861 643074 147271 645542
rect 169646 645502 242046 645542
rect 145861 643050 147495 643074
rect 145861 641640 146061 643050
rect 147471 641640 147495 643050
rect 145861 641616 147495 641640
rect 145861 636919 147271 641616
rect 150477 641265 151715 641289
rect 150477 640075 150501 641265
rect 151691 641262 151715 641265
rect 255446 641262 257886 662842
rect 151691 640075 257886 641262
rect 150477 640072 257886 640075
rect 150477 640051 151751 640072
rect 145477 636895 147271 636919
rect 145477 635485 145501 636895
rect 146911 635485 147271 636895
rect 145477 635461 147271 635485
rect 141488 632106 143126 632130
rect 141488 630798 141512 632106
rect 142820 630798 143126 632106
rect 145861 630856 147271 635461
rect 150561 634869 151751 640051
rect 171216 639902 257886 640072
rect 150377 634845 151751 634869
rect 150377 633655 150401 634845
rect 151591 633655 151751 634845
rect 150377 633631 151751 633655
rect 141488 630774 143126 630798
rect 141818 625710 143126 630774
rect 145597 630832 147271 630856
rect 145597 629422 145621 630832
rect 147031 629422 147271 630832
rect 145597 629398 147271 629422
rect 141728 625686 143126 625710
rect 141728 624378 141752 625686
rect 143060 624378 143126 625686
rect 141728 624354 143126 624378
rect 141818 621138 143126 624354
rect 145861 624336 147271 629398
rect 150561 628401 151751 633631
rect 150237 628377 151751 628401
rect 150237 627187 150261 628377
rect 151451 627187 151751 628377
rect 150237 627163 151751 627187
rect 145817 624312 147275 624336
rect 145817 622902 145841 624312
rect 147251 622902 147275 624312
rect 145817 622878 147275 622902
rect 141508 621114 143126 621138
rect 141508 619806 141532 621114
rect 142840 619806 143126 621114
rect 141508 619782 143126 619806
rect 141818 613688 143126 619782
rect 141638 613664 143126 613688
rect 141638 612356 141662 613664
rect 142970 612356 143126 613664
rect 141638 612332 143126 612356
rect 141818 607638 143126 612332
rect 145861 619254 147271 622878
rect 150561 622761 151751 627163
rect 150327 622737 151751 622761
rect 150327 621547 150351 622737
rect 151541 621547 151751 622737
rect 150327 621523 151751 621547
rect 145861 619230 147465 619254
rect 145861 617820 146031 619230
rect 147441 617820 147465 619230
rect 145861 617796 147465 617820
rect 145861 611804 147271 617796
rect 150561 617293 151751 621523
rect 150273 617269 151751 617293
rect 150273 616031 150297 617269
rect 151535 616031 151751 617269
rect 150273 616007 151751 616031
rect 145687 611780 147271 611804
rect 145687 610370 145711 611780
rect 147121 610370 147271 611780
rect 145687 610346 147271 610370
rect 141668 607614 143126 607638
rect 141668 606306 141692 607614
rect 143000 606306 143126 607614
rect 141668 606282 143126 606306
rect 141818 601378 143126 606282
rect 145861 605704 147271 610346
rect 150561 609819 151751 616007
rect 150561 609795 151995 609819
rect 150561 608605 150781 609795
rect 151971 608605 151995 609795
rect 150561 608581 151995 608605
rect 145861 605680 147385 605704
rect 145861 604270 145951 605680
rect 147361 604270 147385 605680
rect 145861 604246 147385 604270
rect 141818 601354 143244 601378
rect 141818 600046 141912 601354
rect 143220 600046 143244 601354
rect 141818 600022 143244 600046
rect 141818 593828 143126 600022
rect 145861 599394 147271 604246
rect 150561 603669 151751 608581
rect 150537 603645 151775 603669
rect 150537 602455 150561 603645
rect 151751 602455 151775 603645
rect 150537 602431 151775 602455
rect 145807 599370 147271 599394
rect 145807 597960 145831 599370
rect 147241 597960 147271 599370
rect 145807 597936 147271 597960
rect 118356 592720 118620 592960
rect 118860 592720 119246 592960
rect 118356 583420 119246 592720
rect 141618 593804 143126 593828
rect 141618 592496 141642 593804
rect 142950 592496 143126 593804
rect 141618 592472 143126 592496
rect 141818 584848 143126 592472
rect 145861 591794 147271 597936
rect 150561 597309 151751 602431
rect 150517 597285 151755 597309
rect 150517 596095 150541 597285
rect 151731 596095 151755 597285
rect 150517 596071 151755 596095
rect 145467 591770 147271 591794
rect 145467 590360 145491 591770
rect 146901 590360 147271 591770
rect 145467 590336 147271 590360
rect 141718 584824 143126 584848
rect 141718 583516 141742 584824
rect 143050 583516 143126 584824
rect 141718 583492 143126 583516
rect 118356 583180 118660 583420
rect 118900 583180 119246 583420
rect 118356 574400 119246 583180
rect 141818 575828 143126 583492
rect 145861 582964 147271 590336
rect 145707 582940 147271 582964
rect 145707 581530 145731 582940
rect 147141 581530 147271 582940
rect 145707 581506 147271 581530
rect 141688 575804 143126 575828
rect 141688 574496 141712 575804
rect 143020 574496 143126 575804
rect 141688 574472 143126 574496
rect 118356 574160 118700 574400
rect 118940 574160 119246 574400
rect 118356 566730 119246 574160
rect 141818 568158 143126 574472
rect 145861 573894 147271 581506
rect 150561 589659 151751 596071
rect 150561 589635 151805 589659
rect 150561 588445 150591 589635
rect 151781 588445 151805 589635
rect 150561 588421 151805 588445
rect 150561 580979 151751 588421
rect 150437 580955 151751 580979
rect 150437 579765 150461 580955
rect 151651 579765 151751 580955
rect 150437 579741 151751 579765
rect 145517 573870 147271 573894
rect 145517 572460 145541 573870
rect 146951 572460 147271 573870
rect 145517 572436 147271 572460
rect 141448 568134 143126 568158
rect 141448 566826 141472 568134
rect 142780 566826 143126 568134
rect 141448 566802 143126 566826
rect 118356 566490 118650 566730
rect 118890 566490 119246 566730
rect 118356 560190 119246 566490
rect 141818 561618 143126 566802
rect 145861 566174 147271 572436
rect 150561 571859 151751 579741
rect 150517 571835 151755 571859
rect 150517 570645 150541 571835
rect 151731 570645 151755 571835
rect 150517 570621 151755 570645
rect 145687 566150 147271 566174
rect 145687 564740 145711 566150
rect 147121 564740 147271 566150
rect 145687 564716 147271 564740
rect 141668 561594 143126 561618
rect 141668 560286 141692 561594
rect 143000 560286 143126 561594
rect 141668 560262 143126 560286
rect 118356 559950 118650 560190
rect 118890 559950 119246 560190
rect 118356 553650 119246 559950
rect 141818 554788 143126 560262
rect 145861 559584 147271 564716
rect 150561 564089 151751 570621
rect 150367 564065 151751 564089
rect 150367 562875 150391 564065
rect 151581 562875 151751 564065
rect 150367 562851 151751 562875
rect 145537 559560 147271 559584
rect 145537 558150 145561 559560
rect 146971 558150 147271 559560
rect 145537 558126 147271 558150
rect 141808 554764 143164 554788
rect 118356 553360 119260 553650
rect 141808 553456 141832 554764
rect 143140 553456 143164 554764
rect 141808 553432 143164 553456
rect 118356 553120 118720 553360
rect 118960 553120 119260 553360
rect 118356 552850 119260 553120
rect 118356 546080 119246 552850
rect 141818 547218 143126 553432
rect 145861 552904 147271 558126
rect 150561 557449 151751 562851
rect 150467 557425 151751 557449
rect 150467 556235 150491 557425
rect 151681 556235 151751 557425
rect 150467 556211 151751 556235
rect 145687 552880 147271 552904
rect 145687 551470 145711 552880
rect 147121 551470 147271 552880
rect 145687 551446 147271 551470
rect 141688 547194 143126 547218
rect 118356 545790 119260 546080
rect 141688 545886 141712 547194
rect 143020 545886 143126 547194
rect 141688 545862 143126 545886
rect 118356 545550 118720 545790
rect 118960 545550 119260 545790
rect 118356 545280 119260 545550
rect 118356 537730 119246 545280
rect 141818 539158 143126 545862
rect 145861 545234 147271 551446
rect 150561 550919 151751 556211
rect 150487 550895 151751 550919
rect 150487 549705 150511 550895
rect 151701 549705 151751 550895
rect 150487 549681 151751 549705
rect 145567 545210 147271 545234
rect 145567 543800 145591 545210
rect 147001 543800 147271 545210
rect 145567 543776 147271 543800
rect 141548 539134 143126 539158
rect 141548 537826 141572 539134
rect 142880 537826 143126 539134
rect 141548 537802 143126 537826
rect 118356 537490 118690 537730
rect 118930 537490 119246 537730
rect 118356 535532 119246 537490
rect 141818 537408 143126 537802
rect 145861 537029 147271 543776
rect 150561 543149 151751 549681
rect 150367 543125 151751 543149
rect 150367 541935 150391 543125
rect 151581 541935 151751 543125
rect 150367 541911 151751 541935
rect 145777 537005 147271 537029
rect 145777 535595 145801 537005
rect 147211 535595 147271 537005
rect 145777 535571 147271 535595
rect 145861 535057 147271 535571
rect 150561 534889 151751 541911
rect 150487 534865 151751 534889
rect 150487 533675 150511 534865
rect 151701 533675 151751 534865
rect 150487 533651 151751 533675
rect 150561 532687 151751 533651
use shift_reg  shift_reg_4 ./shift_reg
timestamp 1636908413
transform 1 0 311096 0 1 62472
box 0 0 60516 62660
use shift_reg  shift_reg_5
timestamp 1636908413
transform 1 0 311096 0 1 125132
box 0 0 60516 62660
use shift_reg  shift_reg_34
timestamp 1636908413
transform -1 0 436416 0 -1 125132
box 0 0 60516 62660
use shift_reg  shift_reg_35
timestamp 1636908413
transform -1 0 436416 0 -1 187792
box 0 0 60516 62660
use shift_reg  shift_reg_12
timestamp 1636908413
transform 1 0 436416 0 1 62472
box 0 0 60516 62660
use shift_reg  shift_reg_13
timestamp 1636908413
transform 1 0 436416 0 1 125132
box 0 0 60516 62660
use shift_reg  shift_reg_32
timestamp 1636908413
transform -1 0 561736 0 -1 187792
box 0 0 60516 62660
use shift_reg  shift_reg_33
timestamp 1636908413
transform -1 0 561736 0 -1 125132
box 0 0 60516 62660
use shift_reg  shift_reg_6
timestamp 1636908413
transform 1 0 311096 0 1 187792
box 0 0 60516 62660
use shift_reg  shift_reg_30
timestamp 1636908413
transform -1 0 436416 0 -1 250452
box 0 0 60516 62660
use shift_reg  shift_reg_14
timestamp 1636908413
transform 1 0 436416 0 1 187792
box 0 0 60516 62660
use shift_reg  shift_reg_28
timestamp 1636908413
transform -1 0 561736 0 -1 250452
box 0 0 60516 62660
use shift_reg  shift_reg_7
timestamp 1636908413
transform 1 0 311096 0 1 250452
box 0 0 60516 62660
use shift_reg  shift_reg_31
timestamp 1636908413
transform -1 0 436416 0 -1 313112
box 0 0 60516 62660
use shift_reg  shift_reg_15
timestamp 1636908413
transform 1 0 436416 0 1 250452
box 0 0 60516 62660
use shift_reg  shift_reg_29
timestamp 1636908413
transform -1 0 561736 0 -1 313112
box 0 0 60516 62660
use shift_reg  shift_reg_8
timestamp 1636908413
transform 1 0 311096 0 1 313112
box 0 0 60516 62660
use shift_reg  shift_reg_9
timestamp 1636908413
transform 1 0 311096 0 1 375772
box 0 0 60516 62660
use shift_reg  shift_reg_25
timestamp 1636908413
transform -1 0 436416 0 -1 375772
box 0 0 60516 62660
use shift_reg  shift_reg_26
timestamp 1636908413
transform -1 0 436416 0 -1 438432
box 0 0 60516 62660
use shift_reg  shift_reg_16
timestamp 1636908413
transform 1 0 436416 0 1 313112
box 0 0 60516 62660
use shift_reg  shift_reg_17
timestamp 1636908413
transform 1 0 436416 0 1 375772
box 0 0 60516 62660
use shift_reg  shift_reg_22
timestamp 1636908413
transform -1 0 561736 0 -1 375772
box 0 0 60516 62660
use shift_reg  shift_reg_23
timestamp 1636908413
transform -1 0 561736 0 -1 438432
box 0 0 60516 62660
use shift_reg  shift_reg_10
timestamp 1636908413
transform 1 0 311096 0 1 438432
box 0 0 60516 62660
use shift_reg  shift_reg_27
timestamp 1636908413
transform -1 0 436416 0 -1 501092
box 0 0 60516 62660
use shift_reg  shift_reg_18
timestamp 1636908413
transform 1 0 436416 0 1 438432
box 0 0 60516 62660
use shift_reg  shift_reg_24
timestamp 1636908413
transform -1 0 561736 0 -1 501092
box 0 0 60516 62660
use shift_reg  shift_reg_11
timestamp 1636908413
transform 1 0 311096 0 1 501092
box 0 0 60516 62660
use shift_reg  shift_reg_21
timestamp 1636908413
transform -1 0 436416 0 -1 563752
box 0 0 60516 62660
use shift_reg  shift_reg_19
timestamp 1636908413
transform 1 0 436416 0 1 501092
box 0 0 60516 62660
use shift_reg  shift_reg_20
timestamp 1636908413
transform -1 0 561736 0 -1 563752
box 0 0 60516 62660
use switch-small  switch-small_5
timestamp 1640659972
transform 1 0 -10820 0 1 43090
box 129220 556910 131680 558120
use switch-small  switch-small_3
timestamp 1640659972
transform 1 0 -10820 0 1 68690
box 129220 556910 131680 558120
use switch-small  switch-small_2
timestamp 1640659972
transform 1 0 -10820 0 1 75090
box 129220 556910 131680 558120
use switch-small  switch-small_4
timestamp 1640659972
transform 1 0 -10820 0 1 49490
box 129220 556910 131680 558120
use switch-small  switch-small_6
timestamp 1640659972
transform 1 0 -10820 0 1 55890
box 129220 556910 131680 558120
use switch-small  switch-small_7
timestamp 1640659972
transform 1 0 -10820 0 1 62290
box 129220 556910 131680 558120
use switch-small  switch-small_1
timestamp 1640659972
transform 1 0 -10820 0 1 81490
box 129220 556910 131680 558120
use switch-small  switch-small_0
timestamp 1640659972
transform 1 0 -10820 0 1 87890
box 129220 556910 131680 558120
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 83096 0 1 686690
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 82782 0 1 686690
box -38 -48 314 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 83594 0 1 686690
box -38 -48 1510 592
use analog_switch_decoder  analog_switch_decoder_0 analog_switch_decoder
timestamp 1640660022
transform 1 0 101350 0 1 636810
box 0 0 15020 17164
use ring-osc-flat  ring-osc-flat_0 ../../sky-radtol
timestamp 1640269035
transform 1 0 81064 0 1 686642
box -396 -544 1728 640
<< labels >>
rlabel comment s 115242 640074 115242 640074 6 decap_3
rlabel comment s 115242 641162 115242 641162 6 decap_3
rlabel comment s 115242 642250 115242 642250 6 decap_3
rlabel comment s 115242 643338 115242 643338 6 decap_3
rlabel comment s 115242 644426 115242 644426 6 decap_3
rlabel comment s 115242 645514 115242 645514 6 decap_3
rlabel comment s 115242 646602 115242 646602 6 decap_3
rlabel comment s 115242 647690 115242 647690 6 decap_3
rlabel comment s 115242 648778 115242 648778 6 decap_3
rlabel comment s 115242 649866 115242 649866 6 decap_3
rlabel comment s 115242 650954 115242 650954 6 decap_3
rlabel comment s 370436 65736 370436 65736 6 decap_3
rlabel comment s 370436 66824 370436 66824 6 decap_3
rlabel comment s 370436 67912 370436 67912 6 decap_3
rlabel comment s 370436 69000 370436 69000 6 decap_3
rlabel comment s 370436 70088 370436 70088 6 decap_3
rlabel comment s 370436 71176 370436 71176 6 decap_3
rlabel comment s 370436 72264 370436 72264 6 decap_3
rlabel comment s 370436 73352 370436 73352 6 decap_3
rlabel comment s 370436 74440 370436 74440 6 decap_3
rlabel comment s 370436 75528 370436 75528 6 decap_3
rlabel comment s 370436 76616 370436 76616 6 decap_3
rlabel comment s 370436 77704 370436 77704 6 decap_3
rlabel comment s 370436 78792 370436 78792 6 decap_3
rlabel comment s 370436 79880 370436 79880 6 decap_3
rlabel comment s 370436 80968 370436 80968 6 decap_3
rlabel comment s 370436 82056 370436 82056 6 decap_3
rlabel comment s 370436 83144 370436 83144 6 decap_3
rlabel comment s 370436 84232 370436 84232 6 decap_3
rlabel comment s 370436 85320 370436 85320 6 decap_3
rlabel comment s 370436 86408 370436 86408 6 decap_3
rlabel comment s 370436 87496 370436 87496 6 decap_3
rlabel comment s 370436 88584 370436 88584 6 decap_3
rlabel comment s 370436 89672 370436 89672 6 decap_3
rlabel comment s 370436 90760 370436 90760 6 decap_3
rlabel comment s 370436 91848 370436 91848 6 decap_3
rlabel comment s 370436 92936 370436 92936 6 decap_3
rlabel comment s 370436 94024 370436 94024 6 decap_3
rlabel comment s 370436 95112 370436 95112 6 decap_3
rlabel comment s 370436 96200 370436 96200 6 decap_3
rlabel comment s 370436 97288 370436 97288 6 decap_3
rlabel comment s 370436 98376 370436 98376 6 decap_3
rlabel comment s 370436 99464 370436 99464 6 decap_3
rlabel comment s 370436 100552 370436 100552 6 decap_3
rlabel comment s 370436 101640 370436 101640 6 decap_3
rlabel comment s 370436 102728 370436 102728 6 decap_3
rlabel comment s 370436 103816 370436 103816 6 decap_3
rlabel comment s 370436 104904 370436 104904 6 decap_3
rlabel comment s 370436 105992 370436 105992 6 decap_3
rlabel comment s 370436 107080 370436 107080 6 decap_3
rlabel comment s 370436 108168 370436 108168 6 decap_3
rlabel comment s 370436 109256 370436 109256 6 decap_3
rlabel comment s 370436 110344 370436 110344 6 decap_3
rlabel comment s 370436 111432 370436 111432 6 decap_3
rlabel comment s 370436 112520 370436 112520 6 decap_3
rlabel comment s 370436 113608 370436 113608 6 decap_3
rlabel comment s 370436 114696 370436 114696 6 decap_3
rlabel comment s 370436 115784 370436 115784 6 decap_3
rlabel comment s 370436 116872 370436 116872 6 decap_3
rlabel comment s 370436 117960 370436 117960 6 decap_3
rlabel comment s 370436 119048 370436 119048 6 decap_3
rlabel comment s 370436 120136 370436 120136 6 decap_3
rlabel comment s 370436 121224 370436 121224 6 decap_3
rlabel comment s 370436 122312 370436 122312 6 decap_3
rlabel comment s 370436 128396 370436 128396 6 decap_3
rlabel comment s 370436 129484 370436 129484 6 decap_3
rlabel comment s 370436 130572 370436 130572 6 decap_3
rlabel comment s 370436 131660 370436 131660 6 decap_3
rlabel comment s 370436 132748 370436 132748 6 decap_3
rlabel comment s 370436 133836 370436 133836 6 decap_3
rlabel comment s 370436 134924 370436 134924 6 decap_3
rlabel comment s 370436 136012 370436 136012 6 decap_3
rlabel comment s 370436 137100 370436 137100 6 decap_3
rlabel comment s 370436 138188 370436 138188 6 decap_3
rlabel comment s 370436 139276 370436 139276 6 decap_3
rlabel comment s 370436 140364 370436 140364 6 decap_3
rlabel comment s 370436 141452 370436 141452 6 decap_3
rlabel comment s 370436 142540 370436 142540 6 decap_3
rlabel comment s 370436 143628 370436 143628 6 decap_3
rlabel comment s 370436 144716 370436 144716 6 decap_3
rlabel comment s 370436 145804 370436 145804 6 decap_3
rlabel comment s 370436 146892 370436 146892 6 decap_3
rlabel comment s 370436 147980 370436 147980 6 decap_3
rlabel comment s 370436 149068 370436 149068 6 decap_3
rlabel comment s 370436 150156 370436 150156 6 decap_3
rlabel comment s 370436 151244 370436 151244 6 decap_3
rlabel comment s 370436 152332 370436 152332 6 decap_3
rlabel comment s 370436 153420 370436 153420 6 decap_3
rlabel comment s 370436 154508 370436 154508 6 decap_3
rlabel comment s 370436 155596 370436 155596 6 decap_3
rlabel comment s 370436 156684 370436 156684 6 decap_3
rlabel comment s 370436 157772 370436 157772 6 decap_3
rlabel comment s 370436 158860 370436 158860 6 decap_3
rlabel comment s 370436 159948 370436 159948 6 decap_3
rlabel comment s 370436 161036 370436 161036 6 decap_3
rlabel comment s 370436 162124 370436 162124 6 decap_3
rlabel comment s 370436 163212 370436 163212 6 decap_3
rlabel comment s 370436 164300 370436 164300 6 decap_3
rlabel comment s 370436 165388 370436 165388 6 decap_3
rlabel comment s 370436 166476 370436 166476 6 decap_3
rlabel comment s 370436 167564 370436 167564 6 decap_3
rlabel comment s 370436 168652 370436 168652 6 decap_3
rlabel comment s 370436 169740 370436 169740 6 decap_3
rlabel comment s 370436 170828 370436 170828 6 decap_3
rlabel comment s 370436 171916 370436 171916 6 decap_3
rlabel comment s 370436 173004 370436 173004 6 decap_3
rlabel comment s 370436 174092 370436 174092 6 decap_3
rlabel comment s 370436 175180 370436 175180 6 decap_3
rlabel comment s 370436 176268 370436 176268 6 decap_3
rlabel comment s 370436 177356 370436 177356 6 decap_3
rlabel comment s 370436 178444 370436 178444 6 decap_3
rlabel comment s 370436 179532 370436 179532 6 decap_3
rlabel comment s 370436 180620 370436 180620 6 decap_3
rlabel comment s 370436 181708 370436 181708 6 decap_3
rlabel comment s 370436 182796 370436 182796 6 decap_3
rlabel comment s 370436 183884 370436 183884 6 decap_3
rlabel comment s 370436 184972 370436 184972 6 decap_3
rlabel comment s 370436 191056 370436 191056 6 decap_3
rlabel comment s 370436 192144 370436 192144 6 decap_3
rlabel comment s 370436 193232 370436 193232 6 decap_3
rlabel comment s 370436 194320 370436 194320 6 decap_3
rlabel comment s 370436 195408 370436 195408 6 decap_3
rlabel comment s 370436 196496 370436 196496 6 decap_3
rlabel comment s 370436 197584 370436 197584 6 decap_3
rlabel comment s 370436 198672 370436 198672 6 decap_3
rlabel comment s 370436 199760 370436 199760 6 decap_3
rlabel comment s 370436 200848 370436 200848 6 decap_3
rlabel comment s 370436 201936 370436 201936 6 decap_3
rlabel comment s 370436 203024 370436 203024 6 decap_3
rlabel comment s 370436 204112 370436 204112 6 decap_3
rlabel comment s 370436 205200 370436 205200 6 decap_3
rlabel comment s 370436 206288 370436 206288 6 decap_3
rlabel comment s 370436 207376 370436 207376 6 decap_3
rlabel comment s 370436 208464 370436 208464 6 decap_3
rlabel comment s 370436 209552 370436 209552 6 decap_3
rlabel comment s 370436 210640 370436 210640 6 decap_3
rlabel comment s 370436 211728 370436 211728 6 decap_3
rlabel comment s 370436 212816 370436 212816 6 decap_3
rlabel comment s 370436 213904 370436 213904 6 decap_3
rlabel comment s 370436 214992 370436 214992 6 decap_3
rlabel comment s 370436 216080 370436 216080 6 decap_3
rlabel comment s 370436 217168 370436 217168 6 decap_3
rlabel comment s 370436 218256 370436 218256 6 decap_3
rlabel comment s 370436 219344 370436 219344 6 decap_3
rlabel comment s 370436 220432 370436 220432 6 decap_3
rlabel comment s 370436 221520 370436 221520 6 decap_3
rlabel comment s 370436 222608 370436 222608 6 decap_3
rlabel comment s 370436 223696 370436 223696 6 decap_3
rlabel comment s 370436 224784 370436 224784 6 decap_3
rlabel comment s 370436 225872 370436 225872 6 decap_3
rlabel comment s 370436 226960 370436 226960 6 decap_3
rlabel comment s 370436 228048 370436 228048 6 decap_3
rlabel comment s 370436 229136 370436 229136 6 decap_3
rlabel comment s 370436 230224 370436 230224 6 decap_3
rlabel comment s 370436 231312 370436 231312 6 decap_3
rlabel comment s 370436 232400 370436 232400 6 decap_3
rlabel comment s 370436 233488 370436 233488 6 decap_3
rlabel comment s 370436 234576 370436 234576 6 decap_3
rlabel comment s 370436 235664 370436 235664 6 decap_3
rlabel comment s 370436 236752 370436 236752 6 decap_3
rlabel comment s 370436 237840 370436 237840 6 decap_3
rlabel comment s 370436 238928 370436 238928 6 decap_3
rlabel comment s 370436 240016 370436 240016 6 decap_3
rlabel comment s 370436 241104 370436 241104 6 decap_3
rlabel comment s 370436 242192 370436 242192 6 decap_3
rlabel comment s 370436 243280 370436 243280 6 decap_3
rlabel comment s 370436 244368 370436 244368 6 decap_3
rlabel comment s 370436 245456 370436 245456 6 decap_3
rlabel comment s 370436 246544 370436 246544 6 decap_3
rlabel comment s 370436 247632 370436 247632 6 decap_3
rlabel comment s 370436 253716 370436 253716 6 decap_3
rlabel comment s 370436 254804 370436 254804 6 decap_3
rlabel comment s 370436 255892 370436 255892 6 decap_3
rlabel comment s 370436 256980 370436 256980 6 decap_3
rlabel comment s 370436 258068 370436 258068 6 decap_3
rlabel comment s 370436 259156 370436 259156 6 decap_3
rlabel comment s 370436 260244 370436 260244 6 decap_3
rlabel comment s 370436 261332 370436 261332 6 decap_3
rlabel comment s 370436 262420 370436 262420 6 decap_3
rlabel comment s 370436 263508 370436 263508 6 decap_3
rlabel comment s 370436 264596 370436 264596 6 decap_3
rlabel comment s 370436 265684 370436 265684 6 decap_3
rlabel comment s 370436 266772 370436 266772 6 decap_3
rlabel comment s 370436 267860 370436 267860 6 decap_3
rlabel comment s 370436 268948 370436 268948 6 decap_3
rlabel comment s 370436 270036 370436 270036 6 decap_3
rlabel comment s 370436 271124 370436 271124 6 decap_3
rlabel comment s 370436 272212 370436 272212 6 decap_3
rlabel comment s 370436 273300 370436 273300 6 decap_3
rlabel comment s 370436 274388 370436 274388 6 decap_3
rlabel comment s 370436 275476 370436 275476 6 decap_3
rlabel comment s 370436 276564 370436 276564 6 decap_3
rlabel comment s 370436 277652 370436 277652 6 decap_3
rlabel comment s 370436 278740 370436 278740 6 decap_3
rlabel comment s 370436 279828 370436 279828 6 decap_3
rlabel comment s 370436 280916 370436 280916 6 decap_3
rlabel comment s 370436 282004 370436 282004 6 decap_3
rlabel comment s 370436 283092 370436 283092 6 decap_3
rlabel comment s 370436 284180 370436 284180 6 decap_3
rlabel comment s 370436 285268 370436 285268 6 decap_3
rlabel comment s 370436 286356 370436 286356 6 decap_3
rlabel comment s 370436 287444 370436 287444 6 decap_3
rlabel comment s 370436 288532 370436 288532 6 decap_3
rlabel comment s 370436 289620 370436 289620 6 decap_3
rlabel comment s 370436 290708 370436 290708 6 decap_3
rlabel comment s 370436 291796 370436 291796 6 decap_3
rlabel comment s 370436 292884 370436 292884 6 decap_3
rlabel comment s 370436 293972 370436 293972 6 decap_3
rlabel comment s 370436 295060 370436 295060 6 decap_3
rlabel comment s 370436 296148 370436 296148 6 decap_3
rlabel comment s 370436 297236 370436 297236 6 decap_3
rlabel comment s 370436 298324 370436 298324 6 decap_3
rlabel comment s 370436 299412 370436 299412 6 decap_3
rlabel comment s 370436 300500 370436 300500 6 decap_3
rlabel comment s 370436 301588 370436 301588 6 decap_3
rlabel comment s 370436 302676 370436 302676 6 decap_3
rlabel comment s 370436 303764 370436 303764 6 decap_3
rlabel comment s 370436 304852 370436 304852 6 decap_3
rlabel comment s 370436 305940 370436 305940 6 decap_3
rlabel comment s 370436 307028 370436 307028 6 decap_3
rlabel comment s 370436 308116 370436 308116 6 decap_3
rlabel comment s 370436 309204 370436 309204 6 decap_3
rlabel comment s 370436 310292 370436 310292 6 decap_3
rlabel comment s 370436 316376 370436 316376 6 decap_3
rlabel comment s 370436 317464 370436 317464 6 decap_3
rlabel comment s 370436 318552 370436 318552 6 decap_3
rlabel comment s 370436 319640 370436 319640 6 decap_3
rlabel comment s 370436 320728 370436 320728 6 decap_3
rlabel comment s 370436 321816 370436 321816 6 decap_3
rlabel comment s 370436 322904 370436 322904 6 decap_3
rlabel comment s 370436 323992 370436 323992 6 decap_3
rlabel comment s 370436 325080 370436 325080 6 decap_3
rlabel comment s 370436 326168 370436 326168 6 decap_3
rlabel comment s 370436 327256 370436 327256 6 decap_3
rlabel comment s 370436 328344 370436 328344 6 decap_3
rlabel comment s 370436 329432 370436 329432 6 decap_3
rlabel comment s 370436 330520 370436 330520 6 decap_3
rlabel comment s 370436 331608 370436 331608 6 decap_3
rlabel comment s 370436 332696 370436 332696 6 decap_3
rlabel comment s 370436 333784 370436 333784 6 decap_3
rlabel comment s 370436 334872 370436 334872 6 decap_3
rlabel comment s 370436 335960 370436 335960 6 decap_3
rlabel comment s 370436 337048 370436 337048 6 decap_3
rlabel comment s 370436 338136 370436 338136 6 decap_3
rlabel comment s 370436 339224 370436 339224 6 decap_3
rlabel comment s 370436 340312 370436 340312 6 decap_3
rlabel comment s 370436 341400 370436 341400 6 decap_3
rlabel comment s 370436 342488 370436 342488 6 decap_3
rlabel comment s 370436 343576 370436 343576 6 decap_3
rlabel comment s 370436 344664 370436 344664 6 decap_3
rlabel comment s 370436 345752 370436 345752 6 decap_3
rlabel comment s 370436 346840 370436 346840 6 decap_3
rlabel comment s 370436 347928 370436 347928 6 decap_3
rlabel comment s 370436 349016 370436 349016 6 decap_3
rlabel comment s 370436 350104 370436 350104 6 decap_3
rlabel comment s 370436 351192 370436 351192 6 decap_3
rlabel comment s 370436 352280 370436 352280 6 decap_3
rlabel comment s 370436 353368 370436 353368 6 decap_3
rlabel comment s 370436 354456 370436 354456 6 decap_3
rlabel comment s 370436 355544 370436 355544 6 decap_3
rlabel comment s 370436 356632 370436 356632 6 decap_3
rlabel comment s 370436 357720 370436 357720 6 decap_3
rlabel comment s 370436 358808 370436 358808 6 decap_3
rlabel comment s 370436 359896 370436 359896 6 decap_3
rlabel comment s 370436 360984 370436 360984 6 decap_3
rlabel comment s 370436 362072 370436 362072 6 decap_3
rlabel comment s 370436 363160 370436 363160 6 decap_3
rlabel comment s 370436 364248 370436 364248 6 decap_3
rlabel comment s 370436 365336 370436 365336 6 decap_3
rlabel comment s 370436 366424 370436 366424 6 decap_3
rlabel comment s 370436 367512 370436 367512 6 decap_3
rlabel comment s 370436 368600 370436 368600 6 decap_3
rlabel comment s 370436 369688 370436 369688 6 decap_3
rlabel comment s 370436 370776 370436 370776 6 decap_3
rlabel comment s 370436 371864 370436 371864 6 decap_3
rlabel comment s 370436 372952 370436 372952 6 decap_3
rlabel comment s 370436 379036 370436 379036 6 decap_3
rlabel comment s 370436 380124 370436 380124 6 decap_3
rlabel comment s 370436 381212 370436 381212 6 decap_3
rlabel comment s 370436 382300 370436 382300 6 decap_3
rlabel comment s 370436 383388 370436 383388 6 decap_3
rlabel comment s 370436 384476 370436 384476 6 decap_3
rlabel comment s 370436 385564 370436 385564 6 decap_3
rlabel comment s 370436 386652 370436 386652 6 decap_3
rlabel comment s 370436 387740 370436 387740 6 decap_3
rlabel comment s 370436 388828 370436 388828 6 decap_3
rlabel comment s 370436 389916 370436 389916 6 decap_3
rlabel comment s 370436 391004 370436 391004 6 decap_3
rlabel comment s 370436 392092 370436 392092 6 decap_3
rlabel comment s 370436 393180 370436 393180 6 decap_3
rlabel comment s 370436 394268 370436 394268 6 decap_3
rlabel comment s 370436 395356 370436 395356 6 decap_3
rlabel comment s 370436 396444 370436 396444 6 decap_3
rlabel comment s 370436 397532 370436 397532 6 decap_3
rlabel comment s 370436 398620 370436 398620 6 decap_3
rlabel comment s 370436 399708 370436 399708 6 decap_3
rlabel comment s 370436 400796 370436 400796 6 decap_3
rlabel comment s 370436 401884 370436 401884 6 decap_3
rlabel comment s 370436 402972 370436 402972 6 decap_3
rlabel comment s 370436 404060 370436 404060 6 decap_3
rlabel comment s 370436 405148 370436 405148 6 decap_3
rlabel comment s 370436 406236 370436 406236 6 decap_3
rlabel comment s 370436 407324 370436 407324 6 decap_3
rlabel comment s 370436 408412 370436 408412 6 decap_3
rlabel comment s 370436 409500 370436 409500 6 decap_3
rlabel comment s 370436 410588 370436 410588 6 decap_3
rlabel comment s 370436 411676 370436 411676 6 decap_3
rlabel comment s 370436 412764 370436 412764 6 decap_3
rlabel comment s 370436 413852 370436 413852 6 decap_3
rlabel comment s 370436 414940 370436 414940 6 decap_3
rlabel comment s 370436 416028 370436 416028 6 decap_3
rlabel comment s 370436 417116 370436 417116 6 decap_3
rlabel comment s 370436 418204 370436 418204 6 decap_3
rlabel comment s 370436 419292 370436 419292 6 decap_3
rlabel comment s 370436 420380 370436 420380 6 decap_3
rlabel comment s 370436 421468 370436 421468 6 decap_3
rlabel comment s 370436 422556 370436 422556 6 decap_3
rlabel comment s 370436 423644 370436 423644 6 decap_3
rlabel comment s 370436 424732 370436 424732 6 decap_3
rlabel comment s 370436 425820 370436 425820 6 decap_3
rlabel comment s 370436 426908 370436 426908 6 decap_3
rlabel comment s 370436 427996 370436 427996 6 decap_3
rlabel comment s 370436 429084 370436 429084 6 decap_3
rlabel comment s 370436 430172 370436 430172 6 decap_3
rlabel comment s 370436 431260 370436 431260 6 decap_3
rlabel comment s 370436 432348 370436 432348 6 decap_3
rlabel comment s 370436 433436 370436 433436 6 decap_3
rlabel comment s 370436 434524 370436 434524 6 decap_3
rlabel comment s 370436 435612 370436 435612 6 decap_3
rlabel comment s 370436 441696 370436 441696 6 decap_3
rlabel comment s 370436 442784 370436 442784 6 decap_3
rlabel comment s 370436 443872 370436 443872 6 decap_3
rlabel comment s 370436 444960 370436 444960 6 decap_3
rlabel comment s 370436 446048 370436 446048 6 decap_3
rlabel comment s 370436 447136 370436 447136 6 decap_3
rlabel comment s 370436 448224 370436 448224 6 decap_3
rlabel comment s 370436 449312 370436 449312 6 decap_3
rlabel comment s 370436 450400 370436 450400 6 decap_3
rlabel comment s 370436 451488 370436 451488 6 decap_3
rlabel comment s 370436 452576 370436 452576 6 decap_3
rlabel comment s 370436 453664 370436 453664 6 decap_3
rlabel comment s 370436 454752 370436 454752 6 decap_3
rlabel comment s 370436 455840 370436 455840 6 decap_3
rlabel comment s 370436 456928 370436 456928 6 decap_3
rlabel comment s 370436 458016 370436 458016 6 decap_3
rlabel comment s 370436 459104 370436 459104 6 decap_3
rlabel comment s 370436 460192 370436 460192 6 decap_3
rlabel comment s 370436 461280 370436 461280 6 decap_3
rlabel comment s 370436 462368 370436 462368 6 decap_3
rlabel comment s 370436 463456 370436 463456 6 decap_3
rlabel comment s 370436 464544 370436 464544 6 decap_3
rlabel comment s 370436 465632 370436 465632 6 decap_3
rlabel comment s 370436 466720 370436 466720 6 decap_3
rlabel comment s 370436 467808 370436 467808 6 decap_3
rlabel comment s 370436 468896 370436 468896 6 decap_3
rlabel comment s 370436 469984 370436 469984 6 decap_3
rlabel comment s 370436 471072 370436 471072 6 decap_3
rlabel comment s 370436 472160 370436 472160 6 decap_3
rlabel comment s 370436 473248 370436 473248 6 decap_3
rlabel comment s 370436 474336 370436 474336 6 decap_3
rlabel comment s 370436 475424 370436 475424 6 decap_3
rlabel comment s 370436 476512 370436 476512 6 decap_3
rlabel comment s 370436 477600 370436 477600 6 decap_3
rlabel comment s 370436 478688 370436 478688 6 decap_3
rlabel comment s 370436 479776 370436 479776 6 decap_3
rlabel comment s 370436 480864 370436 480864 6 decap_3
rlabel comment s 370436 481952 370436 481952 6 decap_3
rlabel comment s 370436 483040 370436 483040 6 decap_3
rlabel comment s 370436 484128 370436 484128 6 decap_3
rlabel comment s 370436 485216 370436 485216 6 decap_3
rlabel comment s 370436 486304 370436 486304 6 decap_3
rlabel comment s 370436 487392 370436 487392 6 decap_3
rlabel comment s 370436 488480 370436 488480 6 decap_3
rlabel comment s 370436 489568 370436 489568 6 decap_3
rlabel comment s 370436 490656 370436 490656 6 decap_3
rlabel comment s 370436 491744 370436 491744 6 decap_3
rlabel comment s 370436 492832 370436 492832 6 decap_3
rlabel comment s 370436 493920 370436 493920 6 decap_3
rlabel comment s 370436 495008 370436 495008 6 decap_3
rlabel comment s 370436 496096 370436 496096 6 decap_3
rlabel comment s 370436 497184 370436 497184 6 decap_3
rlabel comment s 370436 498272 370436 498272 6 decap_3
rlabel comment s 370436 504356 370436 504356 6 decap_3
rlabel comment s 370436 505444 370436 505444 6 decap_3
rlabel comment s 370436 506532 370436 506532 6 decap_3
rlabel comment s 370436 507620 370436 507620 6 decap_3
rlabel comment s 370436 508708 370436 508708 6 decap_3
rlabel comment s 370436 509796 370436 509796 6 decap_3
rlabel comment s 370436 510884 370436 510884 6 decap_3
rlabel comment s 370436 511972 370436 511972 6 decap_3
rlabel comment s 370436 513060 370436 513060 6 decap_3
rlabel comment s 370436 514148 370436 514148 6 decap_3
rlabel comment s 370436 515236 370436 515236 6 decap_3
rlabel comment s 370436 516324 370436 516324 6 decap_3
rlabel comment s 370436 517412 370436 517412 6 decap_3
rlabel comment s 370436 518500 370436 518500 6 decap_3
rlabel comment s 370436 519588 370436 519588 6 decap_3
rlabel comment s 370436 520676 370436 520676 6 decap_3
rlabel comment s 370436 521764 370436 521764 6 decap_3
rlabel comment s 370436 522852 370436 522852 6 decap_3
rlabel comment s 370436 523940 370436 523940 6 decap_3
rlabel comment s 370436 525028 370436 525028 6 decap_3
rlabel comment s 370436 526116 370436 526116 6 decap_3
rlabel comment s 370436 527204 370436 527204 6 decap_3
rlabel comment s 370436 528292 370436 528292 6 decap_3
rlabel comment s 370436 529380 370436 529380 6 decap_3
rlabel comment s 370436 530468 370436 530468 6 decap_3
rlabel comment s 370436 531556 370436 531556 6 decap_3
rlabel comment s 370436 532644 370436 532644 6 decap_3
rlabel comment s 370436 533732 370436 533732 6 decap_3
rlabel comment s 370436 534820 370436 534820 6 decap_3
rlabel comment s 370436 535908 370436 535908 6 decap_3
rlabel comment s 370436 536996 370436 536996 6 decap_3
rlabel comment s 370436 538084 370436 538084 6 decap_3
rlabel comment s 370436 539172 370436 539172 6 decap_3
rlabel comment s 370436 540260 370436 540260 6 decap_3
rlabel comment s 370436 541348 370436 541348 6 decap_3
rlabel comment s 370436 542436 370436 542436 6 decap_3
rlabel comment s 370436 543524 370436 543524 6 decap_3
rlabel comment s 370436 544612 370436 544612 6 decap_3
rlabel comment s 370436 545700 370436 545700 6 decap_3
rlabel comment s 370436 546788 370436 546788 6 decap_3
rlabel comment s 370436 547876 370436 547876 6 decap_3
rlabel comment s 370436 548964 370436 548964 6 decap_3
rlabel comment s 370436 550052 370436 550052 6 decap_3
rlabel comment s 370436 551140 370436 551140 6 decap_3
rlabel comment s 370436 552228 370436 552228 6 decap_3
rlabel comment s 370436 553316 370436 553316 6 decap_3
rlabel comment s 370436 554404 370436 554404 6 decap_3
rlabel comment s 370436 555492 370436 555492 6 decap_3
rlabel comment s 370436 556580 370436 556580 6 decap_3
rlabel comment s 370436 557668 370436 557668 6 decap_3
rlabel comment s 370436 558756 370436 558756 6 decap_3
rlabel comment s 370436 559844 370436 559844 6 decap_3
rlabel comment s 370436 560932 370436 560932 6 decap_3
rlabel comment s 495756 65736 495756 65736 6 decap_3
rlabel comment s 495756 66824 495756 66824 6 decap_3
rlabel comment s 495756 67912 495756 67912 6 decap_3
rlabel comment s 495756 69000 495756 69000 6 decap_3
rlabel comment s 495756 70088 495756 70088 6 decap_3
rlabel comment s 495756 71176 495756 71176 6 decap_3
rlabel comment s 495756 72264 495756 72264 6 decap_3
rlabel comment s 495756 73352 495756 73352 6 decap_3
rlabel comment s 495756 74440 495756 74440 6 decap_3
rlabel comment s 495756 75528 495756 75528 6 decap_3
rlabel comment s 495756 76616 495756 76616 6 decap_3
rlabel comment s 495756 77704 495756 77704 6 decap_3
rlabel comment s 495756 78792 495756 78792 6 decap_3
rlabel comment s 495756 79880 495756 79880 6 decap_3
rlabel comment s 495756 80968 495756 80968 6 decap_3
rlabel comment s 495756 82056 495756 82056 6 decap_3
rlabel comment s 495756 83144 495756 83144 6 decap_3
rlabel comment s 495756 84232 495756 84232 6 decap_3
rlabel comment s 495756 85320 495756 85320 6 decap_3
rlabel comment s 495756 86408 495756 86408 6 decap_3
rlabel comment s 495756 87496 495756 87496 6 decap_3
rlabel comment s 495756 88584 495756 88584 6 decap_3
rlabel comment s 495756 89672 495756 89672 6 decap_3
rlabel comment s 495756 90760 495756 90760 6 decap_3
rlabel comment s 495756 91848 495756 91848 6 decap_3
rlabel comment s 495756 92936 495756 92936 6 decap_3
rlabel comment s 495756 94024 495756 94024 6 decap_3
rlabel comment s 495756 95112 495756 95112 6 decap_3
rlabel comment s 495756 96200 495756 96200 6 decap_3
rlabel comment s 495756 97288 495756 97288 6 decap_3
rlabel comment s 495756 98376 495756 98376 6 decap_3
rlabel comment s 495756 99464 495756 99464 6 decap_3
rlabel comment s 495756 100552 495756 100552 6 decap_3
rlabel comment s 495756 101640 495756 101640 6 decap_3
rlabel comment s 495756 102728 495756 102728 6 decap_3
rlabel comment s 495756 103816 495756 103816 6 decap_3
rlabel comment s 495756 104904 495756 104904 6 decap_3
rlabel comment s 495756 105992 495756 105992 6 decap_3
rlabel comment s 495756 107080 495756 107080 6 decap_3
rlabel comment s 495756 108168 495756 108168 6 decap_3
rlabel comment s 495756 109256 495756 109256 6 decap_3
rlabel comment s 495756 110344 495756 110344 6 decap_3
rlabel comment s 495756 111432 495756 111432 6 decap_3
rlabel comment s 495756 112520 495756 112520 6 decap_3
rlabel comment s 495756 113608 495756 113608 6 decap_3
rlabel comment s 495756 114696 495756 114696 6 decap_3
rlabel comment s 495756 115784 495756 115784 6 decap_3
rlabel comment s 495756 116872 495756 116872 6 decap_3
rlabel comment s 495756 117960 495756 117960 6 decap_3
rlabel comment s 495756 119048 495756 119048 6 decap_3
rlabel comment s 495756 120136 495756 120136 6 decap_3
rlabel comment s 495756 121224 495756 121224 6 decap_3
rlabel comment s 495756 122312 495756 122312 6 decap_3
rlabel comment s 495756 128396 495756 128396 6 decap_3
rlabel comment s 495756 129484 495756 129484 6 decap_3
rlabel comment s 495756 130572 495756 130572 6 decap_3
rlabel comment s 495756 131660 495756 131660 6 decap_3
rlabel comment s 495756 132748 495756 132748 6 decap_3
rlabel comment s 495756 133836 495756 133836 6 decap_3
rlabel comment s 495756 134924 495756 134924 6 decap_3
rlabel comment s 495756 136012 495756 136012 6 decap_3
rlabel comment s 495756 137100 495756 137100 6 decap_3
rlabel comment s 495756 138188 495756 138188 6 decap_3
rlabel comment s 495756 139276 495756 139276 6 decap_3
rlabel comment s 495756 140364 495756 140364 6 decap_3
rlabel comment s 495756 141452 495756 141452 6 decap_3
rlabel comment s 495756 142540 495756 142540 6 decap_3
rlabel comment s 495756 143628 495756 143628 6 decap_3
rlabel comment s 495756 144716 495756 144716 6 decap_3
rlabel comment s 495756 145804 495756 145804 6 decap_3
rlabel comment s 495756 146892 495756 146892 6 decap_3
rlabel comment s 495756 147980 495756 147980 6 decap_3
rlabel comment s 495756 149068 495756 149068 6 decap_3
rlabel comment s 495756 150156 495756 150156 6 decap_3
rlabel comment s 495756 151244 495756 151244 6 decap_3
rlabel comment s 495756 152332 495756 152332 6 decap_3
rlabel comment s 495756 153420 495756 153420 6 decap_3
rlabel comment s 495756 154508 495756 154508 6 decap_3
rlabel comment s 495756 155596 495756 155596 6 decap_3
rlabel comment s 495756 156684 495756 156684 6 decap_3
rlabel comment s 495756 157772 495756 157772 6 decap_3
rlabel comment s 495756 158860 495756 158860 6 decap_3
rlabel comment s 495756 159948 495756 159948 6 decap_3
rlabel comment s 495756 161036 495756 161036 6 decap_3
rlabel comment s 495756 162124 495756 162124 6 decap_3
rlabel comment s 495756 163212 495756 163212 6 decap_3
rlabel comment s 495756 164300 495756 164300 6 decap_3
rlabel comment s 495756 165388 495756 165388 6 decap_3
rlabel comment s 495756 166476 495756 166476 6 decap_3
rlabel comment s 495756 167564 495756 167564 6 decap_3
rlabel comment s 495756 168652 495756 168652 6 decap_3
rlabel comment s 495756 169740 495756 169740 6 decap_3
rlabel comment s 495756 170828 495756 170828 6 decap_3
rlabel comment s 495756 171916 495756 171916 6 decap_3
rlabel comment s 495756 173004 495756 173004 6 decap_3
rlabel comment s 495756 174092 495756 174092 6 decap_3
rlabel comment s 495756 175180 495756 175180 6 decap_3
rlabel comment s 495756 176268 495756 176268 6 decap_3
rlabel comment s 495756 177356 495756 177356 6 decap_3
rlabel comment s 495756 178444 495756 178444 6 decap_3
rlabel comment s 495756 179532 495756 179532 6 decap_3
rlabel comment s 495756 180620 495756 180620 6 decap_3
rlabel comment s 495756 181708 495756 181708 6 decap_3
rlabel comment s 495756 182796 495756 182796 6 decap_3
rlabel comment s 495756 183884 495756 183884 6 decap_3
rlabel comment s 495756 184972 495756 184972 6 decap_3
rlabel comment s 495756 191056 495756 191056 6 decap_3
rlabel comment s 495756 192144 495756 192144 6 decap_3
rlabel comment s 495756 193232 495756 193232 6 decap_3
rlabel comment s 495756 194320 495756 194320 6 decap_3
rlabel comment s 495756 195408 495756 195408 6 decap_3
rlabel comment s 495756 196496 495756 196496 6 decap_3
rlabel comment s 495756 197584 495756 197584 6 decap_3
rlabel comment s 495756 198672 495756 198672 6 decap_3
rlabel comment s 495756 199760 495756 199760 6 decap_3
rlabel comment s 495756 200848 495756 200848 6 decap_3
rlabel comment s 495756 201936 495756 201936 6 decap_3
rlabel comment s 495756 203024 495756 203024 6 decap_3
rlabel comment s 495756 204112 495756 204112 6 decap_3
rlabel comment s 495756 205200 495756 205200 6 decap_3
rlabel comment s 495756 206288 495756 206288 6 decap_3
rlabel comment s 495756 207376 495756 207376 6 decap_3
rlabel comment s 495756 208464 495756 208464 6 decap_3
rlabel comment s 495756 209552 495756 209552 6 decap_3
rlabel comment s 495756 210640 495756 210640 6 decap_3
rlabel comment s 495756 211728 495756 211728 6 decap_3
rlabel comment s 495756 212816 495756 212816 6 decap_3
rlabel comment s 495756 213904 495756 213904 6 decap_3
rlabel comment s 495756 214992 495756 214992 6 decap_3
rlabel comment s 495756 216080 495756 216080 6 decap_3
rlabel comment s 495756 217168 495756 217168 6 decap_3
rlabel comment s 495756 218256 495756 218256 6 decap_3
rlabel comment s 495756 219344 495756 219344 6 decap_3
rlabel comment s 495756 220432 495756 220432 6 decap_3
rlabel comment s 495756 221520 495756 221520 6 decap_3
rlabel comment s 495756 222608 495756 222608 6 decap_3
rlabel comment s 495756 223696 495756 223696 6 decap_3
rlabel comment s 495756 224784 495756 224784 6 decap_3
rlabel comment s 495756 225872 495756 225872 6 decap_3
rlabel comment s 495756 226960 495756 226960 6 decap_3
rlabel comment s 495756 228048 495756 228048 6 decap_3
rlabel comment s 495756 229136 495756 229136 6 decap_3
rlabel comment s 495756 230224 495756 230224 6 decap_3
rlabel comment s 495756 231312 495756 231312 6 decap_3
rlabel comment s 495756 232400 495756 232400 6 decap_3
rlabel comment s 495756 233488 495756 233488 6 decap_3
rlabel comment s 495756 234576 495756 234576 6 decap_3
rlabel comment s 495756 235664 495756 235664 6 decap_3
rlabel comment s 495756 236752 495756 236752 6 decap_3
rlabel comment s 495756 237840 495756 237840 6 decap_3
rlabel comment s 495756 238928 495756 238928 6 decap_3
rlabel comment s 495756 240016 495756 240016 6 decap_3
rlabel comment s 495756 241104 495756 241104 6 decap_3
rlabel comment s 495756 242192 495756 242192 6 decap_3
rlabel comment s 495756 243280 495756 243280 6 decap_3
rlabel comment s 495756 244368 495756 244368 6 decap_3
rlabel comment s 495756 245456 495756 245456 6 decap_3
rlabel comment s 495756 246544 495756 246544 6 decap_3
rlabel comment s 495756 247632 495756 247632 6 decap_3
rlabel comment s 495756 253716 495756 253716 6 decap_3
rlabel comment s 495756 254804 495756 254804 6 decap_3
rlabel comment s 495756 255892 495756 255892 6 decap_3
rlabel comment s 495756 256980 495756 256980 6 decap_3
rlabel comment s 495756 258068 495756 258068 6 decap_3
rlabel comment s 495756 259156 495756 259156 6 decap_3
rlabel comment s 495756 260244 495756 260244 6 decap_3
rlabel comment s 495756 261332 495756 261332 6 decap_3
rlabel comment s 495756 262420 495756 262420 6 decap_3
rlabel comment s 495756 263508 495756 263508 6 decap_3
rlabel comment s 495756 264596 495756 264596 6 decap_3
rlabel comment s 495756 265684 495756 265684 6 decap_3
rlabel comment s 495756 266772 495756 266772 6 decap_3
rlabel comment s 495756 267860 495756 267860 6 decap_3
rlabel comment s 495756 268948 495756 268948 6 decap_3
rlabel comment s 495756 270036 495756 270036 6 decap_3
rlabel comment s 495756 271124 495756 271124 6 decap_3
rlabel comment s 495756 272212 495756 272212 6 decap_3
rlabel comment s 495756 273300 495756 273300 6 decap_3
rlabel comment s 495756 274388 495756 274388 6 decap_3
rlabel comment s 495756 275476 495756 275476 6 decap_3
rlabel comment s 495756 276564 495756 276564 6 decap_3
rlabel comment s 495756 277652 495756 277652 6 decap_3
rlabel comment s 495756 278740 495756 278740 6 decap_3
rlabel comment s 495756 279828 495756 279828 6 decap_3
rlabel comment s 495756 280916 495756 280916 6 decap_3
rlabel comment s 495756 282004 495756 282004 6 decap_3
rlabel comment s 495756 283092 495756 283092 6 decap_3
rlabel comment s 495756 284180 495756 284180 6 decap_3
rlabel comment s 495756 285268 495756 285268 6 decap_3
rlabel comment s 495756 286356 495756 286356 6 decap_3
rlabel comment s 495756 287444 495756 287444 6 decap_3
rlabel comment s 495756 288532 495756 288532 6 decap_3
rlabel comment s 495756 289620 495756 289620 6 decap_3
rlabel comment s 495756 290708 495756 290708 6 decap_3
rlabel comment s 495756 291796 495756 291796 6 decap_3
rlabel comment s 495756 292884 495756 292884 6 decap_3
rlabel comment s 495756 293972 495756 293972 6 decap_3
rlabel comment s 495756 295060 495756 295060 6 decap_3
rlabel comment s 495756 296148 495756 296148 6 decap_3
rlabel comment s 495756 297236 495756 297236 6 decap_3
rlabel comment s 495756 298324 495756 298324 6 decap_3
rlabel comment s 495756 299412 495756 299412 6 decap_3
rlabel comment s 495756 300500 495756 300500 6 decap_3
rlabel comment s 495756 301588 495756 301588 6 decap_3
rlabel comment s 495756 302676 495756 302676 6 decap_3
rlabel comment s 495756 303764 495756 303764 6 decap_3
rlabel comment s 495756 304852 495756 304852 6 decap_3
rlabel comment s 495756 305940 495756 305940 6 decap_3
rlabel comment s 495756 307028 495756 307028 6 decap_3
rlabel comment s 495756 308116 495756 308116 6 decap_3
rlabel comment s 495756 309204 495756 309204 6 decap_3
rlabel comment s 495756 310292 495756 310292 6 decap_3
rlabel comment s 495756 316376 495756 316376 6 decap_3
rlabel comment s 495756 317464 495756 317464 6 decap_3
rlabel comment s 495756 318552 495756 318552 6 decap_3
rlabel comment s 495756 319640 495756 319640 6 decap_3
rlabel comment s 495756 320728 495756 320728 6 decap_3
rlabel comment s 495756 321816 495756 321816 6 decap_3
rlabel comment s 495756 322904 495756 322904 6 decap_3
rlabel comment s 495756 323992 495756 323992 6 decap_3
rlabel comment s 495756 325080 495756 325080 6 decap_3
rlabel comment s 495756 326168 495756 326168 6 decap_3
rlabel comment s 495756 327256 495756 327256 6 decap_3
rlabel comment s 495756 328344 495756 328344 6 decap_3
rlabel comment s 495756 329432 495756 329432 6 decap_3
rlabel comment s 495756 330520 495756 330520 6 decap_3
rlabel comment s 495756 331608 495756 331608 6 decap_3
rlabel comment s 495756 332696 495756 332696 6 decap_3
rlabel comment s 495756 333784 495756 333784 6 decap_3
rlabel comment s 495756 334872 495756 334872 6 decap_3
rlabel comment s 495756 335960 495756 335960 6 decap_3
rlabel comment s 495756 337048 495756 337048 6 decap_3
rlabel comment s 495756 338136 495756 338136 6 decap_3
rlabel comment s 495756 339224 495756 339224 6 decap_3
rlabel comment s 495756 340312 495756 340312 6 decap_3
rlabel comment s 495756 341400 495756 341400 6 decap_3
rlabel comment s 495756 342488 495756 342488 6 decap_3
rlabel comment s 495756 343576 495756 343576 6 decap_3
rlabel comment s 495756 344664 495756 344664 6 decap_3
rlabel comment s 495756 345752 495756 345752 6 decap_3
rlabel comment s 495756 346840 495756 346840 6 decap_3
rlabel comment s 495756 347928 495756 347928 6 decap_3
rlabel comment s 495756 349016 495756 349016 6 decap_3
rlabel comment s 495756 350104 495756 350104 6 decap_3
rlabel comment s 495756 351192 495756 351192 6 decap_3
rlabel comment s 495756 352280 495756 352280 6 decap_3
rlabel comment s 495756 353368 495756 353368 6 decap_3
rlabel comment s 495756 354456 495756 354456 6 decap_3
rlabel comment s 495756 355544 495756 355544 6 decap_3
rlabel comment s 495756 356632 495756 356632 6 decap_3
rlabel comment s 495756 357720 495756 357720 6 decap_3
rlabel comment s 495756 358808 495756 358808 6 decap_3
rlabel comment s 495756 359896 495756 359896 6 decap_3
rlabel comment s 495756 360984 495756 360984 6 decap_3
rlabel comment s 495756 362072 495756 362072 6 decap_3
rlabel comment s 495756 363160 495756 363160 6 decap_3
rlabel comment s 495756 364248 495756 364248 6 decap_3
rlabel comment s 495756 365336 495756 365336 6 decap_3
rlabel comment s 495756 366424 495756 366424 6 decap_3
rlabel comment s 495756 367512 495756 367512 6 decap_3
rlabel comment s 495756 368600 495756 368600 6 decap_3
rlabel comment s 495756 369688 495756 369688 6 decap_3
rlabel comment s 495756 370776 495756 370776 6 decap_3
rlabel comment s 495756 371864 495756 371864 6 decap_3
rlabel comment s 495756 372952 495756 372952 6 decap_3
rlabel comment s 495756 379036 495756 379036 6 decap_3
rlabel comment s 495756 380124 495756 380124 6 decap_3
rlabel comment s 495756 381212 495756 381212 6 decap_3
rlabel comment s 495756 382300 495756 382300 6 decap_3
rlabel comment s 495756 383388 495756 383388 6 decap_3
rlabel comment s 495756 384476 495756 384476 6 decap_3
rlabel comment s 495756 385564 495756 385564 6 decap_3
rlabel comment s 495756 386652 495756 386652 6 decap_3
rlabel comment s 495756 387740 495756 387740 6 decap_3
rlabel comment s 495756 388828 495756 388828 6 decap_3
rlabel comment s 495756 389916 495756 389916 6 decap_3
rlabel comment s 495756 391004 495756 391004 6 decap_3
rlabel comment s 495756 392092 495756 392092 6 decap_3
rlabel comment s 495756 393180 495756 393180 6 decap_3
rlabel comment s 495756 394268 495756 394268 6 decap_3
rlabel comment s 495756 395356 495756 395356 6 decap_3
rlabel comment s 495756 396444 495756 396444 6 decap_3
rlabel comment s 495756 397532 495756 397532 6 decap_3
rlabel comment s 495756 398620 495756 398620 6 decap_3
rlabel comment s 495756 399708 495756 399708 6 decap_3
rlabel comment s 495756 400796 495756 400796 6 decap_3
rlabel comment s 495756 401884 495756 401884 6 decap_3
rlabel comment s 495756 402972 495756 402972 6 decap_3
rlabel comment s 495756 404060 495756 404060 6 decap_3
rlabel comment s 495756 405148 495756 405148 6 decap_3
rlabel comment s 495756 406236 495756 406236 6 decap_3
rlabel comment s 495756 407324 495756 407324 6 decap_3
rlabel comment s 495756 408412 495756 408412 6 decap_3
rlabel comment s 495756 409500 495756 409500 6 decap_3
rlabel comment s 495756 410588 495756 410588 6 decap_3
rlabel comment s 495756 411676 495756 411676 6 decap_3
rlabel comment s 495756 412764 495756 412764 6 decap_3
rlabel comment s 495756 413852 495756 413852 6 decap_3
rlabel comment s 495756 414940 495756 414940 6 decap_3
rlabel comment s 495756 416028 495756 416028 6 decap_3
rlabel comment s 495756 417116 495756 417116 6 decap_3
rlabel comment s 495756 418204 495756 418204 6 decap_3
rlabel comment s 495756 419292 495756 419292 6 decap_3
rlabel comment s 495756 420380 495756 420380 6 decap_3
rlabel comment s 495756 421468 495756 421468 6 decap_3
rlabel comment s 495756 422556 495756 422556 6 decap_3
rlabel comment s 495756 423644 495756 423644 6 decap_3
rlabel comment s 495756 424732 495756 424732 6 decap_3
rlabel comment s 495756 425820 495756 425820 6 decap_3
rlabel comment s 495756 426908 495756 426908 6 decap_3
rlabel comment s 495756 427996 495756 427996 6 decap_3
rlabel comment s 495756 429084 495756 429084 6 decap_3
rlabel comment s 495756 430172 495756 430172 6 decap_3
rlabel comment s 495756 431260 495756 431260 6 decap_3
rlabel comment s 495756 432348 495756 432348 6 decap_3
rlabel comment s 495756 433436 495756 433436 6 decap_3
rlabel comment s 495756 434524 495756 434524 6 decap_3
rlabel comment s 495756 435612 495756 435612 6 decap_3
rlabel comment s 495756 441696 495756 441696 6 decap_3
rlabel comment s 495756 442784 495756 442784 6 decap_3
rlabel comment s 495756 443872 495756 443872 6 decap_3
rlabel comment s 495756 444960 495756 444960 6 decap_3
rlabel comment s 495756 446048 495756 446048 6 decap_3
rlabel comment s 495756 447136 495756 447136 6 decap_3
rlabel comment s 495756 448224 495756 448224 6 decap_3
rlabel comment s 495756 449312 495756 449312 6 decap_3
rlabel comment s 495756 450400 495756 450400 6 decap_3
rlabel comment s 495756 451488 495756 451488 6 decap_3
rlabel comment s 495756 452576 495756 452576 6 decap_3
rlabel comment s 495756 453664 495756 453664 6 decap_3
rlabel comment s 495756 454752 495756 454752 6 decap_3
rlabel comment s 495756 455840 495756 455840 6 decap_3
rlabel comment s 495756 456928 495756 456928 6 decap_3
rlabel comment s 495756 458016 495756 458016 6 decap_3
rlabel comment s 495756 459104 495756 459104 6 decap_3
rlabel comment s 495756 460192 495756 460192 6 decap_3
rlabel comment s 495756 461280 495756 461280 6 decap_3
rlabel comment s 495756 462368 495756 462368 6 decap_3
rlabel comment s 495756 463456 495756 463456 6 decap_3
rlabel comment s 495756 464544 495756 464544 6 decap_3
rlabel comment s 495756 465632 495756 465632 6 decap_3
rlabel comment s 495756 466720 495756 466720 6 decap_3
rlabel comment s 495756 467808 495756 467808 6 decap_3
rlabel comment s 495756 468896 495756 468896 6 decap_3
rlabel comment s 495756 469984 495756 469984 6 decap_3
rlabel comment s 495756 471072 495756 471072 6 decap_3
rlabel comment s 495756 472160 495756 472160 6 decap_3
rlabel comment s 495756 473248 495756 473248 6 decap_3
rlabel comment s 495756 474336 495756 474336 6 decap_3
rlabel comment s 495756 475424 495756 475424 6 decap_3
rlabel comment s 495756 476512 495756 476512 6 decap_3
rlabel comment s 495756 477600 495756 477600 6 decap_3
rlabel comment s 495756 478688 495756 478688 6 decap_3
rlabel comment s 495756 479776 495756 479776 6 decap_3
rlabel comment s 495756 480864 495756 480864 6 decap_3
rlabel comment s 495756 481952 495756 481952 6 decap_3
rlabel comment s 495756 483040 495756 483040 6 decap_3
rlabel comment s 495756 484128 495756 484128 6 decap_3
rlabel comment s 495756 485216 495756 485216 6 decap_3
rlabel comment s 495756 486304 495756 486304 6 decap_3
rlabel comment s 495756 487392 495756 487392 6 decap_3
rlabel comment s 495756 488480 495756 488480 6 decap_3
rlabel comment s 495756 489568 495756 489568 6 decap_3
rlabel comment s 495756 490656 495756 490656 6 decap_3
rlabel comment s 495756 491744 495756 491744 6 decap_3
rlabel comment s 495756 492832 495756 492832 6 decap_3
rlabel comment s 495756 493920 495756 493920 6 decap_3
rlabel comment s 495756 495008 495756 495008 6 decap_3
rlabel comment s 495756 496096 495756 496096 6 decap_3
rlabel comment s 495756 497184 495756 497184 6 decap_3
rlabel comment s 495756 498272 495756 498272 6 decap_3
rlabel comment s 495756 504356 495756 504356 6 decap_3
rlabel comment s 495756 505444 495756 505444 6 decap_3
rlabel comment s 495756 506532 495756 506532 6 decap_3
rlabel comment s 495756 507620 495756 507620 6 decap_3
rlabel comment s 495756 508708 495756 508708 6 decap_3
rlabel comment s 495756 509796 495756 509796 6 decap_3
rlabel comment s 495756 510884 495756 510884 6 decap_3
rlabel comment s 495756 511972 495756 511972 6 decap_3
rlabel comment s 495756 513060 495756 513060 6 decap_3
rlabel comment s 495756 514148 495756 514148 6 decap_3
rlabel comment s 495756 515236 495756 515236 6 decap_3
rlabel comment s 495756 516324 495756 516324 6 decap_3
rlabel comment s 495756 517412 495756 517412 6 decap_3
rlabel comment s 495756 518500 495756 518500 6 decap_3
rlabel comment s 495756 519588 495756 519588 6 decap_3
rlabel comment s 495756 520676 495756 520676 6 decap_3
rlabel comment s 495756 521764 495756 521764 6 decap_3
rlabel comment s 495756 522852 495756 522852 6 decap_3
rlabel comment s 495756 523940 495756 523940 6 decap_3
rlabel comment s 495756 525028 495756 525028 6 decap_3
rlabel comment s 495756 526116 495756 526116 6 decap_3
rlabel comment s 495756 527204 495756 527204 6 decap_3
rlabel comment s 495756 528292 495756 528292 6 decap_3
rlabel comment s 495756 529380 495756 529380 6 decap_3
rlabel comment s 495756 530468 495756 530468 6 decap_3
rlabel comment s 495756 531556 495756 531556 6 decap_3
rlabel comment s 495756 532644 495756 532644 6 decap_3
rlabel comment s 495756 533732 495756 533732 6 decap_3
rlabel comment s 495756 534820 495756 534820 6 decap_3
rlabel comment s 495756 535908 495756 535908 6 decap_3
rlabel comment s 495756 536996 495756 536996 6 decap_3
rlabel comment s 495756 538084 495756 538084 6 decap_3
rlabel comment s 495756 539172 495756 539172 6 decap_3
rlabel comment s 495756 540260 495756 540260 6 decap_3
rlabel comment s 495756 541348 495756 541348 6 decap_3
rlabel comment s 495756 542436 495756 542436 6 decap_3
rlabel comment s 495756 543524 495756 543524 6 decap_3
rlabel comment s 495756 544612 495756 544612 6 decap_3
rlabel comment s 495756 545700 495756 545700 6 decap_3
rlabel comment s 495756 546788 495756 546788 6 decap_3
rlabel comment s 495756 547876 495756 547876 6 decap_3
rlabel comment s 495756 548964 495756 548964 6 decap_3
rlabel comment s 495756 550052 495756 550052 6 decap_3
rlabel comment s 495756 551140 495756 551140 6 decap_3
rlabel comment s 495756 552228 495756 552228 6 decap_3
rlabel comment s 495756 553316 495756 553316 6 decap_3
rlabel comment s 495756 554404 495756 554404 6 decap_3
rlabel comment s 495756 555492 495756 555492 6 decap_3
rlabel comment s 495756 556580 495756 556580 6 decap_3
rlabel comment s 495756 557668 495756 557668 6 decap_3
rlabel comment s 495756 558756 495756 558756 6 decap_3
rlabel comment s 495756 559844 495756 559844 6 decap_3
rlabel comment s 495756 560932 495756 560932 6 decap_3
rlabel comment s 502396 560488 502396 560488 2 decap_3
rlabel comment s 502396 559400 502396 559400 2 decap_3
rlabel comment s 502396 558312 502396 558312 2 decap_3
rlabel comment s 502396 557224 502396 557224 2 decap_3
rlabel comment s 502396 556136 502396 556136 2 decap_3
rlabel comment s 502396 555048 502396 555048 2 decap_3
rlabel comment s 502396 553960 502396 553960 2 decap_3
rlabel comment s 502396 552872 502396 552872 2 decap_3
rlabel comment s 502396 551784 502396 551784 2 decap_3
rlabel comment s 502396 550696 502396 550696 2 decap_3
rlabel comment s 502396 549608 502396 549608 2 decap_3
rlabel comment s 502396 548520 502396 548520 2 decap_3
rlabel comment s 502396 547432 502396 547432 2 decap_3
rlabel comment s 502396 546344 502396 546344 2 decap_3
rlabel comment s 502396 545256 502396 545256 2 decap_3
rlabel comment s 502396 544168 502396 544168 2 decap_3
rlabel comment s 502396 543080 502396 543080 2 decap_3
rlabel comment s 502396 541992 502396 541992 2 decap_3
rlabel comment s 502396 540904 502396 540904 2 decap_3
rlabel comment s 502396 539816 502396 539816 2 decap_3
rlabel comment s 502396 538728 502396 538728 2 decap_3
rlabel comment s 502396 537640 502396 537640 2 decap_3
rlabel comment s 502396 536552 502396 536552 2 decap_3
rlabel comment s 502396 535464 502396 535464 2 decap_3
rlabel comment s 502396 534376 502396 534376 2 decap_3
rlabel comment s 502396 533288 502396 533288 2 decap_3
rlabel comment s 502396 532200 502396 532200 2 decap_3
rlabel comment s 502396 531112 502396 531112 2 decap_3
rlabel comment s 502396 530024 502396 530024 2 decap_3
rlabel comment s 502396 528936 502396 528936 2 decap_3
rlabel comment s 502396 527848 502396 527848 2 decap_3
rlabel comment s 502396 526760 502396 526760 2 decap_3
rlabel comment s 502396 525672 502396 525672 2 decap_3
rlabel comment s 502396 524584 502396 524584 2 decap_3
rlabel comment s 502396 523496 502396 523496 2 decap_3
rlabel comment s 502396 522408 502396 522408 2 decap_3
rlabel comment s 502396 521320 502396 521320 2 decap_3
rlabel comment s 502396 520232 502396 520232 2 decap_3
rlabel comment s 502396 519144 502396 519144 2 decap_3
rlabel comment s 502396 518056 502396 518056 2 decap_3
rlabel comment s 502396 516968 502396 516968 2 decap_3
rlabel comment s 502396 515880 502396 515880 2 decap_3
rlabel comment s 502396 514792 502396 514792 2 decap_3
rlabel comment s 502396 513704 502396 513704 2 decap_3
rlabel comment s 502396 512616 502396 512616 2 decap_3
rlabel comment s 502396 511528 502396 511528 2 decap_3
rlabel comment s 502396 510440 502396 510440 2 decap_3
rlabel comment s 502396 509352 502396 509352 2 decap_3
rlabel comment s 502396 508264 502396 508264 2 decap_3
rlabel comment s 502396 507176 502396 507176 2 decap_3
rlabel comment s 502396 506088 502396 506088 2 decap_3
rlabel comment s 502396 505000 502396 505000 2 decap_3
rlabel comment s 502396 503912 502396 503912 2 decap_3
rlabel comment s 502396 497828 502396 497828 2 decap_3
rlabel comment s 502396 496740 502396 496740 2 decap_3
rlabel comment s 502396 495652 502396 495652 2 decap_3
rlabel comment s 502396 494564 502396 494564 2 decap_3
rlabel comment s 502396 493476 502396 493476 2 decap_3
rlabel comment s 502396 492388 502396 492388 2 decap_3
rlabel comment s 502396 491300 502396 491300 2 decap_3
rlabel comment s 502396 490212 502396 490212 2 decap_3
rlabel comment s 502396 489124 502396 489124 2 decap_3
rlabel comment s 502396 488036 502396 488036 2 decap_3
rlabel comment s 502396 486948 502396 486948 2 decap_3
rlabel comment s 502396 485860 502396 485860 2 decap_3
rlabel comment s 502396 484772 502396 484772 2 decap_3
rlabel comment s 502396 483684 502396 483684 2 decap_3
rlabel comment s 502396 482596 502396 482596 2 decap_3
rlabel comment s 502396 481508 502396 481508 2 decap_3
rlabel comment s 502396 480420 502396 480420 2 decap_3
rlabel comment s 502396 479332 502396 479332 2 decap_3
rlabel comment s 502396 478244 502396 478244 2 decap_3
rlabel comment s 502396 477156 502396 477156 2 decap_3
rlabel comment s 502396 476068 502396 476068 2 decap_3
rlabel comment s 502396 474980 502396 474980 2 decap_3
rlabel comment s 502396 473892 502396 473892 2 decap_3
rlabel comment s 502396 472804 502396 472804 2 decap_3
rlabel comment s 502396 471716 502396 471716 2 decap_3
rlabel comment s 502396 470628 502396 470628 2 decap_3
rlabel comment s 502396 469540 502396 469540 2 decap_3
rlabel comment s 502396 468452 502396 468452 2 decap_3
rlabel comment s 502396 467364 502396 467364 2 decap_3
rlabel comment s 502396 466276 502396 466276 2 decap_3
rlabel comment s 502396 465188 502396 465188 2 decap_3
rlabel comment s 502396 464100 502396 464100 2 decap_3
rlabel comment s 502396 463012 502396 463012 2 decap_3
rlabel comment s 502396 461924 502396 461924 2 decap_3
rlabel comment s 502396 460836 502396 460836 2 decap_3
rlabel comment s 502396 459748 502396 459748 2 decap_3
rlabel comment s 502396 458660 502396 458660 2 decap_3
rlabel comment s 502396 457572 502396 457572 2 decap_3
rlabel comment s 502396 456484 502396 456484 2 decap_3
rlabel comment s 502396 455396 502396 455396 2 decap_3
rlabel comment s 502396 454308 502396 454308 2 decap_3
rlabel comment s 502396 453220 502396 453220 2 decap_3
rlabel comment s 502396 452132 502396 452132 2 decap_3
rlabel comment s 502396 451044 502396 451044 2 decap_3
rlabel comment s 502396 449956 502396 449956 2 decap_3
rlabel comment s 502396 448868 502396 448868 2 decap_3
rlabel comment s 502396 447780 502396 447780 2 decap_3
rlabel comment s 502396 446692 502396 446692 2 decap_3
rlabel comment s 502396 445604 502396 445604 2 decap_3
rlabel comment s 502396 444516 502396 444516 2 decap_3
rlabel comment s 502396 443428 502396 443428 2 decap_3
rlabel comment s 502396 442340 502396 442340 2 decap_3
rlabel comment s 502396 441252 502396 441252 2 decap_3
rlabel comment s 502396 435168 502396 435168 2 decap_3
rlabel comment s 502396 434080 502396 434080 2 decap_3
rlabel comment s 502396 432992 502396 432992 2 decap_3
rlabel comment s 502396 431904 502396 431904 2 decap_3
rlabel comment s 502396 430816 502396 430816 2 decap_3
rlabel comment s 502396 429728 502396 429728 2 decap_3
rlabel comment s 502396 428640 502396 428640 2 decap_3
rlabel comment s 502396 427552 502396 427552 2 decap_3
rlabel comment s 502396 426464 502396 426464 2 decap_3
rlabel comment s 502396 425376 502396 425376 2 decap_3
rlabel comment s 502396 424288 502396 424288 2 decap_3
rlabel comment s 502396 423200 502396 423200 2 decap_3
rlabel comment s 502396 422112 502396 422112 2 decap_3
rlabel comment s 502396 421024 502396 421024 2 decap_3
rlabel comment s 502396 419936 502396 419936 2 decap_3
rlabel comment s 502396 418848 502396 418848 2 decap_3
rlabel comment s 502396 417760 502396 417760 2 decap_3
rlabel comment s 502396 416672 502396 416672 2 decap_3
rlabel comment s 502396 415584 502396 415584 2 decap_3
rlabel comment s 502396 414496 502396 414496 2 decap_3
rlabel comment s 502396 413408 502396 413408 2 decap_3
rlabel comment s 502396 412320 502396 412320 2 decap_3
rlabel comment s 502396 411232 502396 411232 2 decap_3
rlabel comment s 502396 410144 502396 410144 2 decap_3
rlabel comment s 502396 409056 502396 409056 2 decap_3
rlabel comment s 502396 407968 502396 407968 2 decap_3
rlabel comment s 502396 406880 502396 406880 2 decap_3
rlabel comment s 502396 405792 502396 405792 2 decap_3
rlabel comment s 502396 404704 502396 404704 2 decap_3
rlabel comment s 502396 403616 502396 403616 2 decap_3
rlabel comment s 502396 402528 502396 402528 2 decap_3
rlabel comment s 502396 401440 502396 401440 2 decap_3
rlabel comment s 502396 400352 502396 400352 2 decap_3
rlabel comment s 502396 399264 502396 399264 2 decap_3
rlabel comment s 502396 398176 502396 398176 2 decap_3
rlabel comment s 502396 397088 502396 397088 2 decap_3
rlabel comment s 502396 396000 502396 396000 2 decap_3
rlabel comment s 502396 394912 502396 394912 2 decap_3
rlabel comment s 502396 393824 502396 393824 2 decap_3
rlabel comment s 502396 392736 502396 392736 2 decap_3
rlabel comment s 502396 391648 502396 391648 2 decap_3
rlabel comment s 502396 390560 502396 390560 2 decap_3
rlabel comment s 502396 389472 502396 389472 2 decap_3
rlabel comment s 502396 388384 502396 388384 2 decap_3
rlabel comment s 502396 387296 502396 387296 2 decap_3
rlabel comment s 502396 386208 502396 386208 2 decap_3
rlabel comment s 502396 385120 502396 385120 2 decap_3
rlabel comment s 502396 384032 502396 384032 2 decap_3
rlabel comment s 502396 382944 502396 382944 2 decap_3
rlabel comment s 502396 381856 502396 381856 2 decap_3
rlabel comment s 502396 380768 502396 380768 2 decap_3
rlabel comment s 502396 379680 502396 379680 2 decap_3
rlabel comment s 502396 378592 502396 378592 2 decap_3
rlabel comment s 502396 372508 502396 372508 2 decap_3
rlabel comment s 502396 371420 502396 371420 2 decap_3
rlabel comment s 502396 370332 502396 370332 2 decap_3
rlabel comment s 502396 369244 502396 369244 2 decap_3
rlabel comment s 502396 368156 502396 368156 2 decap_3
rlabel comment s 502396 367068 502396 367068 2 decap_3
rlabel comment s 502396 365980 502396 365980 2 decap_3
rlabel comment s 502396 364892 502396 364892 2 decap_3
rlabel comment s 502396 363804 502396 363804 2 decap_3
rlabel comment s 502396 362716 502396 362716 2 decap_3
rlabel comment s 502396 361628 502396 361628 2 decap_3
rlabel comment s 502396 360540 502396 360540 2 decap_3
rlabel comment s 502396 359452 502396 359452 2 decap_3
rlabel comment s 502396 358364 502396 358364 2 decap_3
rlabel comment s 502396 357276 502396 357276 2 decap_3
rlabel comment s 502396 356188 502396 356188 2 decap_3
rlabel comment s 502396 355100 502396 355100 2 decap_3
rlabel comment s 502396 354012 502396 354012 2 decap_3
rlabel comment s 502396 352924 502396 352924 2 decap_3
rlabel comment s 502396 351836 502396 351836 2 decap_3
rlabel comment s 502396 350748 502396 350748 2 decap_3
rlabel comment s 502396 349660 502396 349660 2 decap_3
rlabel comment s 502396 348572 502396 348572 2 decap_3
rlabel comment s 502396 347484 502396 347484 2 decap_3
rlabel comment s 502396 346396 502396 346396 2 decap_3
rlabel comment s 502396 345308 502396 345308 2 decap_3
rlabel comment s 502396 344220 502396 344220 2 decap_3
rlabel comment s 502396 343132 502396 343132 2 decap_3
rlabel comment s 502396 342044 502396 342044 2 decap_3
rlabel comment s 502396 340956 502396 340956 2 decap_3
rlabel comment s 502396 339868 502396 339868 2 decap_3
rlabel comment s 502396 338780 502396 338780 2 decap_3
rlabel comment s 502396 337692 502396 337692 2 decap_3
rlabel comment s 502396 336604 502396 336604 2 decap_3
rlabel comment s 502396 335516 502396 335516 2 decap_3
rlabel comment s 502396 334428 502396 334428 2 decap_3
rlabel comment s 502396 333340 502396 333340 2 decap_3
rlabel comment s 502396 332252 502396 332252 2 decap_3
rlabel comment s 502396 331164 502396 331164 2 decap_3
rlabel comment s 502396 330076 502396 330076 2 decap_3
rlabel comment s 502396 328988 502396 328988 2 decap_3
rlabel comment s 502396 327900 502396 327900 2 decap_3
rlabel comment s 502396 326812 502396 326812 2 decap_3
rlabel comment s 502396 325724 502396 325724 2 decap_3
rlabel comment s 502396 324636 502396 324636 2 decap_3
rlabel comment s 502396 323548 502396 323548 2 decap_3
rlabel comment s 502396 322460 502396 322460 2 decap_3
rlabel comment s 502396 321372 502396 321372 2 decap_3
rlabel comment s 502396 320284 502396 320284 2 decap_3
rlabel comment s 502396 319196 502396 319196 2 decap_3
rlabel comment s 502396 318108 502396 318108 2 decap_3
rlabel comment s 502396 317020 502396 317020 2 decap_3
rlabel comment s 502396 315932 502396 315932 2 decap_3
rlabel comment s 502396 309848 502396 309848 2 decap_3
rlabel comment s 502396 308760 502396 308760 2 decap_3
rlabel comment s 502396 307672 502396 307672 2 decap_3
rlabel comment s 502396 306584 502396 306584 2 decap_3
rlabel comment s 502396 305496 502396 305496 2 decap_3
rlabel comment s 502396 304408 502396 304408 2 decap_3
rlabel comment s 502396 303320 502396 303320 2 decap_3
rlabel comment s 502396 302232 502396 302232 2 decap_3
rlabel comment s 502396 301144 502396 301144 2 decap_3
rlabel comment s 502396 300056 502396 300056 2 decap_3
rlabel comment s 502396 298968 502396 298968 2 decap_3
rlabel comment s 502396 297880 502396 297880 2 decap_3
rlabel comment s 502396 296792 502396 296792 2 decap_3
rlabel comment s 502396 295704 502396 295704 2 decap_3
rlabel comment s 502396 294616 502396 294616 2 decap_3
rlabel comment s 502396 293528 502396 293528 2 decap_3
rlabel comment s 502396 292440 502396 292440 2 decap_3
rlabel comment s 502396 291352 502396 291352 2 decap_3
rlabel comment s 502396 290264 502396 290264 2 decap_3
rlabel comment s 502396 289176 502396 289176 2 decap_3
rlabel comment s 502396 288088 502396 288088 2 decap_3
rlabel comment s 502396 287000 502396 287000 2 decap_3
rlabel comment s 502396 285912 502396 285912 2 decap_3
rlabel comment s 502396 284824 502396 284824 2 decap_3
rlabel comment s 502396 283736 502396 283736 2 decap_3
rlabel comment s 502396 282648 502396 282648 2 decap_3
rlabel comment s 502396 281560 502396 281560 2 decap_3
rlabel comment s 502396 280472 502396 280472 2 decap_3
rlabel comment s 502396 279384 502396 279384 2 decap_3
rlabel comment s 502396 278296 502396 278296 2 decap_3
rlabel comment s 502396 277208 502396 277208 2 decap_3
rlabel comment s 502396 276120 502396 276120 2 decap_3
rlabel comment s 502396 275032 502396 275032 2 decap_3
rlabel comment s 502396 273944 502396 273944 2 decap_3
rlabel comment s 502396 272856 502396 272856 2 decap_3
rlabel comment s 502396 271768 502396 271768 2 decap_3
rlabel comment s 502396 270680 502396 270680 2 decap_3
rlabel comment s 502396 269592 502396 269592 2 decap_3
rlabel comment s 502396 268504 502396 268504 2 decap_3
rlabel comment s 502396 267416 502396 267416 2 decap_3
rlabel comment s 502396 266328 502396 266328 2 decap_3
rlabel comment s 502396 265240 502396 265240 2 decap_3
rlabel comment s 502396 264152 502396 264152 2 decap_3
rlabel comment s 502396 263064 502396 263064 2 decap_3
rlabel comment s 502396 261976 502396 261976 2 decap_3
rlabel comment s 502396 260888 502396 260888 2 decap_3
rlabel comment s 502396 259800 502396 259800 2 decap_3
rlabel comment s 502396 258712 502396 258712 2 decap_3
rlabel comment s 502396 257624 502396 257624 2 decap_3
rlabel comment s 502396 256536 502396 256536 2 decap_3
rlabel comment s 502396 255448 502396 255448 2 decap_3
rlabel comment s 502396 254360 502396 254360 2 decap_3
rlabel comment s 502396 253272 502396 253272 2 decap_3
rlabel comment s 502396 247188 502396 247188 2 decap_3
rlabel comment s 502396 246100 502396 246100 2 decap_3
rlabel comment s 502396 245012 502396 245012 2 decap_3
rlabel comment s 502396 243924 502396 243924 2 decap_3
rlabel comment s 502396 242836 502396 242836 2 decap_3
rlabel comment s 502396 241748 502396 241748 2 decap_3
rlabel comment s 502396 240660 502396 240660 2 decap_3
rlabel comment s 502396 239572 502396 239572 2 decap_3
rlabel comment s 502396 238484 502396 238484 2 decap_3
rlabel comment s 502396 237396 502396 237396 2 decap_3
rlabel comment s 502396 236308 502396 236308 2 decap_3
rlabel comment s 502396 235220 502396 235220 2 decap_3
rlabel comment s 502396 234132 502396 234132 2 decap_3
rlabel comment s 502396 233044 502396 233044 2 decap_3
rlabel comment s 502396 231956 502396 231956 2 decap_3
rlabel comment s 502396 230868 502396 230868 2 decap_3
rlabel comment s 502396 229780 502396 229780 2 decap_3
rlabel comment s 502396 228692 502396 228692 2 decap_3
rlabel comment s 502396 227604 502396 227604 2 decap_3
rlabel comment s 502396 226516 502396 226516 2 decap_3
rlabel comment s 502396 225428 502396 225428 2 decap_3
rlabel comment s 502396 224340 502396 224340 2 decap_3
rlabel comment s 502396 223252 502396 223252 2 decap_3
rlabel comment s 502396 222164 502396 222164 2 decap_3
rlabel comment s 502396 221076 502396 221076 2 decap_3
rlabel comment s 502396 219988 502396 219988 2 decap_3
rlabel comment s 502396 218900 502396 218900 2 decap_3
rlabel comment s 502396 217812 502396 217812 2 decap_3
rlabel comment s 502396 216724 502396 216724 2 decap_3
rlabel comment s 502396 215636 502396 215636 2 decap_3
rlabel comment s 502396 214548 502396 214548 2 decap_3
rlabel comment s 502396 213460 502396 213460 2 decap_3
rlabel comment s 502396 212372 502396 212372 2 decap_3
rlabel comment s 502396 211284 502396 211284 2 decap_3
rlabel comment s 502396 210196 502396 210196 2 decap_3
rlabel comment s 502396 209108 502396 209108 2 decap_3
rlabel comment s 502396 208020 502396 208020 2 decap_3
rlabel comment s 502396 206932 502396 206932 2 decap_3
rlabel comment s 502396 205844 502396 205844 2 decap_3
rlabel comment s 502396 204756 502396 204756 2 decap_3
rlabel comment s 502396 203668 502396 203668 2 decap_3
rlabel comment s 502396 202580 502396 202580 2 decap_3
rlabel comment s 502396 201492 502396 201492 2 decap_3
rlabel comment s 502396 200404 502396 200404 2 decap_3
rlabel comment s 502396 199316 502396 199316 2 decap_3
rlabel comment s 502396 198228 502396 198228 2 decap_3
rlabel comment s 502396 197140 502396 197140 2 decap_3
rlabel comment s 502396 196052 502396 196052 2 decap_3
rlabel comment s 502396 194964 502396 194964 2 decap_3
rlabel comment s 502396 193876 502396 193876 2 decap_3
rlabel comment s 502396 192788 502396 192788 2 decap_3
rlabel comment s 502396 191700 502396 191700 2 decap_3
rlabel comment s 502396 190612 502396 190612 2 decap_3
rlabel comment s 502396 184528 502396 184528 2 decap_3
rlabel comment s 502396 183440 502396 183440 2 decap_3
rlabel comment s 502396 182352 502396 182352 2 decap_3
rlabel comment s 502396 181264 502396 181264 2 decap_3
rlabel comment s 502396 180176 502396 180176 2 decap_3
rlabel comment s 502396 179088 502396 179088 2 decap_3
rlabel comment s 502396 178000 502396 178000 2 decap_3
rlabel comment s 502396 176912 502396 176912 2 decap_3
rlabel comment s 502396 175824 502396 175824 2 decap_3
rlabel comment s 502396 174736 502396 174736 2 decap_3
rlabel comment s 502396 173648 502396 173648 2 decap_3
rlabel comment s 502396 172560 502396 172560 2 decap_3
rlabel comment s 502396 171472 502396 171472 2 decap_3
rlabel comment s 502396 170384 502396 170384 2 decap_3
rlabel comment s 502396 169296 502396 169296 2 decap_3
rlabel comment s 502396 168208 502396 168208 2 decap_3
rlabel comment s 502396 167120 502396 167120 2 decap_3
rlabel comment s 502396 166032 502396 166032 2 decap_3
rlabel comment s 502396 164944 502396 164944 2 decap_3
rlabel comment s 502396 163856 502396 163856 2 decap_3
rlabel comment s 502396 162768 502396 162768 2 decap_3
rlabel comment s 502396 161680 502396 161680 2 decap_3
rlabel comment s 502396 160592 502396 160592 2 decap_3
rlabel comment s 502396 159504 502396 159504 2 decap_3
rlabel comment s 502396 158416 502396 158416 2 decap_3
rlabel comment s 502396 157328 502396 157328 2 decap_3
rlabel comment s 502396 156240 502396 156240 2 decap_3
rlabel comment s 502396 155152 502396 155152 2 decap_3
rlabel comment s 502396 154064 502396 154064 2 decap_3
rlabel comment s 502396 152976 502396 152976 2 decap_3
rlabel comment s 502396 151888 502396 151888 2 decap_3
rlabel comment s 502396 150800 502396 150800 2 decap_3
rlabel comment s 502396 149712 502396 149712 2 decap_3
rlabel comment s 502396 148624 502396 148624 2 decap_3
rlabel comment s 502396 147536 502396 147536 2 decap_3
rlabel comment s 502396 146448 502396 146448 2 decap_3
rlabel comment s 502396 145360 502396 145360 2 decap_3
rlabel comment s 502396 144272 502396 144272 2 decap_3
rlabel comment s 502396 143184 502396 143184 2 decap_3
rlabel comment s 502396 142096 502396 142096 2 decap_3
rlabel comment s 502396 141008 502396 141008 2 decap_3
rlabel comment s 502396 139920 502396 139920 2 decap_3
rlabel comment s 502396 138832 502396 138832 2 decap_3
rlabel comment s 502396 137744 502396 137744 2 decap_3
rlabel comment s 502396 136656 502396 136656 2 decap_3
rlabel comment s 502396 135568 502396 135568 2 decap_3
rlabel comment s 502396 134480 502396 134480 2 decap_3
rlabel comment s 502396 133392 502396 133392 2 decap_3
rlabel comment s 502396 132304 502396 132304 2 decap_3
rlabel comment s 502396 131216 502396 131216 2 decap_3
rlabel comment s 502396 130128 502396 130128 2 decap_3
rlabel comment s 502396 129040 502396 129040 2 decap_3
rlabel comment s 502396 127952 502396 127952 2 decap_3
rlabel comment s 502396 121868 502396 121868 2 decap_3
rlabel comment s 502396 120780 502396 120780 2 decap_3
rlabel comment s 502396 119692 502396 119692 2 decap_3
rlabel comment s 502396 118604 502396 118604 2 decap_3
rlabel comment s 502396 117516 502396 117516 2 decap_3
rlabel comment s 502396 116428 502396 116428 2 decap_3
rlabel comment s 502396 115340 502396 115340 2 decap_3
rlabel comment s 502396 114252 502396 114252 2 decap_3
rlabel comment s 502396 113164 502396 113164 2 decap_3
rlabel comment s 502396 112076 502396 112076 2 decap_3
rlabel comment s 502396 110988 502396 110988 2 decap_3
rlabel comment s 502396 109900 502396 109900 2 decap_3
rlabel comment s 502396 108812 502396 108812 2 decap_3
rlabel comment s 502396 107724 502396 107724 2 decap_3
rlabel comment s 502396 106636 502396 106636 2 decap_3
rlabel comment s 502396 105548 502396 105548 2 decap_3
rlabel comment s 502396 104460 502396 104460 2 decap_3
rlabel comment s 502396 103372 502396 103372 2 decap_3
rlabel comment s 502396 102284 502396 102284 2 decap_3
rlabel comment s 502396 101196 502396 101196 2 decap_3
rlabel comment s 502396 100108 502396 100108 2 decap_3
rlabel comment s 502396 99020 502396 99020 2 decap_3
rlabel comment s 502396 97932 502396 97932 2 decap_3
rlabel comment s 502396 96844 502396 96844 2 decap_3
rlabel comment s 502396 95756 502396 95756 2 decap_3
rlabel comment s 502396 94668 502396 94668 2 decap_3
rlabel comment s 502396 93580 502396 93580 2 decap_3
rlabel comment s 502396 92492 502396 92492 2 decap_3
rlabel comment s 502396 91404 502396 91404 2 decap_3
rlabel comment s 502396 90316 502396 90316 2 decap_3
rlabel comment s 502396 89228 502396 89228 2 decap_3
rlabel comment s 502396 88140 502396 88140 2 decap_3
rlabel comment s 502396 87052 502396 87052 2 decap_3
rlabel comment s 502396 85964 502396 85964 2 decap_3
rlabel comment s 502396 84876 502396 84876 2 decap_3
rlabel comment s 502396 83788 502396 83788 2 decap_3
rlabel comment s 502396 82700 502396 82700 2 decap_3
rlabel comment s 502396 81612 502396 81612 2 decap_3
rlabel comment s 502396 80524 502396 80524 2 decap_3
rlabel comment s 502396 79436 502396 79436 2 decap_3
rlabel comment s 502396 78348 502396 78348 2 decap_3
rlabel comment s 502396 77260 502396 77260 2 decap_3
rlabel comment s 502396 76172 502396 76172 2 decap_3
rlabel comment s 502396 75084 502396 75084 2 decap_3
rlabel comment s 502396 73996 502396 73996 2 decap_3
rlabel comment s 502396 72908 502396 72908 2 decap_3
rlabel comment s 502396 71820 502396 71820 2 decap_3
rlabel comment s 502396 70732 502396 70732 2 decap_3
rlabel comment s 502396 69644 502396 69644 2 decap_3
rlabel comment s 502396 68556 502396 68556 2 decap_3
rlabel comment s 502396 67468 502396 67468 2 decap_3
rlabel comment s 502396 66380 502396 66380 2 decap_3
rlabel comment s 502396 65292 502396 65292 2 decap_3
rlabel comment s 377076 560488 377076 560488 2 decap_3
rlabel comment s 377076 559400 377076 559400 2 decap_3
rlabel comment s 377076 558312 377076 558312 2 decap_3
rlabel comment s 377076 557224 377076 557224 2 decap_3
rlabel comment s 377076 556136 377076 556136 2 decap_3
rlabel comment s 377076 555048 377076 555048 2 decap_3
rlabel comment s 377076 553960 377076 553960 2 decap_3
rlabel comment s 377076 552872 377076 552872 2 decap_3
rlabel comment s 377076 551784 377076 551784 2 decap_3
rlabel comment s 377076 550696 377076 550696 2 decap_3
rlabel comment s 377076 549608 377076 549608 2 decap_3
rlabel comment s 377076 548520 377076 548520 2 decap_3
rlabel comment s 377076 547432 377076 547432 2 decap_3
rlabel comment s 377076 546344 377076 546344 2 decap_3
rlabel comment s 377076 545256 377076 545256 2 decap_3
rlabel comment s 377076 544168 377076 544168 2 decap_3
rlabel comment s 377076 543080 377076 543080 2 decap_3
rlabel comment s 377076 541992 377076 541992 2 decap_3
rlabel comment s 377076 540904 377076 540904 2 decap_3
rlabel comment s 377076 539816 377076 539816 2 decap_3
rlabel comment s 377076 538728 377076 538728 2 decap_3
rlabel comment s 377076 537640 377076 537640 2 decap_3
rlabel comment s 377076 536552 377076 536552 2 decap_3
rlabel comment s 377076 535464 377076 535464 2 decap_3
rlabel comment s 377076 534376 377076 534376 2 decap_3
rlabel comment s 377076 533288 377076 533288 2 decap_3
rlabel comment s 377076 532200 377076 532200 2 decap_3
rlabel comment s 377076 531112 377076 531112 2 decap_3
rlabel comment s 377076 530024 377076 530024 2 decap_3
rlabel comment s 377076 528936 377076 528936 2 decap_3
rlabel comment s 377076 527848 377076 527848 2 decap_3
rlabel comment s 377076 526760 377076 526760 2 decap_3
rlabel comment s 377076 525672 377076 525672 2 decap_3
rlabel comment s 377076 524584 377076 524584 2 decap_3
rlabel comment s 377076 523496 377076 523496 2 decap_3
rlabel comment s 377076 522408 377076 522408 2 decap_3
rlabel comment s 377076 521320 377076 521320 2 decap_3
rlabel comment s 377076 520232 377076 520232 2 decap_3
rlabel comment s 377076 519144 377076 519144 2 decap_3
rlabel comment s 377076 518056 377076 518056 2 decap_3
rlabel comment s 377076 516968 377076 516968 2 decap_3
rlabel comment s 377076 515880 377076 515880 2 decap_3
rlabel comment s 377076 514792 377076 514792 2 decap_3
rlabel comment s 377076 513704 377076 513704 2 decap_3
rlabel comment s 377076 512616 377076 512616 2 decap_3
rlabel comment s 377076 511528 377076 511528 2 decap_3
rlabel comment s 377076 510440 377076 510440 2 decap_3
rlabel comment s 377076 509352 377076 509352 2 decap_3
rlabel comment s 377076 508264 377076 508264 2 decap_3
rlabel comment s 377076 507176 377076 507176 2 decap_3
rlabel comment s 377076 506088 377076 506088 2 decap_3
rlabel comment s 377076 505000 377076 505000 2 decap_3
rlabel comment s 377076 503912 377076 503912 2 decap_3
rlabel comment s 377076 497828 377076 497828 2 decap_3
rlabel comment s 377076 496740 377076 496740 2 decap_3
rlabel comment s 377076 495652 377076 495652 2 decap_3
rlabel comment s 377076 494564 377076 494564 2 decap_3
rlabel comment s 377076 493476 377076 493476 2 decap_3
rlabel comment s 377076 492388 377076 492388 2 decap_3
rlabel comment s 377076 491300 377076 491300 2 decap_3
rlabel comment s 377076 490212 377076 490212 2 decap_3
rlabel comment s 377076 489124 377076 489124 2 decap_3
rlabel comment s 377076 488036 377076 488036 2 decap_3
rlabel comment s 377076 486948 377076 486948 2 decap_3
rlabel comment s 377076 485860 377076 485860 2 decap_3
rlabel comment s 377076 484772 377076 484772 2 decap_3
rlabel comment s 377076 483684 377076 483684 2 decap_3
rlabel comment s 377076 482596 377076 482596 2 decap_3
rlabel comment s 377076 481508 377076 481508 2 decap_3
rlabel comment s 377076 480420 377076 480420 2 decap_3
rlabel comment s 377076 479332 377076 479332 2 decap_3
rlabel comment s 377076 478244 377076 478244 2 decap_3
rlabel comment s 377076 477156 377076 477156 2 decap_3
rlabel comment s 377076 476068 377076 476068 2 decap_3
rlabel comment s 377076 474980 377076 474980 2 decap_3
rlabel comment s 377076 473892 377076 473892 2 decap_3
rlabel comment s 377076 472804 377076 472804 2 decap_3
rlabel comment s 377076 471716 377076 471716 2 decap_3
rlabel comment s 377076 470628 377076 470628 2 decap_3
rlabel comment s 377076 469540 377076 469540 2 decap_3
rlabel comment s 377076 468452 377076 468452 2 decap_3
rlabel comment s 377076 467364 377076 467364 2 decap_3
rlabel comment s 377076 466276 377076 466276 2 decap_3
rlabel comment s 377076 465188 377076 465188 2 decap_3
rlabel comment s 377076 464100 377076 464100 2 decap_3
rlabel comment s 377076 463012 377076 463012 2 decap_3
rlabel comment s 377076 461924 377076 461924 2 decap_3
rlabel comment s 377076 460836 377076 460836 2 decap_3
rlabel comment s 377076 459748 377076 459748 2 decap_3
rlabel comment s 377076 458660 377076 458660 2 decap_3
rlabel comment s 377076 457572 377076 457572 2 decap_3
rlabel comment s 377076 456484 377076 456484 2 decap_3
rlabel comment s 377076 455396 377076 455396 2 decap_3
rlabel comment s 377076 454308 377076 454308 2 decap_3
rlabel comment s 377076 453220 377076 453220 2 decap_3
rlabel comment s 377076 452132 377076 452132 2 decap_3
rlabel comment s 377076 451044 377076 451044 2 decap_3
rlabel comment s 377076 449956 377076 449956 2 decap_3
rlabel comment s 377076 448868 377076 448868 2 decap_3
rlabel comment s 377076 447780 377076 447780 2 decap_3
rlabel comment s 377076 446692 377076 446692 2 decap_3
rlabel comment s 377076 445604 377076 445604 2 decap_3
rlabel comment s 377076 444516 377076 444516 2 decap_3
rlabel comment s 377076 443428 377076 443428 2 decap_3
rlabel comment s 377076 442340 377076 442340 2 decap_3
rlabel comment s 377076 441252 377076 441252 2 decap_3
rlabel comment s 377076 435168 377076 435168 2 decap_3
rlabel comment s 377076 434080 377076 434080 2 decap_3
rlabel comment s 377076 432992 377076 432992 2 decap_3
rlabel comment s 377076 431904 377076 431904 2 decap_3
rlabel comment s 377076 430816 377076 430816 2 decap_3
rlabel comment s 377076 429728 377076 429728 2 decap_3
rlabel comment s 377076 428640 377076 428640 2 decap_3
rlabel comment s 377076 427552 377076 427552 2 decap_3
rlabel comment s 377076 426464 377076 426464 2 decap_3
rlabel comment s 377076 425376 377076 425376 2 decap_3
rlabel comment s 377076 424288 377076 424288 2 decap_3
rlabel comment s 377076 423200 377076 423200 2 decap_3
rlabel comment s 377076 422112 377076 422112 2 decap_3
rlabel comment s 377076 421024 377076 421024 2 decap_3
rlabel comment s 377076 419936 377076 419936 2 decap_3
rlabel comment s 377076 418848 377076 418848 2 decap_3
rlabel comment s 377076 417760 377076 417760 2 decap_3
rlabel comment s 377076 416672 377076 416672 2 decap_3
rlabel comment s 377076 415584 377076 415584 2 decap_3
rlabel comment s 377076 414496 377076 414496 2 decap_3
rlabel comment s 377076 413408 377076 413408 2 decap_3
rlabel comment s 377076 412320 377076 412320 2 decap_3
rlabel comment s 377076 411232 377076 411232 2 decap_3
rlabel comment s 377076 410144 377076 410144 2 decap_3
rlabel comment s 377076 409056 377076 409056 2 decap_3
rlabel comment s 377076 407968 377076 407968 2 decap_3
rlabel comment s 377076 406880 377076 406880 2 decap_3
rlabel comment s 377076 405792 377076 405792 2 decap_3
rlabel comment s 377076 404704 377076 404704 2 decap_3
rlabel comment s 377076 403616 377076 403616 2 decap_3
rlabel comment s 377076 402528 377076 402528 2 decap_3
rlabel comment s 377076 401440 377076 401440 2 decap_3
rlabel comment s 377076 400352 377076 400352 2 decap_3
rlabel comment s 377076 399264 377076 399264 2 decap_3
rlabel comment s 377076 398176 377076 398176 2 decap_3
rlabel comment s 377076 397088 377076 397088 2 decap_3
rlabel comment s 377076 396000 377076 396000 2 decap_3
rlabel comment s 377076 394912 377076 394912 2 decap_3
rlabel comment s 377076 393824 377076 393824 2 decap_3
rlabel comment s 377076 392736 377076 392736 2 decap_3
rlabel comment s 377076 391648 377076 391648 2 decap_3
rlabel comment s 377076 390560 377076 390560 2 decap_3
rlabel comment s 377076 389472 377076 389472 2 decap_3
rlabel comment s 377076 388384 377076 388384 2 decap_3
rlabel comment s 377076 387296 377076 387296 2 decap_3
rlabel comment s 377076 386208 377076 386208 2 decap_3
rlabel comment s 377076 385120 377076 385120 2 decap_3
rlabel comment s 377076 384032 377076 384032 2 decap_3
rlabel comment s 377076 382944 377076 382944 2 decap_3
rlabel comment s 377076 381856 377076 381856 2 decap_3
rlabel comment s 377076 380768 377076 380768 2 decap_3
rlabel comment s 377076 379680 377076 379680 2 decap_3
rlabel comment s 377076 378592 377076 378592 2 decap_3
rlabel comment s 377076 372508 377076 372508 2 decap_3
rlabel comment s 377076 371420 377076 371420 2 decap_3
rlabel comment s 377076 370332 377076 370332 2 decap_3
rlabel comment s 377076 369244 377076 369244 2 decap_3
rlabel comment s 377076 368156 377076 368156 2 decap_3
rlabel comment s 377076 367068 377076 367068 2 decap_3
rlabel comment s 377076 365980 377076 365980 2 decap_3
rlabel comment s 377076 364892 377076 364892 2 decap_3
rlabel comment s 377076 363804 377076 363804 2 decap_3
rlabel comment s 377076 362716 377076 362716 2 decap_3
rlabel comment s 377076 361628 377076 361628 2 decap_3
rlabel comment s 377076 360540 377076 360540 2 decap_3
rlabel comment s 377076 359452 377076 359452 2 decap_3
rlabel comment s 377076 358364 377076 358364 2 decap_3
rlabel comment s 377076 357276 377076 357276 2 decap_3
rlabel comment s 377076 356188 377076 356188 2 decap_3
rlabel comment s 377076 355100 377076 355100 2 decap_3
rlabel comment s 377076 354012 377076 354012 2 decap_3
rlabel comment s 377076 352924 377076 352924 2 decap_3
rlabel comment s 377076 351836 377076 351836 2 decap_3
rlabel comment s 377076 350748 377076 350748 2 decap_3
rlabel comment s 377076 349660 377076 349660 2 decap_3
rlabel comment s 377076 348572 377076 348572 2 decap_3
rlabel comment s 377076 347484 377076 347484 2 decap_3
rlabel comment s 377076 346396 377076 346396 2 decap_3
rlabel comment s 377076 345308 377076 345308 2 decap_3
rlabel comment s 377076 344220 377076 344220 2 decap_3
rlabel comment s 377076 343132 377076 343132 2 decap_3
rlabel comment s 377076 342044 377076 342044 2 decap_3
rlabel comment s 377076 340956 377076 340956 2 decap_3
rlabel comment s 377076 339868 377076 339868 2 decap_3
rlabel comment s 377076 338780 377076 338780 2 decap_3
rlabel comment s 377076 337692 377076 337692 2 decap_3
rlabel comment s 377076 336604 377076 336604 2 decap_3
rlabel comment s 377076 335516 377076 335516 2 decap_3
rlabel comment s 377076 334428 377076 334428 2 decap_3
rlabel comment s 377076 333340 377076 333340 2 decap_3
rlabel comment s 377076 332252 377076 332252 2 decap_3
rlabel comment s 377076 331164 377076 331164 2 decap_3
rlabel comment s 377076 330076 377076 330076 2 decap_3
rlabel comment s 377076 328988 377076 328988 2 decap_3
rlabel comment s 377076 327900 377076 327900 2 decap_3
rlabel comment s 377076 326812 377076 326812 2 decap_3
rlabel comment s 377076 325724 377076 325724 2 decap_3
rlabel comment s 377076 324636 377076 324636 2 decap_3
rlabel comment s 377076 323548 377076 323548 2 decap_3
rlabel comment s 377076 322460 377076 322460 2 decap_3
rlabel comment s 377076 321372 377076 321372 2 decap_3
rlabel comment s 377076 320284 377076 320284 2 decap_3
rlabel comment s 377076 319196 377076 319196 2 decap_3
rlabel comment s 377076 318108 377076 318108 2 decap_3
rlabel comment s 377076 317020 377076 317020 2 decap_3
rlabel comment s 377076 315932 377076 315932 2 decap_3
rlabel comment s 377076 309848 377076 309848 2 decap_3
rlabel comment s 377076 308760 377076 308760 2 decap_3
rlabel comment s 377076 307672 377076 307672 2 decap_3
rlabel comment s 377076 306584 377076 306584 2 decap_3
rlabel comment s 377076 305496 377076 305496 2 decap_3
rlabel comment s 377076 304408 377076 304408 2 decap_3
rlabel comment s 377076 303320 377076 303320 2 decap_3
rlabel comment s 377076 302232 377076 302232 2 decap_3
rlabel comment s 377076 301144 377076 301144 2 decap_3
rlabel comment s 377076 300056 377076 300056 2 decap_3
rlabel comment s 377076 298968 377076 298968 2 decap_3
rlabel comment s 377076 297880 377076 297880 2 decap_3
rlabel comment s 377076 296792 377076 296792 2 decap_3
rlabel comment s 377076 295704 377076 295704 2 decap_3
rlabel comment s 377076 294616 377076 294616 2 decap_3
rlabel comment s 377076 293528 377076 293528 2 decap_3
rlabel comment s 377076 292440 377076 292440 2 decap_3
rlabel comment s 377076 291352 377076 291352 2 decap_3
rlabel comment s 377076 290264 377076 290264 2 decap_3
rlabel comment s 377076 289176 377076 289176 2 decap_3
rlabel comment s 377076 288088 377076 288088 2 decap_3
rlabel comment s 377076 287000 377076 287000 2 decap_3
rlabel comment s 377076 285912 377076 285912 2 decap_3
rlabel comment s 377076 284824 377076 284824 2 decap_3
rlabel comment s 377076 283736 377076 283736 2 decap_3
rlabel comment s 377076 282648 377076 282648 2 decap_3
rlabel comment s 377076 281560 377076 281560 2 decap_3
rlabel comment s 377076 280472 377076 280472 2 decap_3
rlabel comment s 377076 279384 377076 279384 2 decap_3
rlabel comment s 377076 278296 377076 278296 2 decap_3
rlabel comment s 377076 277208 377076 277208 2 decap_3
rlabel comment s 377076 276120 377076 276120 2 decap_3
rlabel comment s 377076 275032 377076 275032 2 decap_3
rlabel comment s 377076 273944 377076 273944 2 decap_3
rlabel comment s 377076 272856 377076 272856 2 decap_3
rlabel comment s 377076 271768 377076 271768 2 decap_3
rlabel comment s 377076 270680 377076 270680 2 decap_3
rlabel comment s 377076 269592 377076 269592 2 decap_3
rlabel comment s 377076 268504 377076 268504 2 decap_3
rlabel comment s 377076 267416 377076 267416 2 decap_3
rlabel comment s 377076 266328 377076 266328 2 decap_3
rlabel comment s 377076 265240 377076 265240 2 decap_3
rlabel comment s 377076 264152 377076 264152 2 decap_3
rlabel comment s 377076 263064 377076 263064 2 decap_3
rlabel comment s 377076 261976 377076 261976 2 decap_3
rlabel comment s 377076 260888 377076 260888 2 decap_3
rlabel comment s 377076 259800 377076 259800 2 decap_3
rlabel comment s 377076 258712 377076 258712 2 decap_3
rlabel comment s 377076 257624 377076 257624 2 decap_3
rlabel comment s 377076 256536 377076 256536 2 decap_3
rlabel comment s 377076 255448 377076 255448 2 decap_3
rlabel comment s 377076 254360 377076 254360 2 decap_3
rlabel comment s 377076 253272 377076 253272 2 decap_3
rlabel comment s 377076 247188 377076 247188 2 decap_3
rlabel comment s 377076 246100 377076 246100 2 decap_3
rlabel comment s 377076 245012 377076 245012 2 decap_3
rlabel comment s 377076 243924 377076 243924 2 decap_3
rlabel comment s 377076 242836 377076 242836 2 decap_3
rlabel comment s 377076 241748 377076 241748 2 decap_3
rlabel comment s 377076 240660 377076 240660 2 decap_3
rlabel comment s 377076 239572 377076 239572 2 decap_3
rlabel comment s 377076 238484 377076 238484 2 decap_3
rlabel comment s 377076 237396 377076 237396 2 decap_3
rlabel comment s 377076 236308 377076 236308 2 decap_3
rlabel comment s 377076 235220 377076 235220 2 decap_3
rlabel comment s 377076 234132 377076 234132 2 decap_3
rlabel comment s 377076 233044 377076 233044 2 decap_3
rlabel comment s 377076 231956 377076 231956 2 decap_3
rlabel comment s 377076 230868 377076 230868 2 decap_3
rlabel comment s 377076 229780 377076 229780 2 decap_3
rlabel comment s 377076 228692 377076 228692 2 decap_3
rlabel comment s 377076 227604 377076 227604 2 decap_3
rlabel comment s 377076 226516 377076 226516 2 decap_3
rlabel comment s 377076 225428 377076 225428 2 decap_3
rlabel comment s 377076 224340 377076 224340 2 decap_3
rlabel comment s 377076 223252 377076 223252 2 decap_3
rlabel comment s 377076 222164 377076 222164 2 decap_3
rlabel comment s 377076 221076 377076 221076 2 decap_3
rlabel comment s 377076 219988 377076 219988 2 decap_3
rlabel comment s 377076 218900 377076 218900 2 decap_3
rlabel comment s 377076 217812 377076 217812 2 decap_3
rlabel comment s 377076 216724 377076 216724 2 decap_3
rlabel comment s 377076 215636 377076 215636 2 decap_3
rlabel comment s 377076 214548 377076 214548 2 decap_3
rlabel comment s 377076 213460 377076 213460 2 decap_3
rlabel comment s 377076 212372 377076 212372 2 decap_3
rlabel comment s 377076 211284 377076 211284 2 decap_3
rlabel comment s 377076 210196 377076 210196 2 decap_3
rlabel comment s 377076 209108 377076 209108 2 decap_3
rlabel comment s 377076 208020 377076 208020 2 decap_3
rlabel comment s 377076 206932 377076 206932 2 decap_3
rlabel comment s 377076 205844 377076 205844 2 decap_3
rlabel comment s 377076 204756 377076 204756 2 decap_3
rlabel comment s 377076 203668 377076 203668 2 decap_3
rlabel comment s 377076 202580 377076 202580 2 decap_3
rlabel comment s 377076 201492 377076 201492 2 decap_3
rlabel comment s 377076 200404 377076 200404 2 decap_3
rlabel comment s 377076 199316 377076 199316 2 decap_3
rlabel comment s 377076 198228 377076 198228 2 decap_3
rlabel comment s 377076 197140 377076 197140 2 decap_3
rlabel comment s 377076 196052 377076 196052 2 decap_3
rlabel comment s 377076 194964 377076 194964 2 decap_3
rlabel comment s 377076 193876 377076 193876 2 decap_3
rlabel comment s 377076 192788 377076 192788 2 decap_3
rlabel comment s 377076 191700 377076 191700 2 decap_3
rlabel comment s 377076 190612 377076 190612 2 decap_3
rlabel comment s 377076 184528 377076 184528 2 decap_3
rlabel comment s 377076 183440 377076 183440 2 decap_3
rlabel comment s 377076 182352 377076 182352 2 decap_3
rlabel comment s 377076 181264 377076 181264 2 decap_3
rlabel comment s 377076 180176 377076 180176 2 decap_3
rlabel comment s 377076 179088 377076 179088 2 decap_3
rlabel comment s 377076 178000 377076 178000 2 decap_3
rlabel comment s 377076 176912 377076 176912 2 decap_3
rlabel comment s 377076 175824 377076 175824 2 decap_3
rlabel comment s 377076 174736 377076 174736 2 decap_3
rlabel comment s 377076 173648 377076 173648 2 decap_3
rlabel comment s 377076 172560 377076 172560 2 decap_3
rlabel comment s 377076 171472 377076 171472 2 decap_3
rlabel comment s 377076 170384 377076 170384 2 decap_3
rlabel comment s 377076 169296 377076 169296 2 decap_3
rlabel comment s 377076 168208 377076 168208 2 decap_3
rlabel comment s 377076 167120 377076 167120 2 decap_3
rlabel comment s 377076 166032 377076 166032 2 decap_3
rlabel comment s 377076 164944 377076 164944 2 decap_3
rlabel comment s 377076 163856 377076 163856 2 decap_3
rlabel comment s 377076 162768 377076 162768 2 decap_3
rlabel comment s 377076 161680 377076 161680 2 decap_3
rlabel comment s 377076 160592 377076 160592 2 decap_3
rlabel comment s 377076 159504 377076 159504 2 decap_3
rlabel comment s 377076 158416 377076 158416 2 decap_3
rlabel comment s 377076 157328 377076 157328 2 decap_3
rlabel comment s 377076 156240 377076 156240 2 decap_3
rlabel comment s 377076 155152 377076 155152 2 decap_3
rlabel comment s 377076 154064 377076 154064 2 decap_3
rlabel comment s 377076 152976 377076 152976 2 decap_3
rlabel comment s 377076 151888 377076 151888 2 decap_3
rlabel comment s 377076 150800 377076 150800 2 decap_3
rlabel comment s 377076 149712 377076 149712 2 decap_3
rlabel comment s 377076 148624 377076 148624 2 decap_3
rlabel comment s 377076 147536 377076 147536 2 decap_3
rlabel comment s 377076 146448 377076 146448 2 decap_3
rlabel comment s 377076 145360 377076 145360 2 decap_3
rlabel comment s 377076 144272 377076 144272 2 decap_3
rlabel comment s 377076 143184 377076 143184 2 decap_3
rlabel comment s 377076 142096 377076 142096 2 decap_3
rlabel comment s 377076 141008 377076 141008 2 decap_3
rlabel comment s 377076 139920 377076 139920 2 decap_3
rlabel comment s 377076 138832 377076 138832 2 decap_3
rlabel comment s 377076 137744 377076 137744 2 decap_3
rlabel comment s 377076 136656 377076 136656 2 decap_3
rlabel comment s 377076 135568 377076 135568 2 decap_3
rlabel comment s 377076 134480 377076 134480 2 decap_3
rlabel comment s 377076 133392 377076 133392 2 decap_3
rlabel comment s 377076 132304 377076 132304 2 decap_3
rlabel comment s 377076 131216 377076 131216 2 decap_3
rlabel comment s 377076 130128 377076 130128 2 decap_3
rlabel comment s 377076 129040 377076 129040 2 decap_3
rlabel comment s 377076 127952 377076 127952 2 decap_3
rlabel comment s 377076 121868 377076 121868 2 decap_3
rlabel comment s 377076 120780 377076 120780 2 decap_3
rlabel comment s 377076 119692 377076 119692 2 decap_3
rlabel comment s 377076 118604 377076 118604 2 decap_3
rlabel comment s 377076 117516 377076 117516 2 decap_3
rlabel comment s 377076 116428 377076 116428 2 decap_3
rlabel comment s 377076 115340 377076 115340 2 decap_3
rlabel comment s 377076 114252 377076 114252 2 decap_3
rlabel comment s 377076 113164 377076 113164 2 decap_3
rlabel comment s 377076 112076 377076 112076 2 decap_3
rlabel comment s 377076 110988 377076 110988 2 decap_3
rlabel comment s 377076 109900 377076 109900 2 decap_3
rlabel comment s 377076 108812 377076 108812 2 decap_3
rlabel comment s 377076 107724 377076 107724 2 decap_3
rlabel comment s 377076 106636 377076 106636 2 decap_3
rlabel comment s 377076 105548 377076 105548 2 decap_3
rlabel comment s 377076 104460 377076 104460 2 decap_3
rlabel comment s 377076 103372 377076 103372 2 decap_3
rlabel comment s 377076 102284 377076 102284 2 decap_3
rlabel comment s 377076 101196 377076 101196 2 decap_3
rlabel comment s 377076 100108 377076 100108 2 decap_3
rlabel comment s 377076 99020 377076 99020 2 decap_3
rlabel comment s 377076 97932 377076 97932 2 decap_3
rlabel comment s 377076 96844 377076 96844 2 decap_3
rlabel comment s 377076 95756 377076 95756 2 decap_3
rlabel comment s 377076 94668 377076 94668 2 decap_3
rlabel comment s 377076 93580 377076 93580 2 decap_3
rlabel comment s 377076 92492 377076 92492 2 decap_3
rlabel comment s 377076 91404 377076 91404 2 decap_3
rlabel comment s 377076 90316 377076 90316 2 decap_3
rlabel comment s 377076 89228 377076 89228 2 decap_3
rlabel comment s 377076 88140 377076 88140 2 decap_3
rlabel comment s 377076 87052 377076 87052 2 decap_3
rlabel comment s 377076 85964 377076 85964 2 decap_3
rlabel comment s 377076 84876 377076 84876 2 decap_3
rlabel comment s 377076 83788 377076 83788 2 decap_3
rlabel comment s 377076 82700 377076 82700 2 decap_3
rlabel comment s 377076 81612 377076 81612 2 decap_3
rlabel comment s 377076 80524 377076 80524 2 decap_3
rlabel comment s 377076 79436 377076 79436 2 decap_3
rlabel comment s 377076 78348 377076 78348 2 decap_3
rlabel comment s 377076 77260 377076 77260 2 decap_3
rlabel comment s 377076 76172 377076 76172 2 decap_3
rlabel comment s 377076 75084 377076 75084 2 decap_3
rlabel comment s 377076 73996 377076 73996 2 decap_3
rlabel comment s 377076 72908 377076 72908 2 decap_3
rlabel comment s 377076 71820 377076 71820 2 decap_3
rlabel comment s 377076 70732 377076 70732 2 decap_3
rlabel comment s 377076 69644 377076 69644 2 decap_3
rlabel comment s 377076 68556 377076 68556 2 decap_3
rlabel comment s 377076 67468 377076 67468 2 decap_3
rlabel comment s 377076 66380 377076 66380 2 decap_3
rlabel comment s 377076 65292 377076 65292 2 decap_3
rlabel metal1 119182 639676 119182 639676 5 SIgnal
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
