magic
tech sky130A
magscale 1 2
timestamp 1640660022
<< locali >>
rect 14013 10251 14047 13277
rect 14105 8959 14139 14229
rect 14013 3111 14047 6069
rect 14105 2635 14139 5593
<< viali >>
rect 1501 14569 1535 14603
rect 2145 14501 2179 14535
rect 4353 14501 4387 14535
rect 7113 14501 7147 14535
rect 12449 14501 12483 14535
rect 1593 14365 1627 14399
rect 7297 14365 7331 14399
rect 9873 14365 9907 14399
rect 13093 14365 13127 14399
rect 2329 14297 2363 14331
rect 4537 14297 4571 14331
rect 12265 14297 12299 14331
rect 9781 14229 9815 14263
rect 13001 14229 13035 14263
rect 14105 14229 14139 14263
rect 13001 13277 13035 13311
rect 14013 13277 14047 13311
rect 13185 13209 13219 13243
rect 1593 12121 1627 12155
rect 1501 12053 1535 12087
rect 5273 10761 5307 10795
rect 5641 10761 5675 10795
rect 7021 10761 7055 10795
rect 7389 10761 7423 10795
rect 8769 10761 8803 10795
rect 8953 10761 8987 10795
rect 5457 10693 5491 10727
rect 8677 10693 8711 10727
rect 5549 10625 5583 10659
rect 7113 10625 7147 10659
rect 7205 10625 7239 10659
rect 8585 10625 8619 10659
rect 5825 10489 5859 10523
rect 6837 10489 6871 10523
rect 8401 10489 8435 10523
rect 4997 10217 5031 10251
rect 6009 10217 6043 10251
rect 9505 10217 9539 10251
rect 14013 10217 14047 10251
rect 5181 10013 5215 10047
rect 6193 10013 6227 10047
rect 6377 10013 6411 10047
rect 9137 10013 9171 10047
rect 5273 9945 5307 9979
rect 5549 9945 5583 9979
rect 6561 9945 6595 9979
rect 8953 9945 8987 9979
rect 9321 9945 9355 9979
rect 5365 9877 5399 9911
rect 6285 9877 6319 9911
rect 9229 9877 9263 9911
rect 5365 9673 5399 9707
rect 4997 9605 5031 9639
rect 5273 9605 5307 9639
rect 5181 9537 5215 9571
rect 7481 9537 7515 9571
rect 8125 9537 8159 9571
rect 13001 9537 13035 9571
rect 5549 9401 5583 9435
rect 13185 9401 13219 9435
rect 7665 9333 7699 9367
rect 8309 9333 8343 9367
rect 10057 9129 10091 9163
rect 9505 9061 9539 9095
rect 7021 8925 7055 8959
rect 7849 8925 7883 8959
rect 9781 8925 9815 8959
rect 14105 8925 14139 8959
rect 7757 8857 7791 8891
rect 7113 8789 7147 8823
rect 9689 8789 9723 8823
rect 9873 8789 9907 8823
rect 5273 8585 5307 8619
rect 8401 8585 8435 8619
rect 5181 8517 5215 8551
rect 5365 8449 5399 8483
rect 6929 8449 6963 8483
rect 7573 8449 7607 8483
rect 8217 8449 8251 8483
rect 8861 8449 8895 8483
rect 5549 8313 5583 8347
rect 7113 8313 7147 8347
rect 7757 8313 7791 8347
rect 9045 8313 9079 8347
rect 4997 8245 5031 8279
rect 7849 8041 7883 8075
rect 7113 7905 7147 7939
rect 1593 7837 1627 7871
rect 7021 7837 7055 7871
rect 7941 7837 7975 7871
rect 1501 7701 1535 7735
rect 5457 7497 5491 7531
rect 7205 7497 7239 7531
rect 7941 7497 7975 7531
rect 9137 7497 9171 7531
rect 5641 7429 5675 7463
rect 8953 7429 8987 7463
rect 9321 7429 9355 7463
rect 5549 7361 5583 7395
rect 7021 7361 7055 7395
rect 7757 7361 7791 7395
rect 9229 7361 9263 7395
rect 5825 7225 5859 7259
rect 5273 7157 5307 7191
rect 9505 7157 9539 7191
rect 5273 6409 5307 6443
rect 6745 6409 6779 6443
rect 7757 6409 7791 6443
rect 9045 6409 9079 6443
rect 6561 6341 6595 6375
rect 7665 6341 7699 6375
rect 8953 6341 8987 6375
rect 5089 6273 5123 6307
rect 5181 6273 5215 6307
rect 5457 6273 5491 6307
rect 6653 6273 6687 6307
rect 7573 6273 7607 6307
rect 8861 6273 8895 6307
rect 6377 6205 6411 6239
rect 7389 6205 7423 6239
rect 8677 6205 8711 6239
rect 6929 6137 6963 6171
rect 4905 6069 4939 6103
rect 7941 6069 7975 6103
rect 9229 6069 9263 6103
rect 14013 6069 14047 6103
rect 8953 5797 8987 5831
rect 9229 5661 9263 5695
rect 13001 5661 13035 5695
rect 9321 5593 9355 5627
rect 9137 5525 9171 5559
rect 9505 5525 9539 5559
rect 13093 5525 13127 5559
rect 1593 4165 1627 4199
rect 1501 3893 1535 3927
rect 13001 3077 13035 3111
rect 14013 3077 14047 3111
rect 14105 5593 14139 5627
rect 13185 2873 13219 2907
rect 5641 2601 5675 2635
rect 13001 2601 13035 2635
rect 14105 2601 14139 2635
rect 1593 2397 1627 2431
rect 8217 2397 8251 2431
rect 11713 2397 11747 2431
rect 1409 2329 1443 2363
rect 2697 2329 2731 2363
rect 2881 2329 2915 2363
rect 5549 2329 5583 2363
rect 8033 2329 8067 2363
rect 11529 2329 11563 2363
rect 13093 2329 13127 2363
<< metal1 >>
rect 1104 14714 13892 14736
rect 1104 14662 3081 14714
rect 3133 14662 3145 14714
rect 3197 14662 3209 14714
rect 3261 14662 3273 14714
rect 3325 14662 3337 14714
rect 3389 14662 7344 14714
rect 7396 14662 7408 14714
rect 7460 14662 7472 14714
rect 7524 14662 7536 14714
rect 7588 14662 7600 14714
rect 7652 14662 11606 14714
rect 11658 14662 11670 14714
rect 11722 14662 11734 14714
rect 11786 14662 11798 14714
rect 11850 14662 11862 14714
rect 11914 14662 13892 14714
rect 1104 14640 13892 14662
rect 1486 14600 1492 14612
rect 1447 14572 1492 14600
rect 1486 14560 1492 14572
rect 1544 14560 1550 14612
rect 1670 14492 1676 14544
rect 1728 14532 1734 14544
rect 2133 14535 2191 14541
rect 2133 14532 2145 14535
rect 1728 14504 2145 14532
rect 1728 14492 1734 14504
rect 2133 14501 2145 14504
rect 2179 14501 2191 14535
rect 2133 14495 2191 14501
rect 4246 14492 4252 14544
rect 4304 14532 4310 14544
rect 4341 14535 4399 14541
rect 4341 14532 4353 14535
rect 4304 14504 4353 14532
rect 4304 14492 4310 14504
rect 4341 14501 4353 14504
rect 4387 14501 4399 14535
rect 4341 14495 4399 14501
rect 7006 14492 7012 14544
rect 7064 14532 7070 14544
rect 7101 14535 7159 14541
rect 7101 14532 7113 14535
rect 7064 14504 7113 14532
rect 7064 14492 7070 14504
rect 7101 14501 7113 14504
rect 7147 14501 7159 14535
rect 7101 14495 7159 14501
rect 12342 14492 12348 14544
rect 12400 14532 12406 14544
rect 12437 14535 12495 14541
rect 12437 14532 12449 14535
rect 12400 14504 12449 14532
rect 12400 14492 12406 14504
rect 12437 14501 12449 14504
rect 12483 14501 12495 14535
rect 12437 14495 12495 14501
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14396 1639 14399
rect 3786 14396 3792 14408
rect 1627 14368 3792 14396
rect 1627 14365 1639 14368
rect 1581 14359 1639 14365
rect 3786 14356 3792 14368
rect 3844 14356 3850 14408
rect 7190 14356 7196 14408
rect 7248 14396 7254 14408
rect 7285 14399 7343 14405
rect 7285 14396 7297 14399
rect 7248 14368 7297 14396
rect 7248 14356 7254 14368
rect 7285 14365 7297 14368
rect 7331 14365 7343 14399
rect 7285 14359 7343 14365
rect 9674 14356 9680 14408
rect 9732 14396 9738 14408
rect 9861 14399 9919 14405
rect 9861 14396 9873 14399
rect 9732 14368 9873 14396
rect 9732 14356 9738 14368
rect 9861 14365 9873 14368
rect 9907 14365 9919 14399
rect 9861 14359 9919 14365
rect 13081 14399 13139 14405
rect 13081 14365 13093 14399
rect 13127 14396 13139 14399
rect 14918 14396 14924 14408
rect 13127 14368 14924 14396
rect 13127 14365 13139 14368
rect 13081 14359 13139 14365
rect 14918 14356 14924 14368
rect 14976 14356 14982 14408
rect 2317 14331 2375 14337
rect 2317 14297 2329 14331
rect 2363 14328 2375 14331
rect 4062 14328 4068 14340
rect 2363 14300 4068 14328
rect 2363 14297 2375 14300
rect 2317 14291 2375 14297
rect 4062 14288 4068 14300
rect 4120 14288 4126 14340
rect 4525 14331 4583 14337
rect 4525 14297 4537 14331
rect 4571 14328 4583 14331
rect 5994 14328 6000 14340
rect 4571 14300 6000 14328
rect 4571 14297 4583 14300
rect 4525 14291 4583 14297
rect 5994 14288 6000 14300
rect 6052 14288 6058 14340
rect 12250 14328 12256 14340
rect 12211 14300 12256 14328
rect 12250 14288 12256 14300
rect 12308 14288 12314 14340
rect 9769 14263 9827 14269
rect 9769 14229 9781 14263
rect 9815 14260 9827 14263
rect 9858 14260 9864 14272
rect 9815 14232 9864 14260
rect 9815 14229 9827 14232
rect 9769 14223 9827 14229
rect 9858 14220 9864 14232
rect 9916 14220 9922 14272
rect 12989 14263 13047 14269
rect 12989 14229 13001 14263
rect 13035 14260 13047 14263
rect 14093 14263 14151 14269
rect 14093 14260 14105 14263
rect 13035 14232 14105 14260
rect 13035 14229 13047 14232
rect 12989 14223 13047 14229
rect 14093 14229 14105 14232
rect 14139 14229 14151 14263
rect 14093 14223 14151 14229
rect 1104 14170 13892 14192
rect 1104 14118 5212 14170
rect 5264 14118 5276 14170
rect 5328 14118 5340 14170
rect 5392 14118 5404 14170
rect 5456 14118 5468 14170
rect 5520 14118 9475 14170
rect 9527 14118 9539 14170
rect 9591 14118 9603 14170
rect 9655 14118 9667 14170
rect 9719 14118 9731 14170
rect 9783 14118 13892 14170
rect 1104 14096 13892 14118
rect 1104 13626 13892 13648
rect 1104 13574 3081 13626
rect 3133 13574 3145 13626
rect 3197 13574 3209 13626
rect 3261 13574 3273 13626
rect 3325 13574 3337 13626
rect 3389 13574 7344 13626
rect 7396 13574 7408 13626
rect 7460 13574 7472 13626
rect 7524 13574 7536 13626
rect 7588 13574 7600 13626
rect 7652 13574 11606 13626
rect 11658 13574 11670 13626
rect 11722 13574 11734 13626
rect 11786 13574 11798 13626
rect 11850 13574 11862 13626
rect 11914 13574 13892 13626
rect 1104 13552 13892 13574
rect 12989 13311 13047 13317
rect 12989 13277 13001 13311
rect 13035 13308 13047 13311
rect 14001 13311 14059 13317
rect 14001 13308 14013 13311
rect 13035 13280 14013 13308
rect 13035 13277 13047 13280
rect 12989 13271 13047 13277
rect 14001 13277 14013 13280
rect 14047 13277 14059 13311
rect 14001 13271 14059 13277
rect 13170 13240 13176 13252
rect 13131 13212 13176 13240
rect 13170 13200 13176 13212
rect 13228 13200 13234 13252
rect 1104 13082 13892 13104
rect 1104 13030 5212 13082
rect 5264 13030 5276 13082
rect 5328 13030 5340 13082
rect 5392 13030 5404 13082
rect 5456 13030 5468 13082
rect 5520 13030 9475 13082
rect 9527 13030 9539 13082
rect 9591 13030 9603 13082
rect 9655 13030 9667 13082
rect 9719 13030 9731 13082
rect 9783 13030 13892 13082
rect 1104 13008 13892 13030
rect 1104 12538 13892 12560
rect 1104 12486 3081 12538
rect 3133 12486 3145 12538
rect 3197 12486 3209 12538
rect 3261 12486 3273 12538
rect 3325 12486 3337 12538
rect 3389 12486 7344 12538
rect 7396 12486 7408 12538
rect 7460 12486 7472 12538
rect 7524 12486 7536 12538
rect 7588 12486 7600 12538
rect 7652 12486 11606 12538
rect 11658 12486 11670 12538
rect 11722 12486 11734 12538
rect 11786 12486 11798 12538
rect 11850 12486 11862 12538
rect 11914 12486 13892 12538
rect 1104 12464 13892 12486
rect 1581 12155 1639 12161
rect 1581 12121 1593 12155
rect 1627 12152 1639 12155
rect 4982 12152 4988 12164
rect 1627 12124 4988 12152
rect 1627 12121 1639 12124
rect 1581 12115 1639 12121
rect 4982 12112 4988 12124
rect 5040 12112 5046 12164
rect 1486 12084 1492 12096
rect 1447 12056 1492 12084
rect 1486 12044 1492 12056
rect 1544 12044 1550 12096
rect 1104 11994 13892 12016
rect 1104 11942 5212 11994
rect 5264 11942 5276 11994
rect 5328 11942 5340 11994
rect 5392 11942 5404 11994
rect 5456 11942 5468 11994
rect 5520 11942 9475 11994
rect 9527 11942 9539 11994
rect 9591 11942 9603 11994
rect 9655 11942 9667 11994
rect 9719 11942 9731 11994
rect 9783 11942 13892 11994
rect 1104 11920 13892 11942
rect 1104 11450 13892 11472
rect 1104 11398 3081 11450
rect 3133 11398 3145 11450
rect 3197 11398 3209 11450
rect 3261 11398 3273 11450
rect 3325 11398 3337 11450
rect 3389 11398 7344 11450
rect 7396 11398 7408 11450
rect 7460 11398 7472 11450
rect 7524 11398 7536 11450
rect 7588 11398 7600 11450
rect 7652 11398 11606 11450
rect 11658 11398 11670 11450
rect 11722 11398 11734 11450
rect 11786 11398 11798 11450
rect 11850 11398 11862 11450
rect 11914 11398 13892 11450
rect 1104 11376 13892 11398
rect 1104 10906 13892 10928
rect 1104 10854 5212 10906
rect 5264 10854 5276 10906
rect 5328 10854 5340 10906
rect 5392 10854 5404 10906
rect 5456 10854 5468 10906
rect 5520 10854 9475 10906
rect 9527 10854 9539 10906
rect 9591 10854 9603 10906
rect 9655 10854 9667 10906
rect 9719 10854 9731 10906
rect 9783 10854 13892 10906
rect 1104 10832 13892 10854
rect 4062 10752 4068 10804
rect 4120 10792 4126 10804
rect 5261 10795 5319 10801
rect 5261 10792 5273 10795
rect 4120 10764 5273 10792
rect 4120 10752 4126 10764
rect 5261 10761 5273 10764
rect 5307 10761 5319 10795
rect 5261 10755 5319 10761
rect 5629 10795 5687 10801
rect 5629 10761 5641 10795
rect 5675 10792 5687 10795
rect 6914 10792 6920 10804
rect 5675 10764 6920 10792
rect 5675 10761 5687 10764
rect 5629 10755 5687 10761
rect 6914 10752 6920 10764
rect 6972 10752 6978 10804
rect 7006 10752 7012 10804
rect 7064 10792 7070 10804
rect 7064 10764 7109 10792
rect 7064 10752 7070 10764
rect 7190 10752 7196 10804
rect 7248 10792 7254 10804
rect 7377 10795 7435 10801
rect 7377 10792 7389 10795
rect 7248 10764 7389 10792
rect 7248 10752 7254 10764
rect 7377 10761 7389 10764
rect 7423 10761 7435 10795
rect 8757 10795 8815 10801
rect 8757 10792 8769 10795
rect 7377 10755 7435 10761
rect 7760 10764 8769 10792
rect 5445 10727 5503 10733
rect 5445 10693 5457 10727
rect 5491 10724 5503 10727
rect 5491 10696 5672 10724
rect 5491 10693 5503 10696
rect 5445 10687 5503 10693
rect 5644 10668 5672 10696
rect 7760 10668 7788 10764
rect 8757 10761 8769 10764
rect 8803 10761 8815 10795
rect 8757 10755 8815 10761
rect 8941 10795 8999 10801
rect 8941 10761 8953 10795
rect 8987 10792 8999 10795
rect 12250 10792 12256 10804
rect 8987 10764 12256 10792
rect 8987 10761 8999 10764
rect 8941 10755 8999 10761
rect 12250 10752 12256 10764
rect 12308 10752 12314 10804
rect 8202 10684 8208 10736
rect 8260 10724 8266 10736
rect 8665 10727 8723 10733
rect 8665 10724 8677 10727
rect 8260 10696 8677 10724
rect 8260 10684 8266 10696
rect 8665 10693 8677 10696
rect 8711 10693 8723 10727
rect 8665 10687 8723 10693
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10625 5595 10659
rect 5537 10619 5595 10625
rect 5258 10548 5264 10600
rect 5316 10588 5322 10600
rect 5552 10588 5580 10619
rect 5626 10616 5632 10668
rect 5684 10616 5690 10668
rect 7101 10659 7159 10665
rect 7101 10625 7113 10659
rect 7147 10625 7159 10659
rect 7101 10619 7159 10625
rect 7193 10659 7251 10665
rect 7193 10625 7205 10659
rect 7239 10656 7251 10659
rect 7742 10656 7748 10668
rect 7239 10628 7748 10656
rect 7239 10625 7251 10628
rect 7193 10619 7251 10625
rect 7116 10588 7144 10619
rect 7742 10616 7748 10628
rect 7800 10616 7806 10668
rect 8110 10616 8116 10668
rect 8168 10656 8174 10668
rect 8573 10659 8631 10665
rect 8573 10656 8585 10659
rect 8168 10628 8585 10656
rect 8168 10616 8174 10628
rect 8573 10625 8585 10628
rect 8619 10625 8631 10659
rect 8573 10619 8631 10625
rect 7926 10588 7932 10600
rect 5316 10560 7932 10588
rect 5316 10548 5322 10560
rect 7926 10548 7932 10560
rect 7984 10548 7990 10600
rect 5813 10523 5871 10529
rect 5813 10489 5825 10523
rect 5859 10520 5871 10523
rect 6825 10523 6883 10529
rect 5859 10492 6684 10520
rect 5859 10489 5871 10492
rect 5813 10483 5871 10489
rect 6656 10464 6684 10492
rect 6825 10489 6837 10523
rect 6871 10520 6883 10523
rect 7190 10520 7196 10532
rect 6871 10492 7196 10520
rect 6871 10489 6883 10492
rect 6825 10483 6883 10489
rect 7190 10480 7196 10492
rect 7248 10480 7254 10532
rect 8389 10523 8447 10529
rect 8389 10489 8401 10523
rect 8435 10520 8447 10523
rect 8846 10520 8852 10532
rect 8435 10492 8852 10520
rect 8435 10489 8447 10492
rect 8389 10483 8447 10489
rect 6638 10412 6644 10464
rect 6696 10452 6702 10464
rect 8404 10452 8432 10483
rect 8846 10480 8852 10492
rect 8904 10480 8910 10532
rect 6696 10424 8432 10452
rect 6696 10412 6702 10424
rect 1104 10362 13892 10384
rect 1104 10310 3081 10362
rect 3133 10310 3145 10362
rect 3197 10310 3209 10362
rect 3261 10310 3273 10362
rect 3325 10310 3337 10362
rect 3389 10310 7344 10362
rect 7396 10310 7408 10362
rect 7460 10310 7472 10362
rect 7524 10310 7536 10362
rect 7588 10310 7600 10362
rect 7652 10310 11606 10362
rect 11658 10310 11670 10362
rect 11722 10310 11734 10362
rect 11786 10310 11798 10362
rect 11850 10310 11862 10362
rect 11914 10310 13892 10362
rect 1104 10288 13892 10310
rect 3786 10208 3792 10260
rect 3844 10248 3850 10260
rect 4985 10251 5043 10257
rect 4985 10248 4997 10251
rect 3844 10220 4997 10248
rect 3844 10208 3850 10220
rect 4985 10217 4997 10220
rect 5031 10217 5043 10251
rect 5994 10248 6000 10260
rect 5955 10220 6000 10248
rect 4985 10211 5043 10217
rect 5994 10208 6000 10220
rect 6052 10208 6058 10260
rect 8110 10248 8116 10260
rect 6104 10220 8116 10248
rect 5074 10140 5080 10192
rect 5132 10180 5138 10192
rect 6104 10180 6132 10220
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 9493 10251 9551 10257
rect 9493 10217 9505 10251
rect 9539 10248 9551 10251
rect 14001 10251 14059 10257
rect 14001 10248 14013 10251
rect 9539 10220 14013 10248
rect 9539 10217 9551 10220
rect 9493 10211 9551 10217
rect 14001 10217 14013 10220
rect 14047 10217 14059 10251
rect 14001 10211 14059 10217
rect 6822 10180 6828 10192
rect 5132 10152 6132 10180
rect 6196 10152 6828 10180
rect 5132 10140 5138 10152
rect 5169 10047 5227 10053
rect 5169 10013 5181 10047
rect 5215 10044 5227 10047
rect 5994 10044 6000 10056
rect 5215 10016 6000 10044
rect 5215 10013 5227 10016
rect 5169 10007 5227 10013
rect 5994 10004 6000 10016
rect 6052 10004 6058 10056
rect 6196 10053 6224 10152
rect 6822 10140 6828 10152
rect 6880 10180 6886 10192
rect 9858 10180 9864 10192
rect 6880 10152 9864 10180
rect 6880 10140 6886 10152
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 6972 10084 9168 10112
rect 6972 10072 6978 10084
rect 9140 10056 9168 10084
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 6365 10047 6423 10053
rect 6365 10013 6377 10047
rect 6411 10044 6423 10047
rect 7006 10044 7012 10056
rect 6411 10016 7012 10044
rect 6411 10013 6423 10016
rect 6365 10007 6423 10013
rect 7006 10004 7012 10016
rect 7064 10004 7070 10056
rect 9122 10044 9128 10056
rect 9083 10016 9128 10044
rect 9122 10004 9128 10016
rect 9180 10004 9186 10056
rect 5258 9976 5264 9988
rect 5219 9948 5264 9976
rect 5258 9936 5264 9948
rect 5316 9936 5322 9988
rect 5537 9979 5595 9985
rect 5537 9945 5549 9979
rect 5583 9976 5595 9979
rect 6546 9976 6552 9988
rect 5583 9948 6552 9976
rect 5583 9945 5595 9948
rect 5537 9939 5595 9945
rect 6546 9936 6552 9948
rect 6604 9936 6610 9988
rect 8846 9936 8852 9988
rect 8904 9976 8910 9988
rect 8941 9979 8999 9985
rect 8941 9976 8953 9979
rect 8904 9948 8953 9976
rect 8904 9936 8910 9948
rect 8941 9945 8953 9948
rect 8987 9945 8999 9979
rect 8941 9939 8999 9945
rect 9030 9936 9036 9988
rect 9088 9976 9094 9988
rect 9309 9979 9367 9985
rect 9309 9976 9321 9979
rect 9088 9948 9321 9976
rect 9088 9936 9094 9948
rect 9309 9945 9321 9948
rect 9355 9945 9367 9979
rect 9309 9939 9367 9945
rect 5074 9868 5080 9920
rect 5132 9908 5138 9920
rect 5353 9911 5411 9917
rect 5353 9908 5365 9911
rect 5132 9880 5365 9908
rect 5132 9868 5138 9880
rect 5353 9877 5365 9880
rect 5399 9877 5411 9911
rect 5353 9871 5411 9877
rect 6273 9911 6331 9917
rect 6273 9877 6285 9911
rect 6319 9908 6331 9911
rect 6730 9908 6736 9920
rect 6319 9880 6736 9908
rect 6319 9877 6331 9880
rect 6273 9871 6331 9877
rect 6730 9868 6736 9880
rect 6788 9868 6794 9920
rect 9214 9908 9220 9920
rect 9175 9880 9220 9908
rect 9214 9868 9220 9880
rect 9272 9868 9278 9920
rect 1104 9818 13892 9840
rect 1104 9766 5212 9818
rect 5264 9766 5276 9818
rect 5328 9766 5340 9818
rect 5392 9766 5404 9818
rect 5456 9766 5468 9818
rect 5520 9766 9475 9818
rect 9527 9766 9539 9818
rect 9591 9766 9603 9818
rect 9655 9766 9667 9818
rect 9719 9766 9731 9818
rect 9783 9766 13892 9818
rect 1104 9744 13892 9766
rect 5074 9664 5080 9716
rect 5132 9704 5138 9716
rect 5353 9707 5411 9713
rect 5353 9704 5365 9707
rect 5132 9676 5365 9704
rect 5132 9664 5138 9676
rect 5353 9673 5365 9676
rect 5399 9673 5411 9707
rect 5353 9667 5411 9673
rect 4982 9636 4988 9648
rect 4943 9608 4988 9636
rect 4982 9596 4988 9608
rect 5040 9596 5046 9648
rect 5261 9639 5319 9645
rect 5261 9605 5273 9639
rect 5307 9636 5319 9639
rect 8202 9636 8208 9648
rect 5307 9608 8208 9636
rect 5307 9605 5319 9608
rect 5261 9599 5319 9605
rect 8202 9596 8208 9608
rect 8260 9596 8266 9648
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9537 5227 9571
rect 5169 9531 5227 9537
rect 5184 9364 5212 9531
rect 6822 9528 6828 9580
rect 6880 9568 6886 9580
rect 6914 9568 6920 9580
rect 6880 9540 6920 9568
rect 6880 9528 6886 9540
rect 6914 9528 6920 9540
rect 6972 9568 6978 9580
rect 7469 9571 7527 9577
rect 7469 9568 7481 9571
rect 6972 9540 7481 9568
rect 6972 9528 6978 9540
rect 7469 9537 7481 9540
rect 7515 9537 7527 9571
rect 7469 9531 7527 9537
rect 8018 9528 8024 9580
rect 8076 9568 8082 9580
rect 8113 9571 8171 9577
rect 8113 9568 8125 9571
rect 8076 9540 8125 9568
rect 8076 9528 8082 9540
rect 8113 9537 8125 9540
rect 8159 9537 8171 9571
rect 8113 9531 8171 9537
rect 10042 9528 10048 9580
rect 10100 9568 10106 9580
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 10100 9540 13001 9568
rect 10100 9528 10106 9540
rect 12989 9537 13001 9540
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 5537 9435 5595 9441
rect 5537 9401 5549 9435
rect 5583 9432 5595 9435
rect 6546 9432 6552 9444
rect 5583 9404 6552 9432
rect 5583 9401 5595 9404
rect 5537 9395 5595 9401
rect 6546 9392 6552 9404
rect 6604 9432 6610 9444
rect 13170 9432 13176 9444
rect 6604 9404 8340 9432
rect 13131 9404 13176 9432
rect 6604 9392 6610 9404
rect 8312 9376 8340 9404
rect 13170 9392 13176 9404
rect 13228 9392 13234 9444
rect 7653 9367 7711 9373
rect 7653 9364 7665 9367
rect 5184 9336 7665 9364
rect 7653 9333 7665 9336
rect 7699 9364 7711 9367
rect 7742 9364 7748 9376
rect 7699 9336 7748 9364
rect 7699 9333 7711 9336
rect 7653 9327 7711 9333
rect 7742 9324 7748 9336
rect 7800 9324 7806 9376
rect 8294 9364 8300 9376
rect 8255 9336 8300 9364
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 1104 9274 13892 9296
rect 1104 9222 3081 9274
rect 3133 9222 3145 9274
rect 3197 9222 3209 9274
rect 3261 9222 3273 9274
rect 3325 9222 3337 9274
rect 3389 9222 7344 9274
rect 7396 9222 7408 9274
rect 7460 9222 7472 9274
rect 7524 9222 7536 9274
rect 7588 9222 7600 9274
rect 7652 9222 11606 9274
rect 11658 9222 11670 9274
rect 11722 9222 11734 9274
rect 11786 9222 11798 9274
rect 11850 9222 11862 9274
rect 11914 9222 13892 9274
rect 1104 9200 13892 9222
rect 5994 9120 6000 9172
rect 6052 9160 6058 9172
rect 7098 9160 7104 9172
rect 6052 9132 7104 9160
rect 6052 9120 6058 9132
rect 7098 9120 7104 9132
rect 7156 9120 7162 9172
rect 10042 9160 10048 9172
rect 10003 9132 10048 9160
rect 10042 9120 10048 9132
rect 10100 9120 10106 9172
rect 5534 9052 5540 9104
rect 5592 9092 5598 9104
rect 8386 9092 8392 9104
rect 5592 9064 8392 9092
rect 5592 9052 5598 9064
rect 8386 9052 8392 9064
rect 8444 9092 8450 9104
rect 9214 9092 9220 9104
rect 8444 9064 9220 9092
rect 8444 9052 8450 9064
rect 9214 9052 9220 9064
rect 9272 9092 9278 9104
rect 9493 9095 9551 9101
rect 9493 9092 9505 9095
rect 9272 9064 9505 9092
rect 9272 9052 9278 9064
rect 9493 9061 9505 9064
rect 9539 9061 9551 9095
rect 9493 9055 9551 9061
rect 6454 8916 6460 8968
rect 6512 8956 6518 8968
rect 6822 8956 6828 8968
rect 6512 8928 6828 8956
rect 6512 8916 6518 8928
rect 6822 8916 6828 8928
rect 6880 8956 6886 8968
rect 7009 8959 7067 8965
rect 7009 8956 7021 8959
rect 6880 8928 7021 8956
rect 6880 8916 6886 8928
rect 7009 8925 7021 8928
rect 7055 8925 7067 8959
rect 7009 8919 7067 8925
rect 7837 8959 7895 8965
rect 7837 8925 7849 8959
rect 7883 8956 7895 8959
rect 8018 8956 8024 8968
rect 7883 8928 8024 8956
rect 7883 8925 7895 8928
rect 7837 8919 7895 8925
rect 8018 8916 8024 8928
rect 8076 8956 8082 8968
rect 9769 8959 9827 8965
rect 9769 8956 9781 8959
rect 8076 8928 9781 8956
rect 8076 8916 8082 8928
rect 9769 8925 9781 8928
rect 9815 8956 9827 8959
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 9815 8928 14105 8956
rect 9815 8925 9827 8928
rect 9769 8919 9827 8925
rect 14093 8925 14105 8928
rect 14139 8925 14151 8959
rect 14093 8919 14151 8925
rect 6914 8848 6920 8900
rect 6972 8888 6978 8900
rect 7190 8888 7196 8900
rect 6972 8860 7196 8888
rect 6972 8848 6978 8860
rect 7190 8848 7196 8860
rect 7248 8888 7254 8900
rect 7745 8891 7803 8897
rect 7745 8888 7757 8891
rect 7248 8860 7757 8888
rect 7248 8848 7254 8860
rect 7745 8857 7757 8860
rect 7791 8857 7803 8891
rect 7745 8851 7803 8857
rect 7098 8820 7104 8832
rect 7011 8792 7104 8820
rect 7098 8780 7104 8792
rect 7156 8820 7162 8832
rect 8938 8820 8944 8832
rect 7156 8792 8944 8820
rect 7156 8780 7162 8792
rect 8938 8780 8944 8792
rect 8996 8780 9002 8832
rect 9030 8780 9036 8832
rect 9088 8820 9094 8832
rect 9677 8823 9735 8829
rect 9677 8820 9689 8823
rect 9088 8792 9689 8820
rect 9088 8780 9094 8792
rect 9677 8789 9689 8792
rect 9723 8789 9735 8823
rect 9677 8783 9735 8789
rect 9861 8823 9919 8829
rect 9861 8789 9873 8823
rect 9907 8820 9919 8823
rect 9950 8820 9956 8832
rect 9907 8792 9956 8820
rect 9907 8789 9919 8792
rect 9861 8783 9919 8789
rect 9950 8780 9956 8792
rect 10008 8780 10014 8832
rect 1104 8730 13892 8752
rect 1104 8678 5212 8730
rect 5264 8678 5276 8730
rect 5328 8678 5340 8730
rect 5392 8678 5404 8730
rect 5456 8678 5468 8730
rect 5520 8678 9475 8730
rect 9527 8678 9539 8730
rect 9591 8678 9603 8730
rect 9655 8678 9667 8730
rect 9719 8678 9731 8730
rect 9783 8678 13892 8730
rect 1104 8656 13892 8678
rect 5261 8619 5319 8625
rect 5261 8585 5273 8619
rect 5307 8616 5319 8619
rect 5534 8616 5540 8628
rect 5307 8588 5540 8616
rect 5307 8585 5319 8588
rect 5261 8579 5319 8585
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 8386 8616 8392 8628
rect 8347 8588 8392 8616
rect 8386 8576 8392 8588
rect 8444 8576 8450 8628
rect 5169 8551 5227 8557
rect 5169 8517 5181 8551
rect 5215 8548 5227 8551
rect 7742 8548 7748 8560
rect 5215 8520 7748 8548
rect 5215 8517 5227 8520
rect 5169 8511 5227 8517
rect 7742 8508 7748 8520
rect 7800 8508 7806 8560
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8449 5411 8483
rect 5353 8443 5411 8449
rect 5368 8412 5396 8443
rect 6914 8440 6920 8492
rect 6972 8480 6978 8492
rect 6972 8452 7017 8480
rect 6972 8440 6978 8452
rect 7098 8440 7104 8492
rect 7156 8480 7162 8492
rect 7561 8483 7619 8489
rect 7561 8480 7573 8483
rect 7156 8452 7573 8480
rect 7156 8440 7162 8452
rect 7561 8449 7573 8452
rect 7607 8480 7619 8483
rect 7834 8480 7840 8492
rect 7607 8452 7840 8480
rect 7607 8449 7619 8452
rect 7561 8443 7619 8449
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 8202 8480 8208 8492
rect 8163 8452 8208 8480
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 8849 8483 8907 8489
rect 8849 8449 8861 8483
rect 8895 8480 8907 8483
rect 8938 8480 8944 8492
rect 8895 8452 8944 8480
rect 8895 8449 8907 8452
rect 8849 8443 8907 8449
rect 8938 8440 8944 8452
rect 8996 8440 9002 8492
rect 9122 8412 9128 8424
rect 5368 8384 9128 8412
rect 5537 8347 5595 8353
rect 5537 8313 5549 8347
rect 5583 8344 5595 8347
rect 6638 8344 6644 8356
rect 5583 8316 6644 8344
rect 5583 8313 5595 8316
rect 5537 8307 5595 8313
rect 6638 8304 6644 8316
rect 6696 8344 6702 8356
rect 7760 8353 7788 8384
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 7101 8347 7159 8353
rect 7101 8344 7113 8347
rect 6696 8316 7113 8344
rect 6696 8304 6702 8316
rect 7101 8313 7113 8316
rect 7147 8313 7159 8347
rect 7101 8307 7159 8313
rect 7745 8347 7803 8353
rect 7745 8313 7757 8347
rect 7791 8313 7803 8347
rect 7745 8307 7803 8313
rect 8294 8304 8300 8356
rect 8352 8344 8358 8356
rect 9030 8344 9036 8356
rect 8352 8316 9036 8344
rect 8352 8304 8358 8316
rect 9030 8304 9036 8316
rect 9088 8304 9094 8356
rect 4982 8276 4988 8288
rect 4943 8248 4988 8276
rect 4982 8236 4988 8248
rect 5040 8236 5046 8288
rect 1104 8186 13892 8208
rect 1104 8134 3081 8186
rect 3133 8134 3145 8186
rect 3197 8134 3209 8186
rect 3261 8134 3273 8186
rect 3325 8134 3337 8186
rect 3389 8134 7344 8186
rect 7396 8134 7408 8186
rect 7460 8134 7472 8186
rect 7524 8134 7536 8186
rect 7588 8134 7600 8186
rect 7652 8134 11606 8186
rect 11658 8134 11670 8186
rect 11722 8134 11734 8186
rect 11786 8134 11798 8186
rect 11850 8134 11862 8186
rect 11914 8134 13892 8186
rect 1104 8112 13892 8134
rect 7834 8072 7840 8084
rect 7795 8044 7840 8072
rect 7834 8032 7840 8044
rect 7892 8032 7898 8084
rect 5626 7964 5632 8016
rect 5684 8004 5690 8016
rect 8294 8004 8300 8016
rect 5684 7976 8300 8004
rect 5684 7964 5690 7976
rect 8294 7964 8300 7976
rect 8352 7964 8358 8016
rect 7101 7939 7159 7945
rect 7101 7905 7113 7939
rect 7147 7936 7159 7939
rect 8202 7936 8208 7948
rect 7147 7908 8208 7936
rect 7147 7905 7159 7908
rect 7101 7899 7159 7905
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7868 1639 7871
rect 4982 7868 4988 7880
rect 1627 7840 4988 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 4982 7828 4988 7840
rect 5040 7828 5046 7880
rect 6730 7828 6736 7880
rect 6788 7868 6794 7880
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 6788 7840 7021 7868
rect 6788 7828 6794 7840
rect 7009 7837 7021 7840
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7868 7987 7871
rect 8294 7868 8300 7880
rect 7975 7840 8300 7868
rect 7975 7837 7987 7840
rect 7929 7831 7987 7837
rect 8294 7828 8300 7840
rect 8352 7828 8358 7880
rect 1486 7732 1492 7744
rect 1447 7704 1492 7732
rect 1486 7692 1492 7704
rect 1544 7692 1550 7744
rect 1104 7642 13892 7664
rect 1104 7590 5212 7642
rect 5264 7590 5276 7642
rect 5328 7590 5340 7642
rect 5392 7590 5404 7642
rect 5456 7590 5468 7642
rect 5520 7590 9475 7642
rect 9527 7590 9539 7642
rect 9591 7590 9603 7642
rect 9655 7590 9667 7642
rect 9719 7590 9731 7642
rect 9783 7590 13892 7642
rect 1104 7568 13892 7590
rect 5445 7531 5503 7537
rect 5445 7497 5457 7531
rect 5491 7528 5503 7531
rect 7006 7528 7012 7540
rect 5491 7500 7012 7528
rect 5491 7497 5503 7500
rect 5445 7491 5503 7497
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 7193 7531 7251 7537
rect 7193 7497 7205 7531
rect 7239 7528 7251 7531
rect 7834 7528 7840 7540
rect 7239 7500 7840 7528
rect 7239 7497 7251 7500
rect 7193 7491 7251 7497
rect 7834 7488 7840 7500
rect 7892 7488 7898 7540
rect 7929 7531 7987 7537
rect 7929 7497 7941 7531
rect 7975 7528 7987 7531
rect 8110 7528 8116 7540
rect 7975 7500 8116 7528
rect 7975 7497 7987 7500
rect 7929 7491 7987 7497
rect 8110 7488 8116 7500
rect 8168 7528 8174 7540
rect 9125 7531 9183 7537
rect 9125 7528 9137 7531
rect 8168 7500 9137 7528
rect 8168 7488 8174 7500
rect 9125 7497 9137 7500
rect 9171 7497 9183 7531
rect 9125 7491 9183 7497
rect 5626 7460 5632 7472
rect 5587 7432 5632 7460
rect 5626 7420 5632 7432
rect 5684 7460 5690 7472
rect 5902 7460 5908 7472
rect 5684 7432 5908 7460
rect 5684 7420 5690 7432
rect 5902 7420 5908 7432
rect 5960 7420 5966 7472
rect 7852 7460 7880 7488
rect 7852 7432 8432 7460
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 5552 7324 5580 7355
rect 6730 7352 6736 7404
rect 6788 7392 6794 7404
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 6788 7364 7021 7392
rect 6788 7352 6794 7364
rect 7009 7361 7021 7364
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 7745 7395 7803 7401
rect 7745 7361 7757 7395
rect 7791 7392 7803 7395
rect 8294 7392 8300 7404
rect 7791 7364 8300 7392
rect 7791 7361 7803 7364
rect 7745 7355 7803 7361
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 8404 7392 8432 7432
rect 8846 7420 8852 7472
rect 8904 7460 8910 7472
rect 8941 7463 8999 7469
rect 8941 7460 8953 7463
rect 8904 7432 8953 7460
rect 8904 7420 8910 7432
rect 8941 7429 8953 7432
rect 8987 7429 8999 7463
rect 8941 7423 8999 7429
rect 9030 7420 9036 7472
rect 9088 7460 9094 7472
rect 9309 7463 9367 7469
rect 9309 7460 9321 7463
rect 9088 7432 9321 7460
rect 9088 7420 9094 7432
rect 9309 7429 9321 7432
rect 9355 7429 9367 7463
rect 9309 7423 9367 7429
rect 9217 7395 9275 7401
rect 9217 7392 9229 7395
rect 8404 7364 9229 7392
rect 8956 7336 8984 7364
rect 9217 7361 9229 7364
rect 9263 7361 9275 7395
rect 9217 7355 9275 7361
rect 8018 7324 8024 7336
rect 5552 7296 8024 7324
rect 8018 7284 8024 7296
rect 8076 7284 8082 7336
rect 8938 7284 8944 7336
rect 8996 7284 9002 7336
rect 5534 7216 5540 7268
rect 5592 7256 5598 7268
rect 5813 7259 5871 7265
rect 5813 7256 5825 7259
rect 5592 7228 5825 7256
rect 5592 7216 5598 7228
rect 5813 7225 5825 7228
rect 5859 7225 5871 7259
rect 5813 7219 5871 7225
rect 4154 7148 4160 7200
rect 4212 7188 4218 7200
rect 5261 7191 5319 7197
rect 5261 7188 5273 7191
rect 4212 7160 5273 7188
rect 4212 7148 4218 7160
rect 5261 7157 5273 7160
rect 5307 7157 5319 7191
rect 5261 7151 5319 7157
rect 9493 7191 9551 7197
rect 9493 7157 9505 7191
rect 9539 7188 9551 7191
rect 12986 7188 12992 7200
rect 9539 7160 12992 7188
rect 9539 7157 9551 7160
rect 9493 7151 9551 7157
rect 12986 7148 12992 7160
rect 13044 7148 13050 7200
rect 1104 7098 13892 7120
rect 1104 7046 3081 7098
rect 3133 7046 3145 7098
rect 3197 7046 3209 7098
rect 3261 7046 3273 7098
rect 3325 7046 3337 7098
rect 3389 7046 7344 7098
rect 7396 7046 7408 7098
rect 7460 7046 7472 7098
rect 7524 7046 7536 7098
rect 7588 7046 7600 7098
rect 7652 7046 11606 7098
rect 11658 7046 11670 7098
rect 11722 7046 11734 7098
rect 11786 7046 11798 7098
rect 11850 7046 11862 7098
rect 11914 7046 13892 7098
rect 1104 7024 13892 7046
rect 8294 6808 8300 6860
rect 8352 6848 8358 6860
rect 9950 6848 9956 6860
rect 8352 6820 9956 6848
rect 8352 6808 8358 6820
rect 9950 6808 9956 6820
rect 10008 6808 10014 6860
rect 1104 6554 13892 6576
rect 1104 6502 5212 6554
rect 5264 6502 5276 6554
rect 5328 6502 5340 6554
rect 5392 6502 5404 6554
rect 5456 6502 5468 6554
rect 5520 6502 9475 6554
rect 9527 6502 9539 6554
rect 9591 6502 9603 6554
rect 9655 6502 9667 6554
rect 9719 6502 9731 6554
rect 9783 6502 13892 6554
rect 1104 6480 13892 6502
rect 5074 6400 5080 6452
rect 5132 6440 5138 6452
rect 5261 6443 5319 6449
rect 5261 6440 5273 6443
rect 5132 6412 5273 6440
rect 5132 6400 5138 6412
rect 5261 6409 5273 6412
rect 5307 6409 5319 6443
rect 5261 6403 5319 6409
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 6733 6443 6791 6449
rect 6733 6440 6745 6443
rect 5960 6412 6745 6440
rect 5960 6400 5966 6412
rect 6733 6409 6745 6412
rect 6779 6409 6791 6443
rect 7742 6440 7748 6452
rect 7703 6412 7748 6440
rect 6733 6403 6791 6409
rect 7742 6400 7748 6412
rect 7800 6400 7806 6452
rect 9030 6440 9036 6452
rect 8991 6412 9036 6440
rect 9030 6400 9036 6412
rect 9088 6400 9094 6452
rect 6454 6372 6460 6384
rect 5092 6344 6460 6372
rect 5092 6313 5120 6344
rect 6454 6332 6460 6344
rect 6512 6332 6518 6384
rect 6549 6375 6607 6381
rect 6549 6341 6561 6375
rect 6595 6372 6607 6375
rect 7653 6375 7711 6381
rect 6595 6344 7328 6372
rect 6595 6341 6607 6344
rect 6549 6335 6607 6341
rect 5077 6307 5135 6313
rect 5077 6273 5089 6307
rect 5123 6273 5135 6307
rect 5077 6267 5135 6273
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6304 5227 6307
rect 5350 6304 5356 6316
rect 5215 6276 5356 6304
rect 5215 6273 5227 6276
rect 5169 6267 5227 6273
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 5445 6307 5503 6313
rect 5445 6273 5457 6307
rect 5491 6304 5503 6307
rect 6641 6307 6699 6313
rect 6641 6304 6653 6307
rect 5491 6276 6653 6304
rect 5491 6273 5503 6276
rect 5445 6267 5503 6273
rect 6641 6273 6653 6276
rect 6687 6304 6699 6307
rect 6914 6304 6920 6316
rect 6687 6276 6920 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 6914 6264 6920 6276
rect 6972 6264 6978 6316
rect 2866 6196 2872 6248
rect 2924 6236 2930 6248
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 2924 6208 6377 6236
rect 2924 6196 2930 6208
rect 6365 6205 6377 6208
rect 6411 6205 6423 6239
rect 6365 6199 6423 6205
rect 5534 6128 5540 6180
rect 5592 6168 5598 6180
rect 6917 6171 6975 6177
rect 6917 6168 6929 6171
rect 5592 6140 6929 6168
rect 5592 6128 5598 6140
rect 6917 6137 6929 6140
rect 6963 6137 6975 6171
rect 7300 6168 7328 6344
rect 7653 6341 7665 6375
rect 7699 6372 7711 6375
rect 8202 6372 8208 6384
rect 7699 6344 8208 6372
rect 7699 6341 7711 6344
rect 7653 6335 7711 6341
rect 8202 6332 8208 6344
rect 8260 6332 8266 6384
rect 8938 6372 8944 6384
rect 8899 6344 8944 6372
rect 8938 6332 8944 6344
rect 8996 6332 9002 6384
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6304 7619 6307
rect 8849 6307 8907 6313
rect 8849 6304 8861 6307
rect 7607 6276 8861 6304
rect 7607 6273 7619 6276
rect 7561 6267 7619 6273
rect 8849 6273 8861 6276
rect 8895 6304 8907 6307
rect 9122 6304 9128 6316
rect 8895 6276 9128 6304
rect 8895 6273 8907 6276
rect 8849 6267 8907 6273
rect 9122 6264 9128 6276
rect 9180 6264 9186 6316
rect 7377 6239 7435 6245
rect 7377 6205 7389 6239
rect 7423 6236 7435 6239
rect 8386 6236 8392 6248
rect 7423 6208 8392 6236
rect 7423 6205 7435 6208
rect 7377 6199 7435 6205
rect 8386 6196 8392 6208
rect 8444 6236 8450 6248
rect 8665 6239 8723 6245
rect 8665 6236 8677 6239
rect 8444 6208 8677 6236
rect 8444 6196 8450 6208
rect 8665 6205 8677 6208
rect 8711 6205 8723 6239
rect 8665 6199 8723 6205
rect 8294 6168 8300 6180
rect 7300 6140 8300 6168
rect 6917 6131 6975 6137
rect 8294 6128 8300 6140
rect 8352 6128 8358 6180
rect 4890 6100 4896 6112
rect 4851 6072 4896 6100
rect 4890 6060 4896 6072
rect 4948 6060 4954 6112
rect 7929 6103 7987 6109
rect 7929 6069 7941 6103
rect 7975 6100 7987 6103
rect 8202 6100 8208 6112
rect 7975 6072 8208 6100
rect 7975 6069 7987 6072
rect 7929 6063 7987 6069
rect 8202 6060 8208 6072
rect 8260 6060 8266 6112
rect 9217 6103 9275 6109
rect 9217 6069 9229 6103
rect 9263 6100 9275 6103
rect 14001 6103 14059 6109
rect 14001 6100 14013 6103
rect 9263 6072 14013 6100
rect 9263 6069 9275 6072
rect 9217 6063 9275 6069
rect 14001 6069 14013 6072
rect 14047 6069 14059 6103
rect 14001 6063 14059 6069
rect 1104 6010 13892 6032
rect 1104 5958 3081 6010
rect 3133 5958 3145 6010
rect 3197 5958 3209 6010
rect 3261 5958 3273 6010
rect 3325 5958 3337 6010
rect 3389 5958 7344 6010
rect 7396 5958 7408 6010
rect 7460 5958 7472 6010
rect 7524 5958 7536 6010
rect 7588 5958 7600 6010
rect 7652 5958 11606 6010
rect 11658 5958 11670 6010
rect 11722 5958 11734 6010
rect 11786 5958 11798 6010
rect 11850 5958 11862 6010
rect 11914 5958 13892 6010
rect 1104 5936 13892 5958
rect 8110 5788 8116 5840
rect 8168 5828 8174 5840
rect 8941 5831 8999 5837
rect 8941 5828 8953 5831
rect 8168 5800 8953 5828
rect 8168 5788 8174 5800
rect 8941 5797 8953 5800
rect 8987 5797 8999 5831
rect 8941 5791 8999 5797
rect 5534 5720 5540 5772
rect 5592 5760 5598 5772
rect 6822 5760 6828 5772
rect 5592 5732 6828 5760
rect 5592 5720 5598 5732
rect 6822 5720 6828 5732
rect 6880 5760 6886 5772
rect 6880 5732 9260 5760
rect 6880 5720 6886 5732
rect 9232 5701 9260 5732
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5661 9275 5695
rect 12986 5692 12992 5704
rect 12947 5664 12992 5692
rect 9217 5655 9275 5661
rect 12986 5652 12992 5664
rect 13044 5652 13050 5704
rect 9309 5627 9367 5633
rect 9309 5624 9321 5627
rect 9048 5596 9321 5624
rect 6454 5516 6460 5568
rect 6512 5556 6518 5568
rect 9048 5556 9076 5596
rect 9309 5593 9321 5596
rect 9355 5593 9367 5627
rect 9950 5624 9956 5636
rect 9309 5587 9367 5593
rect 9416 5596 9956 5624
rect 6512 5528 9076 5556
rect 9125 5559 9183 5565
rect 6512 5516 6518 5528
rect 9125 5525 9137 5559
rect 9171 5556 9183 5559
rect 9416 5556 9444 5596
rect 9950 5584 9956 5596
rect 10008 5624 10014 5636
rect 14093 5627 14151 5633
rect 14093 5624 14105 5627
rect 10008 5596 14105 5624
rect 10008 5584 10014 5596
rect 14093 5593 14105 5596
rect 14139 5593 14151 5627
rect 14093 5587 14151 5593
rect 9171 5528 9444 5556
rect 9493 5559 9551 5565
rect 9171 5525 9183 5528
rect 9125 5519 9183 5525
rect 9493 5525 9505 5559
rect 9539 5556 9551 5559
rect 10778 5556 10784 5568
rect 9539 5528 10784 5556
rect 9539 5525 9551 5528
rect 9493 5519 9551 5525
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 13078 5556 13084 5568
rect 13039 5528 13084 5556
rect 13078 5516 13084 5528
rect 13136 5516 13142 5568
rect 1104 5466 13892 5488
rect 1104 5414 5212 5466
rect 5264 5414 5276 5466
rect 5328 5414 5340 5466
rect 5392 5414 5404 5466
rect 5456 5414 5468 5466
rect 5520 5414 9475 5466
rect 9527 5414 9539 5466
rect 9591 5414 9603 5466
rect 9655 5414 9667 5466
rect 9719 5414 9731 5466
rect 9783 5414 13892 5466
rect 1104 5392 13892 5414
rect 1104 4922 13892 4944
rect 1104 4870 3081 4922
rect 3133 4870 3145 4922
rect 3197 4870 3209 4922
rect 3261 4870 3273 4922
rect 3325 4870 3337 4922
rect 3389 4870 7344 4922
rect 7396 4870 7408 4922
rect 7460 4870 7472 4922
rect 7524 4870 7536 4922
rect 7588 4870 7600 4922
rect 7652 4870 11606 4922
rect 11658 4870 11670 4922
rect 11722 4870 11734 4922
rect 11786 4870 11798 4922
rect 11850 4870 11862 4922
rect 11914 4870 13892 4922
rect 1104 4848 13892 4870
rect 1104 4378 13892 4400
rect 1104 4326 5212 4378
rect 5264 4326 5276 4378
rect 5328 4326 5340 4378
rect 5392 4326 5404 4378
rect 5456 4326 5468 4378
rect 5520 4326 9475 4378
rect 9527 4326 9539 4378
rect 9591 4326 9603 4378
rect 9655 4326 9667 4378
rect 9719 4326 9731 4378
rect 9783 4326 13892 4378
rect 1104 4304 13892 4326
rect 1581 4199 1639 4205
rect 1581 4165 1593 4199
rect 1627 4196 1639 4199
rect 4154 4196 4160 4208
rect 1627 4168 4160 4196
rect 1627 4165 1639 4168
rect 1581 4159 1639 4165
rect 4154 4156 4160 4168
rect 4212 4156 4218 4208
rect 1486 3924 1492 3936
rect 1447 3896 1492 3924
rect 1486 3884 1492 3896
rect 1544 3884 1550 3936
rect 1104 3834 13892 3856
rect 1104 3782 3081 3834
rect 3133 3782 3145 3834
rect 3197 3782 3209 3834
rect 3261 3782 3273 3834
rect 3325 3782 3337 3834
rect 3389 3782 7344 3834
rect 7396 3782 7408 3834
rect 7460 3782 7472 3834
rect 7524 3782 7536 3834
rect 7588 3782 7600 3834
rect 7652 3782 11606 3834
rect 11658 3782 11670 3834
rect 11722 3782 11734 3834
rect 11786 3782 11798 3834
rect 11850 3782 11862 3834
rect 11914 3782 13892 3834
rect 1104 3760 13892 3782
rect 1104 3290 13892 3312
rect 1104 3238 5212 3290
rect 5264 3238 5276 3290
rect 5328 3238 5340 3290
rect 5392 3238 5404 3290
rect 5456 3238 5468 3290
rect 5520 3238 9475 3290
rect 9527 3238 9539 3290
rect 9591 3238 9603 3290
rect 9655 3238 9667 3290
rect 9719 3238 9731 3290
rect 9783 3238 13892 3290
rect 1104 3216 13892 3238
rect 12989 3111 13047 3117
rect 12989 3077 13001 3111
rect 13035 3108 13047 3111
rect 14001 3111 14059 3117
rect 14001 3108 14013 3111
rect 13035 3080 14013 3108
rect 13035 3077 13047 3080
rect 12989 3071 13047 3077
rect 14001 3077 14013 3080
rect 14047 3077 14059 3111
rect 14001 3071 14059 3077
rect 13173 2907 13231 2913
rect 13173 2873 13185 2907
rect 13219 2904 13231 2907
rect 13262 2904 13268 2916
rect 13219 2876 13268 2904
rect 13219 2873 13231 2876
rect 13173 2867 13231 2873
rect 13262 2864 13268 2876
rect 13320 2864 13326 2916
rect 1104 2746 13892 2768
rect 1104 2694 3081 2746
rect 3133 2694 3145 2746
rect 3197 2694 3209 2746
rect 3261 2694 3273 2746
rect 3325 2694 3337 2746
rect 3389 2694 7344 2746
rect 7396 2694 7408 2746
rect 7460 2694 7472 2746
rect 7524 2694 7536 2746
rect 7588 2694 7600 2746
rect 7652 2694 11606 2746
rect 11658 2694 11670 2746
rect 11722 2694 11734 2746
rect 11786 2694 11798 2746
rect 11850 2694 11862 2746
rect 11914 2694 13892 2746
rect 1104 2672 13892 2694
rect 5534 2592 5540 2644
rect 5592 2632 5598 2644
rect 5629 2635 5687 2641
rect 5629 2632 5641 2635
rect 5592 2604 5641 2632
rect 5592 2592 5598 2604
rect 5629 2601 5641 2604
rect 5675 2601 5687 2635
rect 5629 2595 5687 2601
rect 12989 2635 13047 2641
rect 12989 2601 13001 2635
rect 13035 2632 13047 2635
rect 14093 2635 14151 2641
rect 14093 2632 14105 2635
rect 13035 2604 14105 2632
rect 13035 2601 13047 2604
rect 12989 2595 13047 2601
rect 14093 2601 14105 2604
rect 14139 2601 14151 2635
rect 14093 2595 14151 2601
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2428 1639 2431
rect 4890 2428 4896 2440
rect 1627 2400 4896 2428
rect 1627 2397 1639 2400
rect 1581 2391 1639 2397
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 8202 2428 8208 2440
rect 8163 2400 8208 2428
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 10778 2388 10784 2440
rect 10836 2428 10842 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 10836 2400 11713 2428
rect 10836 2388 10842 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 920 2360 926 2372
rect 917 2332 926 2360
rect 920 2320 926 2332
rect 978 2360 984 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 978 2332 1409 2360
rect 978 2320 984 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 2590 2320 2596 2372
rect 2648 2360 2654 2372
rect 2685 2363 2743 2369
rect 2685 2360 2697 2363
rect 2648 2332 2697 2360
rect 2648 2320 2654 2332
rect 2685 2329 2697 2332
rect 2731 2329 2743 2363
rect 2866 2360 2872 2372
rect 2827 2332 2872 2360
rect 2685 2323 2743 2329
rect 2866 2320 2872 2332
rect 2924 2320 2930 2372
rect 5534 2360 5540 2372
rect 5495 2332 5540 2360
rect 5534 2320 5540 2332
rect 5592 2320 5598 2372
rect 7926 2320 7932 2372
rect 7984 2360 7990 2372
rect 8021 2363 8079 2369
rect 8021 2360 8033 2363
rect 7984 2332 8033 2360
rect 7984 2320 7990 2332
rect 8021 2329 8033 2332
rect 8067 2329 8079 2363
rect 8021 2323 8079 2329
rect 10686 2320 10692 2372
rect 10744 2360 10750 2372
rect 11517 2363 11575 2369
rect 11517 2360 11529 2363
rect 10744 2332 11529 2360
rect 10744 2320 10750 2332
rect 11517 2329 11529 2332
rect 11563 2329 11575 2363
rect 13078 2360 13084 2372
rect 13039 2332 13084 2360
rect 11517 2323 11575 2329
rect 13078 2320 13084 2332
rect 13136 2320 13142 2372
rect 1104 2202 13892 2224
rect 1104 2150 5212 2202
rect 5264 2150 5276 2202
rect 5328 2150 5340 2202
rect 5392 2150 5404 2202
rect 5456 2150 5468 2202
rect 5520 2150 9475 2202
rect 9527 2150 9539 2202
rect 9591 2150 9603 2202
rect 9655 2150 9667 2202
rect 9719 2150 9731 2202
rect 9783 2150 13892 2202
rect 1104 2128 13892 2150
<< via1 >>
rect 3081 14662 3133 14714
rect 3145 14662 3197 14714
rect 3209 14662 3261 14714
rect 3273 14662 3325 14714
rect 3337 14662 3389 14714
rect 7344 14662 7396 14714
rect 7408 14662 7460 14714
rect 7472 14662 7524 14714
rect 7536 14662 7588 14714
rect 7600 14662 7652 14714
rect 11606 14662 11658 14714
rect 11670 14662 11722 14714
rect 11734 14662 11786 14714
rect 11798 14662 11850 14714
rect 11862 14662 11914 14714
rect 1492 14603 1544 14612
rect 1492 14569 1501 14603
rect 1501 14569 1535 14603
rect 1535 14569 1544 14603
rect 1492 14560 1544 14569
rect 1676 14492 1728 14544
rect 4252 14492 4304 14544
rect 7012 14492 7064 14544
rect 12348 14492 12400 14544
rect 3792 14356 3844 14408
rect 7196 14356 7248 14408
rect 9680 14356 9732 14408
rect 14924 14356 14976 14408
rect 4068 14288 4120 14340
rect 6000 14288 6052 14340
rect 12256 14331 12308 14340
rect 12256 14297 12265 14331
rect 12265 14297 12299 14331
rect 12299 14297 12308 14331
rect 12256 14288 12308 14297
rect 9864 14220 9916 14272
rect 5212 14118 5264 14170
rect 5276 14118 5328 14170
rect 5340 14118 5392 14170
rect 5404 14118 5456 14170
rect 5468 14118 5520 14170
rect 9475 14118 9527 14170
rect 9539 14118 9591 14170
rect 9603 14118 9655 14170
rect 9667 14118 9719 14170
rect 9731 14118 9783 14170
rect 3081 13574 3133 13626
rect 3145 13574 3197 13626
rect 3209 13574 3261 13626
rect 3273 13574 3325 13626
rect 3337 13574 3389 13626
rect 7344 13574 7396 13626
rect 7408 13574 7460 13626
rect 7472 13574 7524 13626
rect 7536 13574 7588 13626
rect 7600 13574 7652 13626
rect 11606 13574 11658 13626
rect 11670 13574 11722 13626
rect 11734 13574 11786 13626
rect 11798 13574 11850 13626
rect 11862 13574 11914 13626
rect 13176 13243 13228 13252
rect 13176 13209 13185 13243
rect 13185 13209 13219 13243
rect 13219 13209 13228 13243
rect 13176 13200 13228 13209
rect 5212 13030 5264 13082
rect 5276 13030 5328 13082
rect 5340 13030 5392 13082
rect 5404 13030 5456 13082
rect 5468 13030 5520 13082
rect 9475 13030 9527 13082
rect 9539 13030 9591 13082
rect 9603 13030 9655 13082
rect 9667 13030 9719 13082
rect 9731 13030 9783 13082
rect 3081 12486 3133 12538
rect 3145 12486 3197 12538
rect 3209 12486 3261 12538
rect 3273 12486 3325 12538
rect 3337 12486 3389 12538
rect 7344 12486 7396 12538
rect 7408 12486 7460 12538
rect 7472 12486 7524 12538
rect 7536 12486 7588 12538
rect 7600 12486 7652 12538
rect 11606 12486 11658 12538
rect 11670 12486 11722 12538
rect 11734 12486 11786 12538
rect 11798 12486 11850 12538
rect 11862 12486 11914 12538
rect 4988 12112 5040 12164
rect 1492 12087 1544 12096
rect 1492 12053 1501 12087
rect 1501 12053 1535 12087
rect 1535 12053 1544 12087
rect 1492 12044 1544 12053
rect 5212 11942 5264 11994
rect 5276 11942 5328 11994
rect 5340 11942 5392 11994
rect 5404 11942 5456 11994
rect 5468 11942 5520 11994
rect 9475 11942 9527 11994
rect 9539 11942 9591 11994
rect 9603 11942 9655 11994
rect 9667 11942 9719 11994
rect 9731 11942 9783 11994
rect 3081 11398 3133 11450
rect 3145 11398 3197 11450
rect 3209 11398 3261 11450
rect 3273 11398 3325 11450
rect 3337 11398 3389 11450
rect 7344 11398 7396 11450
rect 7408 11398 7460 11450
rect 7472 11398 7524 11450
rect 7536 11398 7588 11450
rect 7600 11398 7652 11450
rect 11606 11398 11658 11450
rect 11670 11398 11722 11450
rect 11734 11398 11786 11450
rect 11798 11398 11850 11450
rect 11862 11398 11914 11450
rect 5212 10854 5264 10906
rect 5276 10854 5328 10906
rect 5340 10854 5392 10906
rect 5404 10854 5456 10906
rect 5468 10854 5520 10906
rect 9475 10854 9527 10906
rect 9539 10854 9591 10906
rect 9603 10854 9655 10906
rect 9667 10854 9719 10906
rect 9731 10854 9783 10906
rect 4068 10752 4120 10804
rect 6920 10752 6972 10804
rect 7012 10795 7064 10804
rect 7012 10761 7021 10795
rect 7021 10761 7055 10795
rect 7055 10761 7064 10795
rect 7012 10752 7064 10761
rect 7196 10752 7248 10804
rect 12256 10752 12308 10804
rect 8208 10684 8260 10736
rect 5264 10548 5316 10600
rect 5632 10616 5684 10668
rect 7748 10616 7800 10668
rect 8116 10616 8168 10668
rect 7932 10548 7984 10600
rect 7196 10480 7248 10532
rect 6644 10412 6696 10464
rect 8852 10480 8904 10532
rect 3081 10310 3133 10362
rect 3145 10310 3197 10362
rect 3209 10310 3261 10362
rect 3273 10310 3325 10362
rect 3337 10310 3389 10362
rect 7344 10310 7396 10362
rect 7408 10310 7460 10362
rect 7472 10310 7524 10362
rect 7536 10310 7588 10362
rect 7600 10310 7652 10362
rect 11606 10310 11658 10362
rect 11670 10310 11722 10362
rect 11734 10310 11786 10362
rect 11798 10310 11850 10362
rect 11862 10310 11914 10362
rect 3792 10208 3844 10260
rect 6000 10251 6052 10260
rect 6000 10217 6009 10251
rect 6009 10217 6043 10251
rect 6043 10217 6052 10251
rect 6000 10208 6052 10217
rect 5080 10140 5132 10192
rect 8116 10208 8168 10260
rect 6000 10004 6052 10056
rect 6828 10140 6880 10192
rect 9864 10140 9916 10192
rect 6920 10072 6972 10124
rect 7012 10004 7064 10056
rect 9128 10047 9180 10056
rect 9128 10013 9137 10047
rect 9137 10013 9171 10047
rect 9171 10013 9180 10047
rect 9128 10004 9180 10013
rect 5264 9979 5316 9988
rect 5264 9945 5273 9979
rect 5273 9945 5307 9979
rect 5307 9945 5316 9979
rect 5264 9936 5316 9945
rect 6552 9979 6604 9988
rect 6552 9945 6561 9979
rect 6561 9945 6595 9979
rect 6595 9945 6604 9979
rect 6552 9936 6604 9945
rect 8852 9936 8904 9988
rect 9036 9936 9088 9988
rect 5080 9868 5132 9920
rect 6736 9868 6788 9920
rect 9220 9911 9272 9920
rect 9220 9877 9229 9911
rect 9229 9877 9263 9911
rect 9263 9877 9272 9911
rect 9220 9868 9272 9877
rect 5212 9766 5264 9818
rect 5276 9766 5328 9818
rect 5340 9766 5392 9818
rect 5404 9766 5456 9818
rect 5468 9766 5520 9818
rect 9475 9766 9527 9818
rect 9539 9766 9591 9818
rect 9603 9766 9655 9818
rect 9667 9766 9719 9818
rect 9731 9766 9783 9818
rect 5080 9664 5132 9716
rect 4988 9639 5040 9648
rect 4988 9605 4997 9639
rect 4997 9605 5031 9639
rect 5031 9605 5040 9639
rect 4988 9596 5040 9605
rect 8208 9596 8260 9648
rect 6828 9528 6880 9580
rect 6920 9528 6972 9580
rect 8024 9528 8076 9580
rect 10048 9528 10100 9580
rect 6552 9392 6604 9444
rect 13176 9435 13228 9444
rect 13176 9401 13185 9435
rect 13185 9401 13219 9435
rect 13219 9401 13228 9435
rect 13176 9392 13228 9401
rect 7748 9324 7800 9376
rect 8300 9367 8352 9376
rect 8300 9333 8309 9367
rect 8309 9333 8343 9367
rect 8343 9333 8352 9367
rect 8300 9324 8352 9333
rect 3081 9222 3133 9274
rect 3145 9222 3197 9274
rect 3209 9222 3261 9274
rect 3273 9222 3325 9274
rect 3337 9222 3389 9274
rect 7344 9222 7396 9274
rect 7408 9222 7460 9274
rect 7472 9222 7524 9274
rect 7536 9222 7588 9274
rect 7600 9222 7652 9274
rect 11606 9222 11658 9274
rect 11670 9222 11722 9274
rect 11734 9222 11786 9274
rect 11798 9222 11850 9274
rect 11862 9222 11914 9274
rect 6000 9120 6052 9172
rect 7104 9120 7156 9172
rect 10048 9163 10100 9172
rect 10048 9129 10057 9163
rect 10057 9129 10091 9163
rect 10091 9129 10100 9163
rect 10048 9120 10100 9129
rect 5540 9052 5592 9104
rect 8392 9052 8444 9104
rect 9220 9052 9272 9104
rect 6460 8916 6512 8968
rect 6828 8916 6880 8968
rect 8024 8916 8076 8968
rect 6920 8848 6972 8900
rect 7196 8848 7248 8900
rect 7104 8823 7156 8832
rect 7104 8789 7113 8823
rect 7113 8789 7147 8823
rect 7147 8789 7156 8823
rect 7104 8780 7156 8789
rect 8944 8780 8996 8832
rect 9036 8780 9088 8832
rect 9956 8780 10008 8832
rect 5212 8678 5264 8730
rect 5276 8678 5328 8730
rect 5340 8678 5392 8730
rect 5404 8678 5456 8730
rect 5468 8678 5520 8730
rect 9475 8678 9527 8730
rect 9539 8678 9591 8730
rect 9603 8678 9655 8730
rect 9667 8678 9719 8730
rect 9731 8678 9783 8730
rect 5540 8576 5592 8628
rect 8392 8619 8444 8628
rect 8392 8585 8401 8619
rect 8401 8585 8435 8619
rect 8435 8585 8444 8619
rect 8392 8576 8444 8585
rect 7748 8508 7800 8560
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 7104 8440 7156 8492
rect 7840 8440 7892 8492
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 8944 8440 8996 8492
rect 6644 8304 6696 8356
rect 9128 8372 9180 8424
rect 8300 8304 8352 8356
rect 9036 8347 9088 8356
rect 9036 8313 9045 8347
rect 9045 8313 9079 8347
rect 9079 8313 9088 8347
rect 9036 8304 9088 8313
rect 4988 8279 5040 8288
rect 4988 8245 4997 8279
rect 4997 8245 5031 8279
rect 5031 8245 5040 8279
rect 4988 8236 5040 8245
rect 3081 8134 3133 8186
rect 3145 8134 3197 8186
rect 3209 8134 3261 8186
rect 3273 8134 3325 8186
rect 3337 8134 3389 8186
rect 7344 8134 7396 8186
rect 7408 8134 7460 8186
rect 7472 8134 7524 8186
rect 7536 8134 7588 8186
rect 7600 8134 7652 8186
rect 11606 8134 11658 8186
rect 11670 8134 11722 8186
rect 11734 8134 11786 8186
rect 11798 8134 11850 8186
rect 11862 8134 11914 8186
rect 7840 8075 7892 8084
rect 7840 8041 7849 8075
rect 7849 8041 7883 8075
rect 7883 8041 7892 8075
rect 7840 8032 7892 8041
rect 5632 7964 5684 8016
rect 8300 7964 8352 8016
rect 8208 7896 8260 7948
rect 4988 7828 5040 7880
rect 6736 7828 6788 7880
rect 8300 7828 8352 7880
rect 1492 7735 1544 7744
rect 1492 7701 1501 7735
rect 1501 7701 1535 7735
rect 1535 7701 1544 7735
rect 1492 7692 1544 7701
rect 5212 7590 5264 7642
rect 5276 7590 5328 7642
rect 5340 7590 5392 7642
rect 5404 7590 5456 7642
rect 5468 7590 5520 7642
rect 9475 7590 9527 7642
rect 9539 7590 9591 7642
rect 9603 7590 9655 7642
rect 9667 7590 9719 7642
rect 9731 7590 9783 7642
rect 7012 7488 7064 7540
rect 7840 7488 7892 7540
rect 8116 7488 8168 7540
rect 5632 7463 5684 7472
rect 5632 7429 5641 7463
rect 5641 7429 5675 7463
rect 5675 7429 5684 7463
rect 5632 7420 5684 7429
rect 5908 7420 5960 7472
rect 6736 7352 6788 7404
rect 8300 7352 8352 7404
rect 8852 7420 8904 7472
rect 9036 7420 9088 7472
rect 8024 7284 8076 7336
rect 8944 7284 8996 7336
rect 5540 7216 5592 7268
rect 4160 7148 4212 7200
rect 12992 7148 13044 7200
rect 3081 7046 3133 7098
rect 3145 7046 3197 7098
rect 3209 7046 3261 7098
rect 3273 7046 3325 7098
rect 3337 7046 3389 7098
rect 7344 7046 7396 7098
rect 7408 7046 7460 7098
rect 7472 7046 7524 7098
rect 7536 7046 7588 7098
rect 7600 7046 7652 7098
rect 11606 7046 11658 7098
rect 11670 7046 11722 7098
rect 11734 7046 11786 7098
rect 11798 7046 11850 7098
rect 11862 7046 11914 7098
rect 8300 6808 8352 6860
rect 9956 6808 10008 6860
rect 5212 6502 5264 6554
rect 5276 6502 5328 6554
rect 5340 6502 5392 6554
rect 5404 6502 5456 6554
rect 5468 6502 5520 6554
rect 9475 6502 9527 6554
rect 9539 6502 9591 6554
rect 9603 6502 9655 6554
rect 9667 6502 9719 6554
rect 9731 6502 9783 6554
rect 5080 6400 5132 6452
rect 5908 6400 5960 6452
rect 7748 6443 7800 6452
rect 7748 6409 7757 6443
rect 7757 6409 7791 6443
rect 7791 6409 7800 6443
rect 7748 6400 7800 6409
rect 9036 6443 9088 6452
rect 9036 6409 9045 6443
rect 9045 6409 9079 6443
rect 9079 6409 9088 6443
rect 9036 6400 9088 6409
rect 6460 6332 6512 6384
rect 5356 6264 5408 6316
rect 6920 6264 6972 6316
rect 2872 6196 2924 6248
rect 5540 6128 5592 6180
rect 8208 6332 8260 6384
rect 8944 6375 8996 6384
rect 8944 6341 8953 6375
rect 8953 6341 8987 6375
rect 8987 6341 8996 6375
rect 8944 6332 8996 6341
rect 9128 6264 9180 6316
rect 8392 6196 8444 6248
rect 8300 6128 8352 6180
rect 4896 6103 4948 6112
rect 4896 6069 4905 6103
rect 4905 6069 4939 6103
rect 4939 6069 4948 6103
rect 4896 6060 4948 6069
rect 8208 6060 8260 6112
rect 3081 5958 3133 6010
rect 3145 5958 3197 6010
rect 3209 5958 3261 6010
rect 3273 5958 3325 6010
rect 3337 5958 3389 6010
rect 7344 5958 7396 6010
rect 7408 5958 7460 6010
rect 7472 5958 7524 6010
rect 7536 5958 7588 6010
rect 7600 5958 7652 6010
rect 11606 5958 11658 6010
rect 11670 5958 11722 6010
rect 11734 5958 11786 6010
rect 11798 5958 11850 6010
rect 11862 5958 11914 6010
rect 8116 5788 8168 5840
rect 5540 5720 5592 5772
rect 6828 5720 6880 5772
rect 12992 5695 13044 5704
rect 12992 5661 13001 5695
rect 13001 5661 13035 5695
rect 13035 5661 13044 5695
rect 12992 5652 13044 5661
rect 6460 5516 6512 5568
rect 9956 5584 10008 5636
rect 10784 5516 10836 5568
rect 13084 5559 13136 5568
rect 13084 5525 13093 5559
rect 13093 5525 13127 5559
rect 13127 5525 13136 5559
rect 13084 5516 13136 5525
rect 5212 5414 5264 5466
rect 5276 5414 5328 5466
rect 5340 5414 5392 5466
rect 5404 5414 5456 5466
rect 5468 5414 5520 5466
rect 9475 5414 9527 5466
rect 9539 5414 9591 5466
rect 9603 5414 9655 5466
rect 9667 5414 9719 5466
rect 9731 5414 9783 5466
rect 3081 4870 3133 4922
rect 3145 4870 3197 4922
rect 3209 4870 3261 4922
rect 3273 4870 3325 4922
rect 3337 4870 3389 4922
rect 7344 4870 7396 4922
rect 7408 4870 7460 4922
rect 7472 4870 7524 4922
rect 7536 4870 7588 4922
rect 7600 4870 7652 4922
rect 11606 4870 11658 4922
rect 11670 4870 11722 4922
rect 11734 4870 11786 4922
rect 11798 4870 11850 4922
rect 11862 4870 11914 4922
rect 5212 4326 5264 4378
rect 5276 4326 5328 4378
rect 5340 4326 5392 4378
rect 5404 4326 5456 4378
rect 5468 4326 5520 4378
rect 9475 4326 9527 4378
rect 9539 4326 9591 4378
rect 9603 4326 9655 4378
rect 9667 4326 9719 4378
rect 9731 4326 9783 4378
rect 4160 4156 4212 4208
rect 1492 3927 1544 3936
rect 1492 3893 1501 3927
rect 1501 3893 1535 3927
rect 1535 3893 1544 3927
rect 1492 3884 1544 3893
rect 3081 3782 3133 3834
rect 3145 3782 3197 3834
rect 3209 3782 3261 3834
rect 3273 3782 3325 3834
rect 3337 3782 3389 3834
rect 7344 3782 7396 3834
rect 7408 3782 7460 3834
rect 7472 3782 7524 3834
rect 7536 3782 7588 3834
rect 7600 3782 7652 3834
rect 11606 3782 11658 3834
rect 11670 3782 11722 3834
rect 11734 3782 11786 3834
rect 11798 3782 11850 3834
rect 11862 3782 11914 3834
rect 5212 3238 5264 3290
rect 5276 3238 5328 3290
rect 5340 3238 5392 3290
rect 5404 3238 5456 3290
rect 5468 3238 5520 3290
rect 9475 3238 9527 3290
rect 9539 3238 9591 3290
rect 9603 3238 9655 3290
rect 9667 3238 9719 3290
rect 9731 3238 9783 3290
rect 13268 2864 13320 2916
rect 3081 2694 3133 2746
rect 3145 2694 3197 2746
rect 3209 2694 3261 2746
rect 3273 2694 3325 2746
rect 3337 2694 3389 2746
rect 7344 2694 7396 2746
rect 7408 2694 7460 2746
rect 7472 2694 7524 2746
rect 7536 2694 7588 2746
rect 7600 2694 7652 2746
rect 11606 2694 11658 2746
rect 11670 2694 11722 2746
rect 11734 2694 11786 2746
rect 11798 2694 11850 2746
rect 11862 2694 11914 2746
rect 5540 2592 5592 2644
rect 4896 2388 4948 2440
rect 8208 2431 8260 2440
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 8208 2388 8260 2397
rect 10784 2388 10836 2440
rect 926 2320 978 2372
rect 2596 2320 2648 2372
rect 2872 2363 2924 2372
rect 2872 2329 2881 2363
rect 2881 2329 2915 2363
rect 2915 2329 2924 2363
rect 2872 2320 2924 2329
rect 5540 2363 5592 2372
rect 5540 2329 5549 2363
rect 5549 2329 5583 2363
rect 5583 2329 5592 2363
rect 5540 2320 5592 2329
rect 7932 2320 7984 2372
rect 10692 2320 10744 2372
rect 13084 2363 13136 2372
rect 13084 2329 13093 2363
rect 13093 2329 13127 2363
rect 13127 2329 13136 2363
rect 13084 2320 13136 2329
rect 5212 2150 5264 2202
rect 5276 2150 5328 2202
rect 5340 2150 5392 2202
rect 5404 2150 5456 2202
rect 5468 2150 5520 2202
rect 9475 2150 9527 2202
rect 9539 2150 9591 2202
rect 9603 2150 9655 2202
rect 9667 2150 9719 2202
rect 9731 2150 9783 2202
<< metal2 >>
rect 1674 16364 1730 17164
rect 4250 16364 4306 17164
rect 7010 16364 7066 17164
rect 9586 16364 9642 17164
rect 12346 16364 12402 17164
rect 14922 16364 14978 17164
rect 1490 15600 1546 15609
rect 1490 15535 1546 15544
rect 1504 14618 1532 15535
rect 1492 14612 1544 14618
rect 1492 14554 1544 14560
rect 1688 14550 1716 16364
rect 3081 14716 3389 14736
rect 3081 14714 3087 14716
rect 3143 14714 3167 14716
rect 3223 14714 3247 14716
rect 3303 14714 3327 14716
rect 3383 14714 3389 14716
rect 3143 14662 3145 14714
rect 3325 14662 3327 14714
rect 3081 14660 3087 14662
rect 3143 14660 3167 14662
rect 3223 14660 3247 14662
rect 3303 14660 3327 14662
rect 3383 14660 3389 14662
rect 3081 14640 3389 14660
rect 4264 14550 4292 16364
rect 7024 14550 7052 16364
rect 7344 14716 7652 14736
rect 7344 14714 7350 14716
rect 7406 14714 7430 14716
rect 7486 14714 7510 14716
rect 7566 14714 7590 14716
rect 7646 14714 7652 14716
rect 7406 14662 7408 14714
rect 7588 14662 7590 14714
rect 7344 14660 7350 14662
rect 7406 14660 7430 14662
rect 7486 14660 7510 14662
rect 7566 14660 7590 14662
rect 7646 14660 7652 14662
rect 7344 14640 7652 14660
rect 1676 14544 1728 14550
rect 1676 14486 1728 14492
rect 4252 14544 4304 14550
rect 4252 14486 4304 14492
rect 7012 14544 7064 14550
rect 7012 14486 7064 14492
rect 9600 14498 9628 16364
rect 11606 14716 11914 14736
rect 11606 14714 11612 14716
rect 11668 14714 11692 14716
rect 11748 14714 11772 14716
rect 11828 14714 11852 14716
rect 11908 14714 11914 14716
rect 11668 14662 11670 14714
rect 11850 14662 11852 14714
rect 11606 14660 11612 14662
rect 11668 14660 11692 14662
rect 11748 14660 11772 14662
rect 11828 14660 11852 14662
rect 11908 14660 11914 14662
rect 11606 14640 11914 14660
rect 12360 14550 12388 16364
rect 12348 14544 12400 14550
rect 9600 14470 9720 14498
rect 12348 14486 12400 14492
rect 9692 14414 9720 14470
rect 14936 14414 14964 16364
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 14924 14408 14976 14414
rect 14924 14350 14976 14356
rect 3081 13628 3389 13648
rect 3081 13626 3087 13628
rect 3143 13626 3167 13628
rect 3223 13626 3247 13628
rect 3303 13626 3327 13628
rect 3383 13626 3389 13628
rect 3143 13574 3145 13626
rect 3325 13574 3327 13626
rect 3081 13572 3087 13574
rect 3143 13572 3167 13574
rect 3223 13572 3247 13574
rect 3303 13572 3327 13574
rect 3383 13572 3389 13574
rect 3081 13552 3389 13572
rect 3081 12540 3389 12560
rect 3081 12538 3087 12540
rect 3143 12538 3167 12540
rect 3223 12538 3247 12540
rect 3303 12538 3327 12540
rect 3383 12538 3389 12540
rect 3143 12486 3145 12538
rect 3325 12486 3327 12538
rect 3081 12484 3087 12486
rect 3143 12484 3167 12486
rect 3223 12484 3247 12486
rect 3303 12484 3327 12486
rect 3383 12484 3389 12486
rect 3081 12464 3389 12484
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1504 11801 1532 12038
rect 1490 11792 1546 11801
rect 1490 11727 1546 11736
rect 3081 11452 3389 11472
rect 3081 11450 3087 11452
rect 3143 11450 3167 11452
rect 3223 11450 3247 11452
rect 3303 11450 3327 11452
rect 3383 11450 3389 11452
rect 3143 11398 3145 11450
rect 3325 11398 3327 11450
rect 3081 11396 3087 11398
rect 3143 11396 3167 11398
rect 3223 11396 3247 11398
rect 3303 11396 3327 11398
rect 3383 11396 3389 11398
rect 3081 11376 3389 11396
rect 3081 10364 3389 10384
rect 3081 10362 3087 10364
rect 3143 10362 3167 10364
rect 3223 10362 3247 10364
rect 3303 10362 3327 10364
rect 3383 10362 3389 10364
rect 3143 10310 3145 10362
rect 3325 10310 3327 10362
rect 3081 10308 3087 10310
rect 3143 10308 3167 10310
rect 3223 10308 3247 10310
rect 3303 10308 3327 10310
rect 3383 10308 3389 10310
rect 3081 10288 3389 10308
rect 3804 10266 3832 14350
rect 4068 14340 4120 14346
rect 4068 14282 4120 14288
rect 6000 14340 6052 14346
rect 6000 14282 6052 14288
rect 4080 10810 4108 14282
rect 5212 14172 5520 14192
rect 5212 14170 5218 14172
rect 5274 14170 5298 14172
rect 5354 14170 5378 14172
rect 5434 14170 5458 14172
rect 5514 14170 5520 14172
rect 5274 14118 5276 14170
rect 5456 14118 5458 14170
rect 5212 14116 5218 14118
rect 5274 14116 5298 14118
rect 5354 14116 5378 14118
rect 5434 14116 5458 14118
rect 5514 14116 5520 14118
rect 5212 14096 5520 14116
rect 5212 13084 5520 13104
rect 5212 13082 5218 13084
rect 5274 13082 5298 13084
rect 5354 13082 5378 13084
rect 5434 13082 5458 13084
rect 5514 13082 5520 13084
rect 5274 13030 5276 13082
rect 5456 13030 5458 13082
rect 5212 13028 5218 13030
rect 5274 13028 5298 13030
rect 5354 13028 5378 13030
rect 5434 13028 5458 13030
rect 5514 13028 5520 13030
rect 5212 13008 5520 13028
rect 4988 12164 5040 12170
rect 4988 12106 5040 12112
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 5000 9654 5028 12106
rect 5212 11996 5520 12016
rect 5212 11994 5218 11996
rect 5274 11994 5298 11996
rect 5354 11994 5378 11996
rect 5434 11994 5458 11996
rect 5514 11994 5520 11996
rect 5274 11942 5276 11994
rect 5456 11942 5458 11994
rect 5212 11940 5218 11942
rect 5274 11940 5298 11942
rect 5354 11940 5378 11942
rect 5434 11940 5458 11942
rect 5514 11940 5520 11942
rect 5212 11920 5520 11940
rect 5212 10908 5520 10928
rect 5212 10906 5218 10908
rect 5274 10906 5298 10908
rect 5354 10906 5378 10908
rect 5434 10906 5458 10908
rect 5514 10906 5520 10908
rect 5274 10854 5276 10906
rect 5456 10854 5458 10906
rect 5212 10852 5218 10854
rect 5274 10852 5298 10854
rect 5354 10852 5378 10854
rect 5434 10852 5458 10854
rect 5514 10852 5520 10854
rect 5212 10832 5520 10852
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5080 10192 5132 10198
rect 5080 10134 5132 10140
rect 5092 9926 5120 10134
rect 5276 9994 5304 10542
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 5092 9722 5120 9862
rect 5212 9820 5520 9840
rect 5212 9818 5218 9820
rect 5274 9818 5298 9820
rect 5354 9818 5378 9820
rect 5434 9818 5458 9820
rect 5514 9818 5520 9820
rect 5274 9766 5276 9818
rect 5456 9766 5458 9818
rect 5212 9764 5218 9766
rect 5274 9764 5298 9766
rect 5354 9764 5378 9766
rect 5434 9764 5458 9766
rect 5514 9764 5520 9766
rect 5212 9744 5520 9764
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 3081 9276 3389 9296
rect 3081 9274 3087 9276
rect 3143 9274 3167 9276
rect 3223 9274 3247 9276
rect 3303 9274 3327 9276
rect 3383 9274 3389 9276
rect 3143 9222 3145 9274
rect 3325 9222 3327 9274
rect 3081 9220 3087 9222
rect 3143 9220 3167 9222
rect 3223 9220 3247 9222
rect 3303 9220 3327 9222
rect 3383 9220 3389 9222
rect 3081 9200 3389 9220
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 3081 8188 3389 8208
rect 3081 8186 3087 8188
rect 3143 8186 3167 8188
rect 3223 8186 3247 8188
rect 3303 8186 3327 8188
rect 3383 8186 3389 8188
rect 3143 8134 3145 8186
rect 3325 8134 3327 8186
rect 3081 8132 3087 8134
rect 3143 8132 3167 8134
rect 3223 8132 3247 8134
rect 3303 8132 3327 8134
rect 3383 8132 3389 8134
rect 3081 8112 3389 8132
rect 5000 7886 5028 8230
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 1492 7744 1544 7750
rect 1490 7712 1492 7721
rect 1544 7712 1546 7721
rect 1490 7647 1546 7656
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 3081 7100 3389 7120
rect 3081 7098 3087 7100
rect 3143 7098 3167 7100
rect 3223 7098 3247 7100
rect 3303 7098 3327 7100
rect 3383 7098 3389 7100
rect 3143 7046 3145 7098
rect 3325 7046 3327 7098
rect 3081 7044 3087 7046
rect 3143 7044 3167 7046
rect 3223 7044 3247 7046
rect 3303 7044 3327 7046
rect 3383 7044 3389 7046
rect 3081 7024 3389 7044
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 1492 3936 1544 3942
rect 1490 3904 1492 3913
rect 1544 3904 1546 3913
rect 1490 3839 1546 3848
rect 2884 2378 2912 6190
rect 3081 6012 3389 6032
rect 3081 6010 3087 6012
rect 3143 6010 3167 6012
rect 3223 6010 3247 6012
rect 3303 6010 3327 6012
rect 3383 6010 3389 6012
rect 3143 5958 3145 6010
rect 3325 5958 3327 6010
rect 3081 5956 3087 5958
rect 3143 5956 3167 5958
rect 3223 5956 3247 5958
rect 3303 5956 3327 5958
rect 3383 5956 3389 5958
rect 3081 5936 3389 5956
rect 3081 4924 3389 4944
rect 3081 4922 3087 4924
rect 3143 4922 3167 4924
rect 3223 4922 3247 4924
rect 3303 4922 3327 4924
rect 3383 4922 3389 4924
rect 3143 4870 3145 4922
rect 3325 4870 3327 4922
rect 3081 4868 3087 4870
rect 3143 4868 3167 4870
rect 3223 4868 3247 4870
rect 3303 4868 3327 4870
rect 3383 4868 3389 4870
rect 3081 4848 3389 4868
rect 4172 4214 4200 7142
rect 5092 6458 5120 9658
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5212 8732 5520 8752
rect 5212 8730 5218 8732
rect 5274 8730 5298 8732
rect 5354 8730 5378 8732
rect 5434 8730 5458 8732
rect 5514 8730 5520 8732
rect 5274 8678 5276 8730
rect 5456 8678 5458 8730
rect 5212 8676 5218 8678
rect 5274 8676 5298 8678
rect 5354 8676 5378 8678
rect 5434 8676 5458 8678
rect 5514 8676 5520 8678
rect 5212 8656 5520 8676
rect 5552 8634 5580 9046
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5212 7644 5520 7664
rect 5212 7642 5218 7644
rect 5274 7642 5298 7644
rect 5354 7642 5378 7644
rect 5434 7642 5458 7644
rect 5514 7642 5520 7644
rect 5274 7590 5276 7642
rect 5456 7590 5458 7642
rect 5212 7588 5218 7590
rect 5274 7588 5298 7590
rect 5354 7588 5378 7590
rect 5434 7588 5458 7590
rect 5514 7588 5520 7590
rect 5212 7568 5520 7588
rect 5552 7274 5580 8570
rect 5644 8022 5672 10610
rect 6012 10266 6040 14282
rect 7208 10810 7236 14350
rect 12256 14340 12308 14346
rect 12256 14282 12308 14288
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9475 14172 9783 14192
rect 9475 14170 9481 14172
rect 9537 14170 9561 14172
rect 9617 14170 9641 14172
rect 9697 14170 9721 14172
rect 9777 14170 9783 14172
rect 9537 14118 9539 14170
rect 9719 14118 9721 14170
rect 9475 14116 9481 14118
rect 9537 14116 9561 14118
rect 9617 14116 9641 14118
rect 9697 14116 9721 14118
rect 9777 14116 9783 14118
rect 9475 14096 9783 14116
rect 7344 13628 7652 13648
rect 7344 13626 7350 13628
rect 7406 13626 7430 13628
rect 7486 13626 7510 13628
rect 7566 13626 7590 13628
rect 7646 13626 7652 13628
rect 7406 13574 7408 13626
rect 7588 13574 7590 13626
rect 7344 13572 7350 13574
rect 7406 13572 7430 13574
rect 7486 13572 7510 13574
rect 7566 13572 7590 13574
rect 7646 13572 7652 13574
rect 7344 13552 7652 13572
rect 9475 13084 9783 13104
rect 9475 13082 9481 13084
rect 9537 13082 9561 13084
rect 9617 13082 9641 13084
rect 9697 13082 9721 13084
rect 9777 13082 9783 13084
rect 9537 13030 9539 13082
rect 9719 13030 9721 13082
rect 9475 13028 9481 13030
rect 9537 13028 9561 13030
rect 9617 13028 9641 13030
rect 9697 13028 9721 13030
rect 9777 13028 9783 13030
rect 9475 13008 9783 13028
rect 7344 12540 7652 12560
rect 7344 12538 7350 12540
rect 7406 12538 7430 12540
rect 7486 12538 7510 12540
rect 7566 12538 7590 12540
rect 7646 12538 7652 12540
rect 7406 12486 7408 12538
rect 7588 12486 7590 12538
rect 7344 12484 7350 12486
rect 7406 12484 7430 12486
rect 7486 12484 7510 12486
rect 7566 12484 7590 12486
rect 7646 12484 7652 12486
rect 7344 12464 7652 12484
rect 9475 11996 9783 12016
rect 9475 11994 9481 11996
rect 9537 11994 9561 11996
rect 9617 11994 9641 11996
rect 9697 11994 9721 11996
rect 9777 11994 9783 11996
rect 9537 11942 9539 11994
rect 9719 11942 9721 11994
rect 9475 11940 9481 11942
rect 9537 11940 9561 11942
rect 9617 11940 9641 11942
rect 9697 11940 9721 11942
rect 9777 11940 9783 11942
rect 9475 11920 9783 11940
rect 7344 11452 7652 11472
rect 7344 11450 7350 11452
rect 7406 11450 7430 11452
rect 7486 11450 7510 11452
rect 7566 11450 7590 11452
rect 7646 11450 7652 11452
rect 7406 11398 7408 11450
rect 7588 11398 7590 11450
rect 7344 11396 7350 11398
rect 7406 11396 7430 11398
rect 7486 11396 7510 11398
rect 7566 11396 7590 11398
rect 7646 11396 7652 11398
rect 7344 11376 7652 11396
rect 9475 10908 9783 10928
rect 9475 10906 9481 10908
rect 9537 10906 9561 10908
rect 9617 10906 9641 10908
rect 9697 10906 9721 10908
rect 9777 10906 9783 10908
rect 9537 10854 9539 10906
rect 9719 10854 9721 10906
rect 9475 10852 9481 10854
rect 9537 10852 9561 10854
rect 9617 10852 9641 10854
rect 9697 10852 9721 10854
rect 9777 10852 9783 10854
rect 9475 10832 9783 10852
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6012 9178 6040 9998
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6564 9450 6592 9930
rect 6552 9444 6604 9450
rect 6552 9386 6604 9392
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5644 7478 5672 7958
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 5908 7472 5960 7478
rect 5908 7414 5960 7420
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5212 6556 5520 6576
rect 5212 6554 5218 6556
rect 5274 6554 5298 6556
rect 5354 6554 5378 6556
rect 5434 6554 5458 6556
rect 5514 6554 5520 6556
rect 5274 6502 5276 6554
rect 5456 6502 5458 6554
rect 5212 6500 5218 6502
rect 5274 6500 5298 6502
rect 5354 6500 5378 6502
rect 5434 6500 5458 6502
rect 5514 6500 5520 6502
rect 5212 6480 5520 6500
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 5368 6066 5396 6258
rect 5552 6186 5580 7210
rect 5920 6458 5948 7414
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 6472 6390 6500 8910
rect 6656 8362 6684 10406
rect 6828 10192 6880 10198
rect 6828 10134 6880 10140
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6748 7886 6776 9862
rect 6840 9586 6868 10134
rect 6932 10130 6960 10746
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 7024 10062 7052 10746
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 7196 10532 7248 10538
rect 7196 10474 7248 10480
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6932 9330 6960 9522
rect 6840 9302 6960 9330
rect 6840 8974 6868 9302
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6920 8900 6972 8906
rect 6920 8842 6972 8848
rect 6932 8498 6960 8842
rect 7024 8514 7052 9998
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7116 8838 7144 9114
rect 7208 8906 7236 10474
rect 7344 10364 7652 10384
rect 7344 10362 7350 10364
rect 7406 10362 7430 10364
rect 7486 10362 7510 10364
rect 7566 10362 7590 10364
rect 7646 10362 7652 10364
rect 7406 10310 7408 10362
rect 7588 10310 7590 10362
rect 7344 10308 7350 10310
rect 7406 10308 7430 10310
rect 7486 10308 7510 10310
rect 7566 10308 7590 10310
rect 7646 10308 7652 10310
rect 7344 10288 7652 10308
rect 7760 9382 7788 10610
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7344 9276 7652 9296
rect 7344 9274 7350 9276
rect 7406 9274 7430 9276
rect 7486 9274 7510 9276
rect 7566 9274 7590 9276
rect 7646 9274 7652 9276
rect 7406 9222 7408 9274
rect 7588 9222 7590 9274
rect 7344 9220 7350 9222
rect 7406 9220 7430 9222
rect 7486 9220 7510 9222
rect 7566 9220 7590 9222
rect 7646 9220 7652 9222
rect 7344 9200 7652 9220
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7760 8566 7788 9318
rect 7748 8560 7800 8566
rect 7024 8498 7144 8514
rect 7748 8502 7800 8508
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7024 8492 7156 8498
rect 7024 8486 7104 8492
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6748 7410 6776 7822
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6748 6914 6776 7346
rect 6748 6886 6868 6914
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 5540 6180 5592 6186
rect 5540 6122 5592 6128
rect 4160 4208 4212 4214
rect 4160 4150 4212 4156
rect 3081 3836 3389 3856
rect 3081 3834 3087 3836
rect 3143 3834 3167 3836
rect 3223 3834 3247 3836
rect 3303 3834 3327 3836
rect 3383 3834 3389 3836
rect 3143 3782 3145 3834
rect 3325 3782 3327 3834
rect 3081 3780 3087 3782
rect 3143 3780 3167 3782
rect 3223 3780 3247 3782
rect 3303 3780 3327 3782
rect 3383 3780 3389 3782
rect 3081 3760 3389 3780
rect 3081 2748 3389 2768
rect 3081 2746 3087 2748
rect 3143 2746 3167 2748
rect 3223 2746 3247 2748
rect 3303 2746 3327 2748
rect 3383 2746 3389 2748
rect 3143 2694 3145 2746
rect 3325 2694 3327 2746
rect 3081 2692 3087 2694
rect 3143 2692 3167 2694
rect 3223 2692 3247 2694
rect 3303 2692 3327 2694
rect 3383 2692 3389 2694
rect 3081 2672 3389 2692
rect 4908 2446 4936 6054
rect 5368 6038 5580 6066
rect 5552 5778 5580 6038
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5212 5468 5520 5488
rect 5212 5466 5218 5468
rect 5274 5466 5298 5468
rect 5354 5466 5378 5468
rect 5434 5466 5458 5468
rect 5514 5466 5520 5468
rect 5274 5414 5276 5466
rect 5456 5414 5458 5466
rect 5212 5412 5218 5414
rect 5274 5412 5298 5414
rect 5354 5412 5378 5414
rect 5434 5412 5458 5414
rect 5514 5412 5520 5414
rect 5212 5392 5520 5412
rect 5212 4380 5520 4400
rect 5212 4378 5218 4380
rect 5274 4378 5298 4380
rect 5354 4378 5378 4380
rect 5434 4378 5458 4380
rect 5514 4378 5520 4380
rect 5274 4326 5276 4378
rect 5456 4326 5458 4378
rect 5212 4324 5218 4326
rect 5274 4324 5298 4326
rect 5354 4324 5378 4326
rect 5434 4324 5458 4326
rect 5514 4324 5520 4326
rect 5212 4304 5520 4324
rect 5212 3292 5520 3312
rect 5212 3290 5218 3292
rect 5274 3290 5298 3292
rect 5354 3290 5378 3292
rect 5434 3290 5458 3292
rect 5514 3290 5520 3292
rect 5274 3238 5276 3290
rect 5456 3238 5458 3290
rect 5212 3236 5218 3238
rect 5274 3236 5298 3238
rect 5354 3236 5378 3238
rect 5434 3236 5458 3238
rect 5514 3236 5520 3238
rect 5212 3216 5520 3236
rect 5552 2650 5580 5714
rect 6472 5574 6500 6326
rect 6840 5778 6868 6886
rect 6932 6322 6960 8434
rect 7024 7546 7052 8486
rect 7104 8434 7156 8440
rect 7344 8188 7652 8208
rect 7344 8186 7350 8188
rect 7406 8186 7430 8188
rect 7486 8186 7510 8188
rect 7566 8186 7590 8188
rect 7646 8186 7652 8188
rect 7406 8134 7408 8186
rect 7588 8134 7590 8186
rect 7344 8132 7350 8134
rect 7406 8132 7430 8134
rect 7486 8132 7510 8134
rect 7566 8132 7590 8134
rect 7646 8132 7652 8134
rect 7344 8112 7652 8132
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7344 7100 7652 7120
rect 7344 7098 7350 7100
rect 7406 7098 7430 7100
rect 7486 7098 7510 7100
rect 7566 7098 7590 7100
rect 7646 7098 7652 7100
rect 7406 7046 7408 7098
rect 7588 7046 7590 7098
rect 7344 7044 7350 7046
rect 7406 7044 7430 7046
rect 7486 7044 7510 7046
rect 7566 7044 7590 7046
rect 7646 7044 7652 7046
rect 7344 7024 7652 7044
rect 7760 6458 7788 8502
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7852 8090 7880 8434
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7944 7562 7972 10542
rect 8128 10266 8156 10610
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 8036 8974 8064 9522
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 7852 7546 7972 7562
rect 7840 7540 7972 7546
rect 7892 7534 7972 7540
rect 7840 7482 7892 7488
rect 8036 7342 8064 8910
rect 8128 7546 8156 10202
rect 8220 9654 8248 10678
rect 8852 10532 8904 10538
rect 8852 10474 8904 10480
rect 8864 9994 8892 10474
rect 9876 10198 9904 14214
rect 11606 13628 11914 13648
rect 11606 13626 11612 13628
rect 11668 13626 11692 13628
rect 11748 13626 11772 13628
rect 11828 13626 11852 13628
rect 11908 13626 11914 13628
rect 11668 13574 11670 13626
rect 11850 13574 11852 13626
rect 11606 13572 11612 13574
rect 11668 13572 11692 13574
rect 11748 13572 11772 13574
rect 11828 13572 11852 13574
rect 11908 13572 11914 13574
rect 11606 13552 11914 13572
rect 11606 12540 11914 12560
rect 11606 12538 11612 12540
rect 11668 12538 11692 12540
rect 11748 12538 11772 12540
rect 11828 12538 11852 12540
rect 11908 12538 11914 12540
rect 11668 12486 11670 12538
rect 11850 12486 11852 12538
rect 11606 12484 11612 12486
rect 11668 12484 11692 12486
rect 11748 12484 11772 12486
rect 11828 12484 11852 12486
rect 11908 12484 11914 12486
rect 11606 12464 11914 12484
rect 11606 11452 11914 11472
rect 11606 11450 11612 11452
rect 11668 11450 11692 11452
rect 11748 11450 11772 11452
rect 11828 11450 11852 11452
rect 11908 11450 11914 11452
rect 11668 11398 11670 11450
rect 11850 11398 11852 11450
rect 11606 11396 11612 11398
rect 11668 11396 11692 11398
rect 11748 11396 11772 11398
rect 11828 11396 11852 11398
rect 11908 11396 11914 11398
rect 11606 11376 11914 11396
rect 12268 10810 12296 14282
rect 13176 13252 13228 13258
rect 13176 13194 13228 13200
rect 13188 13161 13216 13194
rect 13174 13152 13230 13161
rect 13174 13087 13230 13096
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 11606 10364 11914 10384
rect 11606 10362 11612 10364
rect 11668 10362 11692 10364
rect 11748 10362 11772 10364
rect 11828 10362 11852 10364
rect 11908 10362 11914 10364
rect 11668 10310 11670 10362
rect 11850 10310 11852 10362
rect 11606 10308 11612 10310
rect 11668 10308 11692 10310
rect 11748 10308 11772 10310
rect 11828 10308 11852 10310
rect 11908 10308 11914 10310
rect 11606 10288 11914 10308
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 8852 9988 8904 9994
rect 8852 9930 8904 9936
rect 9036 9988 9088 9994
rect 9036 9930 9088 9936
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8220 8498 8248 9590
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8312 8514 8340 9318
rect 8392 9104 8444 9110
rect 8392 9046 8444 9052
rect 8404 8634 8432 9046
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8208 8492 8260 8498
rect 8312 8486 8432 8514
rect 8208 8434 8260 8440
rect 8220 7954 8248 8434
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8312 8022 8340 8298
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 8036 6914 8064 7278
rect 8036 6886 8156 6914
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 7344 6012 7652 6032
rect 7344 6010 7350 6012
rect 7406 6010 7430 6012
rect 7486 6010 7510 6012
rect 7566 6010 7590 6012
rect 7646 6010 7652 6012
rect 7406 5958 7408 6010
rect 7588 5958 7590 6010
rect 7344 5956 7350 5958
rect 7406 5956 7430 5958
rect 7486 5956 7510 5958
rect 7566 5956 7590 5958
rect 7646 5956 7652 5958
rect 7344 5936 7652 5956
rect 8128 5846 8156 6886
rect 8220 6390 8248 7890
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8312 7410 8340 7822
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8312 6866 8340 7346
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 8312 6186 8340 6802
rect 8404 6254 8432 8486
rect 8864 7478 8892 9930
rect 9048 8838 9076 9930
rect 8944 8832 8996 8838
rect 8944 8774 8996 8780
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 8956 8498 8984 8774
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8956 8242 8984 8434
rect 9048 8362 9076 8774
rect 9140 8430 9168 9998
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9232 9110 9260 9862
rect 9475 9820 9783 9840
rect 9475 9818 9481 9820
rect 9537 9818 9561 9820
rect 9617 9818 9641 9820
rect 9697 9818 9721 9820
rect 9777 9818 9783 9820
rect 9537 9766 9539 9818
rect 9719 9766 9721 9818
rect 9475 9764 9481 9766
rect 9537 9764 9561 9766
rect 9617 9764 9641 9766
rect 9697 9764 9721 9766
rect 9777 9764 9783 9766
rect 9475 9744 9783 9764
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 10060 9178 10088 9522
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 13188 9353 13216 9386
rect 13174 9344 13230 9353
rect 11606 9276 11914 9296
rect 13174 9279 13230 9288
rect 11606 9274 11612 9276
rect 11668 9274 11692 9276
rect 11748 9274 11772 9276
rect 11828 9274 11852 9276
rect 11908 9274 11914 9276
rect 11668 9222 11670 9274
rect 11850 9222 11852 9274
rect 11606 9220 11612 9222
rect 11668 9220 11692 9222
rect 11748 9220 11772 9222
rect 11828 9220 11852 9222
rect 11908 9220 11914 9222
rect 11606 9200 11914 9220
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 9220 9104 9272 9110
rect 9220 9046 9272 9052
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9475 8732 9783 8752
rect 9475 8730 9481 8732
rect 9537 8730 9561 8732
rect 9617 8730 9641 8732
rect 9697 8730 9721 8732
rect 9777 8730 9783 8732
rect 9537 8678 9539 8730
rect 9719 8678 9721 8730
rect 9475 8676 9481 8678
rect 9537 8676 9561 8678
rect 9617 8676 9641 8678
rect 9697 8676 9721 8678
rect 9777 8676 9783 8678
rect 9475 8656 9783 8676
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 8956 8214 9076 8242
rect 9048 7478 9076 8214
rect 8852 7472 8904 7478
rect 8852 7414 8904 7420
rect 9036 7472 9088 7478
rect 9036 7414 9088 7420
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8956 6390 8984 7278
rect 9048 6458 9076 7414
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 8944 6384 8996 6390
rect 8944 6326 8996 6332
rect 9140 6322 9168 8366
rect 9475 7644 9783 7664
rect 9475 7642 9481 7644
rect 9537 7642 9561 7644
rect 9617 7642 9641 7644
rect 9697 7642 9721 7644
rect 9777 7642 9783 7644
rect 9537 7590 9539 7642
rect 9719 7590 9721 7642
rect 9475 7588 9481 7590
rect 9537 7588 9561 7590
rect 9617 7588 9641 7590
rect 9697 7588 9721 7590
rect 9777 7588 9783 7590
rect 9475 7568 9783 7588
rect 9968 6866 9996 8774
rect 11606 8188 11914 8208
rect 11606 8186 11612 8188
rect 11668 8186 11692 8188
rect 11748 8186 11772 8188
rect 11828 8186 11852 8188
rect 11908 8186 11914 8188
rect 11668 8134 11670 8186
rect 11850 8134 11852 8186
rect 11606 8132 11612 8134
rect 11668 8132 11692 8134
rect 11748 8132 11772 8134
rect 11828 8132 11852 8134
rect 11908 8132 11914 8134
rect 11606 8112 11914 8132
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 11606 7100 11914 7120
rect 11606 7098 11612 7100
rect 11668 7098 11692 7100
rect 11748 7098 11772 7100
rect 11828 7098 11852 7100
rect 11908 7098 11914 7100
rect 11668 7046 11670 7098
rect 11850 7046 11852 7098
rect 11606 7044 11612 7046
rect 11668 7044 11692 7046
rect 11748 7044 11772 7046
rect 11828 7044 11852 7046
rect 11908 7044 11914 7046
rect 11606 7024 11914 7044
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9475 6556 9783 6576
rect 9475 6554 9481 6556
rect 9537 6554 9561 6556
rect 9617 6554 9641 6556
rect 9697 6554 9721 6556
rect 9777 6554 9783 6556
rect 9537 6502 9539 6554
rect 9719 6502 9721 6554
rect 9475 6500 9481 6502
rect 9537 6500 9561 6502
rect 9617 6500 9641 6502
rect 9697 6500 9721 6502
rect 9777 6500 9783 6502
rect 9475 6480 9783 6500
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 7344 4924 7652 4944
rect 7344 4922 7350 4924
rect 7406 4922 7430 4924
rect 7486 4922 7510 4924
rect 7566 4922 7590 4924
rect 7646 4922 7652 4924
rect 7406 4870 7408 4922
rect 7588 4870 7590 4922
rect 7344 4868 7350 4870
rect 7406 4868 7430 4870
rect 7486 4868 7510 4870
rect 7566 4868 7590 4870
rect 7646 4868 7652 4870
rect 7344 4848 7652 4868
rect 7344 3836 7652 3856
rect 7344 3834 7350 3836
rect 7406 3834 7430 3836
rect 7486 3834 7510 3836
rect 7566 3834 7590 3836
rect 7646 3834 7652 3836
rect 7406 3782 7408 3834
rect 7588 3782 7590 3834
rect 7344 3780 7350 3782
rect 7406 3780 7430 3782
rect 7486 3780 7510 3782
rect 7566 3780 7590 3782
rect 7646 3780 7652 3782
rect 7344 3760 7652 3780
rect 7344 2748 7652 2768
rect 7344 2746 7350 2748
rect 7406 2746 7430 2748
rect 7486 2746 7510 2748
rect 7566 2746 7590 2748
rect 7646 2746 7652 2748
rect 7406 2694 7408 2746
rect 7588 2694 7590 2746
rect 7344 2692 7350 2694
rect 7406 2692 7430 2694
rect 7486 2692 7510 2694
rect 7566 2692 7590 2694
rect 7646 2692 7652 2694
rect 7344 2672 7652 2692
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 8220 2446 8248 6054
rect 9968 5642 9996 6802
rect 11606 6012 11914 6032
rect 11606 6010 11612 6012
rect 11668 6010 11692 6012
rect 11748 6010 11772 6012
rect 11828 6010 11852 6012
rect 11908 6010 11914 6012
rect 11668 5958 11670 6010
rect 11850 5958 11852 6010
rect 11606 5956 11612 5958
rect 11668 5956 11692 5958
rect 11748 5956 11772 5958
rect 11828 5956 11852 5958
rect 11908 5956 11914 5958
rect 11606 5936 11914 5956
rect 13004 5710 13032 7142
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 9956 5636 10008 5642
rect 9956 5578 10008 5584
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 9475 5468 9783 5488
rect 9475 5466 9481 5468
rect 9537 5466 9561 5468
rect 9617 5466 9641 5468
rect 9697 5466 9721 5468
rect 9777 5466 9783 5468
rect 9537 5414 9539 5466
rect 9719 5414 9721 5466
rect 9475 5412 9481 5414
rect 9537 5412 9561 5414
rect 9617 5412 9641 5414
rect 9697 5412 9721 5414
rect 9777 5412 9783 5414
rect 9475 5392 9783 5412
rect 9475 4380 9783 4400
rect 9475 4378 9481 4380
rect 9537 4378 9561 4380
rect 9617 4378 9641 4380
rect 9697 4378 9721 4380
rect 9777 4378 9783 4380
rect 9537 4326 9539 4378
rect 9719 4326 9721 4378
rect 9475 4324 9481 4326
rect 9537 4324 9561 4326
rect 9617 4324 9641 4326
rect 9697 4324 9721 4326
rect 9777 4324 9783 4326
rect 9475 4304 9783 4324
rect 9475 3292 9783 3312
rect 9475 3290 9481 3292
rect 9537 3290 9561 3292
rect 9617 3290 9641 3292
rect 9697 3290 9721 3292
rect 9777 3290 9783 3292
rect 9537 3238 9539 3290
rect 9719 3238 9721 3290
rect 9475 3236 9481 3238
rect 9537 3236 9561 3238
rect 9617 3236 9641 3238
rect 9697 3236 9721 3238
rect 9777 3236 9783 3238
rect 9475 3216 9783 3236
rect 10796 2446 10824 5510
rect 13096 5273 13124 5510
rect 13082 5264 13138 5273
rect 13082 5199 13138 5208
rect 11606 4924 11914 4944
rect 11606 4922 11612 4924
rect 11668 4922 11692 4924
rect 11748 4922 11772 4924
rect 11828 4922 11852 4924
rect 11908 4922 11914 4924
rect 11668 4870 11670 4922
rect 11850 4870 11852 4922
rect 11606 4868 11612 4870
rect 11668 4868 11692 4870
rect 11748 4868 11772 4870
rect 11828 4868 11852 4870
rect 11908 4868 11914 4870
rect 11606 4848 11914 4868
rect 11606 3836 11914 3856
rect 11606 3834 11612 3836
rect 11668 3834 11692 3836
rect 11748 3834 11772 3836
rect 11828 3834 11852 3836
rect 11908 3834 11914 3836
rect 11668 3782 11670 3834
rect 11850 3782 11852 3834
rect 11606 3780 11612 3782
rect 11668 3780 11692 3782
rect 11748 3780 11772 3782
rect 11828 3780 11852 3782
rect 11908 3780 11914 3782
rect 11606 3760 11914 3780
rect 13268 2916 13320 2922
rect 13268 2858 13320 2864
rect 11606 2748 11914 2768
rect 11606 2746 11612 2748
rect 11668 2746 11692 2748
rect 11748 2746 11772 2748
rect 11828 2746 11852 2748
rect 11908 2746 11914 2748
rect 11668 2694 11670 2746
rect 11850 2694 11852 2746
rect 11606 2692 11612 2694
rect 11668 2692 11692 2694
rect 11748 2692 11772 2694
rect 11828 2692 11852 2694
rect 11908 2692 11914 2694
rect 11606 2672 11914 2692
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 926 2372 978 2378
rect 35 2368 926 2372
rect 32 2335 926 2368
rect 32 2295 61 2335
rect 926 2314 978 2320
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 2872 2372 2924 2378
rect 2872 2314 2924 2320
rect 5540 2372 5592 2378
rect 5540 2314 5592 2320
rect 7932 2372 7984 2378
rect 7932 2314 7984 2320
rect 10692 2372 10744 2378
rect 10692 2314 10744 2320
rect 13084 2372 13136 2378
rect 13084 2314 13136 2320
rect 938 2304 966 2314
rect 32 800 60 2295
rect 2608 800 2636 2314
rect 5212 2204 5520 2224
rect 5212 2202 5218 2204
rect 5274 2202 5298 2204
rect 5354 2202 5378 2204
rect 5434 2202 5458 2204
rect 5514 2202 5520 2204
rect 5274 2150 5276 2202
rect 5456 2150 5458 2202
rect 5212 2148 5218 2150
rect 5274 2148 5298 2150
rect 5354 2148 5378 2150
rect 5434 2148 5458 2150
rect 5514 2148 5520 2150
rect 5212 2128 5520 2148
rect 5552 1442 5580 2314
rect 5368 1414 5580 1442
rect 5368 800 5396 1414
rect 7944 800 7972 2314
rect 9475 2204 9783 2224
rect 9475 2202 9481 2204
rect 9537 2202 9561 2204
rect 9617 2202 9641 2204
rect 9697 2202 9721 2204
rect 9777 2202 9783 2204
rect 9537 2150 9539 2202
rect 9719 2150 9721 2202
rect 9475 2148 9481 2150
rect 9537 2148 9561 2150
rect 9617 2148 9641 2150
rect 9697 2148 9721 2150
rect 9777 2148 9783 2150
rect 9475 2128 9783 2148
rect 10704 800 10732 2314
rect 13096 1465 13124 2314
rect 13082 1391 13138 1465
rect 13280 800 13308 2858
rect 18 0 74 800
rect 2594 0 2650 800
rect 5354 0 5410 800
rect 7930 0 7986 800
rect 10690 0 10746 800
rect 13266 0 13322 800
<< via2 >>
rect 1490 15544 1546 15600
rect 3087 14714 3143 14716
rect 3167 14714 3223 14716
rect 3247 14714 3303 14716
rect 3327 14714 3383 14716
rect 3087 14662 3133 14714
rect 3133 14662 3143 14714
rect 3167 14662 3197 14714
rect 3197 14662 3209 14714
rect 3209 14662 3223 14714
rect 3247 14662 3261 14714
rect 3261 14662 3273 14714
rect 3273 14662 3303 14714
rect 3327 14662 3337 14714
rect 3337 14662 3383 14714
rect 3087 14660 3143 14662
rect 3167 14660 3223 14662
rect 3247 14660 3303 14662
rect 3327 14660 3383 14662
rect 7350 14714 7406 14716
rect 7430 14714 7486 14716
rect 7510 14714 7566 14716
rect 7590 14714 7646 14716
rect 7350 14662 7396 14714
rect 7396 14662 7406 14714
rect 7430 14662 7460 14714
rect 7460 14662 7472 14714
rect 7472 14662 7486 14714
rect 7510 14662 7524 14714
rect 7524 14662 7536 14714
rect 7536 14662 7566 14714
rect 7590 14662 7600 14714
rect 7600 14662 7646 14714
rect 7350 14660 7406 14662
rect 7430 14660 7486 14662
rect 7510 14660 7566 14662
rect 7590 14660 7646 14662
rect 11612 14714 11668 14716
rect 11692 14714 11748 14716
rect 11772 14714 11828 14716
rect 11852 14714 11908 14716
rect 11612 14662 11658 14714
rect 11658 14662 11668 14714
rect 11692 14662 11722 14714
rect 11722 14662 11734 14714
rect 11734 14662 11748 14714
rect 11772 14662 11786 14714
rect 11786 14662 11798 14714
rect 11798 14662 11828 14714
rect 11852 14662 11862 14714
rect 11862 14662 11908 14714
rect 11612 14660 11668 14662
rect 11692 14660 11748 14662
rect 11772 14660 11828 14662
rect 11852 14660 11908 14662
rect 3087 13626 3143 13628
rect 3167 13626 3223 13628
rect 3247 13626 3303 13628
rect 3327 13626 3383 13628
rect 3087 13574 3133 13626
rect 3133 13574 3143 13626
rect 3167 13574 3197 13626
rect 3197 13574 3209 13626
rect 3209 13574 3223 13626
rect 3247 13574 3261 13626
rect 3261 13574 3273 13626
rect 3273 13574 3303 13626
rect 3327 13574 3337 13626
rect 3337 13574 3383 13626
rect 3087 13572 3143 13574
rect 3167 13572 3223 13574
rect 3247 13572 3303 13574
rect 3327 13572 3383 13574
rect 3087 12538 3143 12540
rect 3167 12538 3223 12540
rect 3247 12538 3303 12540
rect 3327 12538 3383 12540
rect 3087 12486 3133 12538
rect 3133 12486 3143 12538
rect 3167 12486 3197 12538
rect 3197 12486 3209 12538
rect 3209 12486 3223 12538
rect 3247 12486 3261 12538
rect 3261 12486 3273 12538
rect 3273 12486 3303 12538
rect 3327 12486 3337 12538
rect 3337 12486 3383 12538
rect 3087 12484 3143 12486
rect 3167 12484 3223 12486
rect 3247 12484 3303 12486
rect 3327 12484 3383 12486
rect 1490 11736 1546 11792
rect 3087 11450 3143 11452
rect 3167 11450 3223 11452
rect 3247 11450 3303 11452
rect 3327 11450 3383 11452
rect 3087 11398 3133 11450
rect 3133 11398 3143 11450
rect 3167 11398 3197 11450
rect 3197 11398 3209 11450
rect 3209 11398 3223 11450
rect 3247 11398 3261 11450
rect 3261 11398 3273 11450
rect 3273 11398 3303 11450
rect 3327 11398 3337 11450
rect 3337 11398 3383 11450
rect 3087 11396 3143 11398
rect 3167 11396 3223 11398
rect 3247 11396 3303 11398
rect 3327 11396 3383 11398
rect 3087 10362 3143 10364
rect 3167 10362 3223 10364
rect 3247 10362 3303 10364
rect 3327 10362 3383 10364
rect 3087 10310 3133 10362
rect 3133 10310 3143 10362
rect 3167 10310 3197 10362
rect 3197 10310 3209 10362
rect 3209 10310 3223 10362
rect 3247 10310 3261 10362
rect 3261 10310 3273 10362
rect 3273 10310 3303 10362
rect 3327 10310 3337 10362
rect 3337 10310 3383 10362
rect 3087 10308 3143 10310
rect 3167 10308 3223 10310
rect 3247 10308 3303 10310
rect 3327 10308 3383 10310
rect 5218 14170 5274 14172
rect 5298 14170 5354 14172
rect 5378 14170 5434 14172
rect 5458 14170 5514 14172
rect 5218 14118 5264 14170
rect 5264 14118 5274 14170
rect 5298 14118 5328 14170
rect 5328 14118 5340 14170
rect 5340 14118 5354 14170
rect 5378 14118 5392 14170
rect 5392 14118 5404 14170
rect 5404 14118 5434 14170
rect 5458 14118 5468 14170
rect 5468 14118 5514 14170
rect 5218 14116 5274 14118
rect 5298 14116 5354 14118
rect 5378 14116 5434 14118
rect 5458 14116 5514 14118
rect 5218 13082 5274 13084
rect 5298 13082 5354 13084
rect 5378 13082 5434 13084
rect 5458 13082 5514 13084
rect 5218 13030 5264 13082
rect 5264 13030 5274 13082
rect 5298 13030 5328 13082
rect 5328 13030 5340 13082
rect 5340 13030 5354 13082
rect 5378 13030 5392 13082
rect 5392 13030 5404 13082
rect 5404 13030 5434 13082
rect 5458 13030 5468 13082
rect 5468 13030 5514 13082
rect 5218 13028 5274 13030
rect 5298 13028 5354 13030
rect 5378 13028 5434 13030
rect 5458 13028 5514 13030
rect 5218 11994 5274 11996
rect 5298 11994 5354 11996
rect 5378 11994 5434 11996
rect 5458 11994 5514 11996
rect 5218 11942 5264 11994
rect 5264 11942 5274 11994
rect 5298 11942 5328 11994
rect 5328 11942 5340 11994
rect 5340 11942 5354 11994
rect 5378 11942 5392 11994
rect 5392 11942 5404 11994
rect 5404 11942 5434 11994
rect 5458 11942 5468 11994
rect 5468 11942 5514 11994
rect 5218 11940 5274 11942
rect 5298 11940 5354 11942
rect 5378 11940 5434 11942
rect 5458 11940 5514 11942
rect 5218 10906 5274 10908
rect 5298 10906 5354 10908
rect 5378 10906 5434 10908
rect 5458 10906 5514 10908
rect 5218 10854 5264 10906
rect 5264 10854 5274 10906
rect 5298 10854 5328 10906
rect 5328 10854 5340 10906
rect 5340 10854 5354 10906
rect 5378 10854 5392 10906
rect 5392 10854 5404 10906
rect 5404 10854 5434 10906
rect 5458 10854 5468 10906
rect 5468 10854 5514 10906
rect 5218 10852 5274 10854
rect 5298 10852 5354 10854
rect 5378 10852 5434 10854
rect 5458 10852 5514 10854
rect 5218 9818 5274 9820
rect 5298 9818 5354 9820
rect 5378 9818 5434 9820
rect 5458 9818 5514 9820
rect 5218 9766 5264 9818
rect 5264 9766 5274 9818
rect 5298 9766 5328 9818
rect 5328 9766 5340 9818
rect 5340 9766 5354 9818
rect 5378 9766 5392 9818
rect 5392 9766 5404 9818
rect 5404 9766 5434 9818
rect 5458 9766 5468 9818
rect 5468 9766 5514 9818
rect 5218 9764 5274 9766
rect 5298 9764 5354 9766
rect 5378 9764 5434 9766
rect 5458 9764 5514 9766
rect 3087 9274 3143 9276
rect 3167 9274 3223 9276
rect 3247 9274 3303 9276
rect 3327 9274 3383 9276
rect 3087 9222 3133 9274
rect 3133 9222 3143 9274
rect 3167 9222 3197 9274
rect 3197 9222 3209 9274
rect 3209 9222 3223 9274
rect 3247 9222 3261 9274
rect 3261 9222 3273 9274
rect 3273 9222 3303 9274
rect 3327 9222 3337 9274
rect 3337 9222 3383 9274
rect 3087 9220 3143 9222
rect 3167 9220 3223 9222
rect 3247 9220 3303 9222
rect 3327 9220 3383 9222
rect 3087 8186 3143 8188
rect 3167 8186 3223 8188
rect 3247 8186 3303 8188
rect 3327 8186 3383 8188
rect 3087 8134 3133 8186
rect 3133 8134 3143 8186
rect 3167 8134 3197 8186
rect 3197 8134 3209 8186
rect 3209 8134 3223 8186
rect 3247 8134 3261 8186
rect 3261 8134 3273 8186
rect 3273 8134 3303 8186
rect 3327 8134 3337 8186
rect 3337 8134 3383 8186
rect 3087 8132 3143 8134
rect 3167 8132 3223 8134
rect 3247 8132 3303 8134
rect 3327 8132 3383 8134
rect 1490 7692 1492 7712
rect 1492 7692 1544 7712
rect 1544 7692 1546 7712
rect 1490 7656 1546 7692
rect 3087 7098 3143 7100
rect 3167 7098 3223 7100
rect 3247 7098 3303 7100
rect 3327 7098 3383 7100
rect 3087 7046 3133 7098
rect 3133 7046 3143 7098
rect 3167 7046 3197 7098
rect 3197 7046 3209 7098
rect 3209 7046 3223 7098
rect 3247 7046 3261 7098
rect 3261 7046 3273 7098
rect 3273 7046 3303 7098
rect 3327 7046 3337 7098
rect 3337 7046 3383 7098
rect 3087 7044 3143 7046
rect 3167 7044 3223 7046
rect 3247 7044 3303 7046
rect 3327 7044 3383 7046
rect 1490 3884 1492 3904
rect 1492 3884 1544 3904
rect 1544 3884 1546 3904
rect 1490 3848 1546 3884
rect 3087 6010 3143 6012
rect 3167 6010 3223 6012
rect 3247 6010 3303 6012
rect 3327 6010 3383 6012
rect 3087 5958 3133 6010
rect 3133 5958 3143 6010
rect 3167 5958 3197 6010
rect 3197 5958 3209 6010
rect 3209 5958 3223 6010
rect 3247 5958 3261 6010
rect 3261 5958 3273 6010
rect 3273 5958 3303 6010
rect 3327 5958 3337 6010
rect 3337 5958 3383 6010
rect 3087 5956 3143 5958
rect 3167 5956 3223 5958
rect 3247 5956 3303 5958
rect 3327 5956 3383 5958
rect 3087 4922 3143 4924
rect 3167 4922 3223 4924
rect 3247 4922 3303 4924
rect 3327 4922 3383 4924
rect 3087 4870 3133 4922
rect 3133 4870 3143 4922
rect 3167 4870 3197 4922
rect 3197 4870 3209 4922
rect 3209 4870 3223 4922
rect 3247 4870 3261 4922
rect 3261 4870 3273 4922
rect 3273 4870 3303 4922
rect 3327 4870 3337 4922
rect 3337 4870 3383 4922
rect 3087 4868 3143 4870
rect 3167 4868 3223 4870
rect 3247 4868 3303 4870
rect 3327 4868 3383 4870
rect 5218 8730 5274 8732
rect 5298 8730 5354 8732
rect 5378 8730 5434 8732
rect 5458 8730 5514 8732
rect 5218 8678 5264 8730
rect 5264 8678 5274 8730
rect 5298 8678 5328 8730
rect 5328 8678 5340 8730
rect 5340 8678 5354 8730
rect 5378 8678 5392 8730
rect 5392 8678 5404 8730
rect 5404 8678 5434 8730
rect 5458 8678 5468 8730
rect 5468 8678 5514 8730
rect 5218 8676 5274 8678
rect 5298 8676 5354 8678
rect 5378 8676 5434 8678
rect 5458 8676 5514 8678
rect 5218 7642 5274 7644
rect 5298 7642 5354 7644
rect 5378 7642 5434 7644
rect 5458 7642 5514 7644
rect 5218 7590 5264 7642
rect 5264 7590 5274 7642
rect 5298 7590 5328 7642
rect 5328 7590 5340 7642
rect 5340 7590 5354 7642
rect 5378 7590 5392 7642
rect 5392 7590 5404 7642
rect 5404 7590 5434 7642
rect 5458 7590 5468 7642
rect 5468 7590 5514 7642
rect 5218 7588 5274 7590
rect 5298 7588 5354 7590
rect 5378 7588 5434 7590
rect 5458 7588 5514 7590
rect 9481 14170 9537 14172
rect 9561 14170 9617 14172
rect 9641 14170 9697 14172
rect 9721 14170 9777 14172
rect 9481 14118 9527 14170
rect 9527 14118 9537 14170
rect 9561 14118 9591 14170
rect 9591 14118 9603 14170
rect 9603 14118 9617 14170
rect 9641 14118 9655 14170
rect 9655 14118 9667 14170
rect 9667 14118 9697 14170
rect 9721 14118 9731 14170
rect 9731 14118 9777 14170
rect 9481 14116 9537 14118
rect 9561 14116 9617 14118
rect 9641 14116 9697 14118
rect 9721 14116 9777 14118
rect 7350 13626 7406 13628
rect 7430 13626 7486 13628
rect 7510 13626 7566 13628
rect 7590 13626 7646 13628
rect 7350 13574 7396 13626
rect 7396 13574 7406 13626
rect 7430 13574 7460 13626
rect 7460 13574 7472 13626
rect 7472 13574 7486 13626
rect 7510 13574 7524 13626
rect 7524 13574 7536 13626
rect 7536 13574 7566 13626
rect 7590 13574 7600 13626
rect 7600 13574 7646 13626
rect 7350 13572 7406 13574
rect 7430 13572 7486 13574
rect 7510 13572 7566 13574
rect 7590 13572 7646 13574
rect 9481 13082 9537 13084
rect 9561 13082 9617 13084
rect 9641 13082 9697 13084
rect 9721 13082 9777 13084
rect 9481 13030 9527 13082
rect 9527 13030 9537 13082
rect 9561 13030 9591 13082
rect 9591 13030 9603 13082
rect 9603 13030 9617 13082
rect 9641 13030 9655 13082
rect 9655 13030 9667 13082
rect 9667 13030 9697 13082
rect 9721 13030 9731 13082
rect 9731 13030 9777 13082
rect 9481 13028 9537 13030
rect 9561 13028 9617 13030
rect 9641 13028 9697 13030
rect 9721 13028 9777 13030
rect 7350 12538 7406 12540
rect 7430 12538 7486 12540
rect 7510 12538 7566 12540
rect 7590 12538 7646 12540
rect 7350 12486 7396 12538
rect 7396 12486 7406 12538
rect 7430 12486 7460 12538
rect 7460 12486 7472 12538
rect 7472 12486 7486 12538
rect 7510 12486 7524 12538
rect 7524 12486 7536 12538
rect 7536 12486 7566 12538
rect 7590 12486 7600 12538
rect 7600 12486 7646 12538
rect 7350 12484 7406 12486
rect 7430 12484 7486 12486
rect 7510 12484 7566 12486
rect 7590 12484 7646 12486
rect 9481 11994 9537 11996
rect 9561 11994 9617 11996
rect 9641 11994 9697 11996
rect 9721 11994 9777 11996
rect 9481 11942 9527 11994
rect 9527 11942 9537 11994
rect 9561 11942 9591 11994
rect 9591 11942 9603 11994
rect 9603 11942 9617 11994
rect 9641 11942 9655 11994
rect 9655 11942 9667 11994
rect 9667 11942 9697 11994
rect 9721 11942 9731 11994
rect 9731 11942 9777 11994
rect 9481 11940 9537 11942
rect 9561 11940 9617 11942
rect 9641 11940 9697 11942
rect 9721 11940 9777 11942
rect 7350 11450 7406 11452
rect 7430 11450 7486 11452
rect 7510 11450 7566 11452
rect 7590 11450 7646 11452
rect 7350 11398 7396 11450
rect 7396 11398 7406 11450
rect 7430 11398 7460 11450
rect 7460 11398 7472 11450
rect 7472 11398 7486 11450
rect 7510 11398 7524 11450
rect 7524 11398 7536 11450
rect 7536 11398 7566 11450
rect 7590 11398 7600 11450
rect 7600 11398 7646 11450
rect 7350 11396 7406 11398
rect 7430 11396 7486 11398
rect 7510 11396 7566 11398
rect 7590 11396 7646 11398
rect 9481 10906 9537 10908
rect 9561 10906 9617 10908
rect 9641 10906 9697 10908
rect 9721 10906 9777 10908
rect 9481 10854 9527 10906
rect 9527 10854 9537 10906
rect 9561 10854 9591 10906
rect 9591 10854 9603 10906
rect 9603 10854 9617 10906
rect 9641 10854 9655 10906
rect 9655 10854 9667 10906
rect 9667 10854 9697 10906
rect 9721 10854 9731 10906
rect 9731 10854 9777 10906
rect 9481 10852 9537 10854
rect 9561 10852 9617 10854
rect 9641 10852 9697 10854
rect 9721 10852 9777 10854
rect 5218 6554 5274 6556
rect 5298 6554 5354 6556
rect 5378 6554 5434 6556
rect 5458 6554 5514 6556
rect 5218 6502 5264 6554
rect 5264 6502 5274 6554
rect 5298 6502 5328 6554
rect 5328 6502 5340 6554
rect 5340 6502 5354 6554
rect 5378 6502 5392 6554
rect 5392 6502 5404 6554
rect 5404 6502 5434 6554
rect 5458 6502 5468 6554
rect 5468 6502 5514 6554
rect 5218 6500 5274 6502
rect 5298 6500 5354 6502
rect 5378 6500 5434 6502
rect 5458 6500 5514 6502
rect 7350 10362 7406 10364
rect 7430 10362 7486 10364
rect 7510 10362 7566 10364
rect 7590 10362 7646 10364
rect 7350 10310 7396 10362
rect 7396 10310 7406 10362
rect 7430 10310 7460 10362
rect 7460 10310 7472 10362
rect 7472 10310 7486 10362
rect 7510 10310 7524 10362
rect 7524 10310 7536 10362
rect 7536 10310 7566 10362
rect 7590 10310 7600 10362
rect 7600 10310 7646 10362
rect 7350 10308 7406 10310
rect 7430 10308 7486 10310
rect 7510 10308 7566 10310
rect 7590 10308 7646 10310
rect 7350 9274 7406 9276
rect 7430 9274 7486 9276
rect 7510 9274 7566 9276
rect 7590 9274 7646 9276
rect 7350 9222 7396 9274
rect 7396 9222 7406 9274
rect 7430 9222 7460 9274
rect 7460 9222 7472 9274
rect 7472 9222 7486 9274
rect 7510 9222 7524 9274
rect 7524 9222 7536 9274
rect 7536 9222 7566 9274
rect 7590 9222 7600 9274
rect 7600 9222 7646 9274
rect 7350 9220 7406 9222
rect 7430 9220 7486 9222
rect 7510 9220 7566 9222
rect 7590 9220 7646 9222
rect 3087 3834 3143 3836
rect 3167 3834 3223 3836
rect 3247 3834 3303 3836
rect 3327 3834 3383 3836
rect 3087 3782 3133 3834
rect 3133 3782 3143 3834
rect 3167 3782 3197 3834
rect 3197 3782 3209 3834
rect 3209 3782 3223 3834
rect 3247 3782 3261 3834
rect 3261 3782 3273 3834
rect 3273 3782 3303 3834
rect 3327 3782 3337 3834
rect 3337 3782 3383 3834
rect 3087 3780 3143 3782
rect 3167 3780 3223 3782
rect 3247 3780 3303 3782
rect 3327 3780 3383 3782
rect 3087 2746 3143 2748
rect 3167 2746 3223 2748
rect 3247 2746 3303 2748
rect 3327 2746 3383 2748
rect 3087 2694 3133 2746
rect 3133 2694 3143 2746
rect 3167 2694 3197 2746
rect 3197 2694 3209 2746
rect 3209 2694 3223 2746
rect 3247 2694 3261 2746
rect 3261 2694 3273 2746
rect 3273 2694 3303 2746
rect 3327 2694 3337 2746
rect 3337 2694 3383 2746
rect 3087 2692 3143 2694
rect 3167 2692 3223 2694
rect 3247 2692 3303 2694
rect 3327 2692 3383 2694
rect 5218 5466 5274 5468
rect 5298 5466 5354 5468
rect 5378 5466 5434 5468
rect 5458 5466 5514 5468
rect 5218 5414 5264 5466
rect 5264 5414 5274 5466
rect 5298 5414 5328 5466
rect 5328 5414 5340 5466
rect 5340 5414 5354 5466
rect 5378 5414 5392 5466
rect 5392 5414 5404 5466
rect 5404 5414 5434 5466
rect 5458 5414 5468 5466
rect 5468 5414 5514 5466
rect 5218 5412 5274 5414
rect 5298 5412 5354 5414
rect 5378 5412 5434 5414
rect 5458 5412 5514 5414
rect 5218 4378 5274 4380
rect 5298 4378 5354 4380
rect 5378 4378 5434 4380
rect 5458 4378 5514 4380
rect 5218 4326 5264 4378
rect 5264 4326 5274 4378
rect 5298 4326 5328 4378
rect 5328 4326 5340 4378
rect 5340 4326 5354 4378
rect 5378 4326 5392 4378
rect 5392 4326 5404 4378
rect 5404 4326 5434 4378
rect 5458 4326 5468 4378
rect 5468 4326 5514 4378
rect 5218 4324 5274 4326
rect 5298 4324 5354 4326
rect 5378 4324 5434 4326
rect 5458 4324 5514 4326
rect 5218 3290 5274 3292
rect 5298 3290 5354 3292
rect 5378 3290 5434 3292
rect 5458 3290 5514 3292
rect 5218 3238 5264 3290
rect 5264 3238 5274 3290
rect 5298 3238 5328 3290
rect 5328 3238 5340 3290
rect 5340 3238 5354 3290
rect 5378 3238 5392 3290
rect 5392 3238 5404 3290
rect 5404 3238 5434 3290
rect 5458 3238 5468 3290
rect 5468 3238 5514 3290
rect 5218 3236 5274 3238
rect 5298 3236 5354 3238
rect 5378 3236 5434 3238
rect 5458 3236 5514 3238
rect 7350 8186 7406 8188
rect 7430 8186 7486 8188
rect 7510 8186 7566 8188
rect 7590 8186 7646 8188
rect 7350 8134 7396 8186
rect 7396 8134 7406 8186
rect 7430 8134 7460 8186
rect 7460 8134 7472 8186
rect 7472 8134 7486 8186
rect 7510 8134 7524 8186
rect 7524 8134 7536 8186
rect 7536 8134 7566 8186
rect 7590 8134 7600 8186
rect 7600 8134 7646 8186
rect 7350 8132 7406 8134
rect 7430 8132 7486 8134
rect 7510 8132 7566 8134
rect 7590 8132 7646 8134
rect 7350 7098 7406 7100
rect 7430 7098 7486 7100
rect 7510 7098 7566 7100
rect 7590 7098 7646 7100
rect 7350 7046 7396 7098
rect 7396 7046 7406 7098
rect 7430 7046 7460 7098
rect 7460 7046 7472 7098
rect 7472 7046 7486 7098
rect 7510 7046 7524 7098
rect 7524 7046 7536 7098
rect 7536 7046 7566 7098
rect 7590 7046 7600 7098
rect 7600 7046 7646 7098
rect 7350 7044 7406 7046
rect 7430 7044 7486 7046
rect 7510 7044 7566 7046
rect 7590 7044 7646 7046
rect 11612 13626 11668 13628
rect 11692 13626 11748 13628
rect 11772 13626 11828 13628
rect 11852 13626 11908 13628
rect 11612 13574 11658 13626
rect 11658 13574 11668 13626
rect 11692 13574 11722 13626
rect 11722 13574 11734 13626
rect 11734 13574 11748 13626
rect 11772 13574 11786 13626
rect 11786 13574 11798 13626
rect 11798 13574 11828 13626
rect 11852 13574 11862 13626
rect 11862 13574 11908 13626
rect 11612 13572 11668 13574
rect 11692 13572 11748 13574
rect 11772 13572 11828 13574
rect 11852 13572 11908 13574
rect 11612 12538 11668 12540
rect 11692 12538 11748 12540
rect 11772 12538 11828 12540
rect 11852 12538 11908 12540
rect 11612 12486 11658 12538
rect 11658 12486 11668 12538
rect 11692 12486 11722 12538
rect 11722 12486 11734 12538
rect 11734 12486 11748 12538
rect 11772 12486 11786 12538
rect 11786 12486 11798 12538
rect 11798 12486 11828 12538
rect 11852 12486 11862 12538
rect 11862 12486 11908 12538
rect 11612 12484 11668 12486
rect 11692 12484 11748 12486
rect 11772 12484 11828 12486
rect 11852 12484 11908 12486
rect 11612 11450 11668 11452
rect 11692 11450 11748 11452
rect 11772 11450 11828 11452
rect 11852 11450 11908 11452
rect 11612 11398 11658 11450
rect 11658 11398 11668 11450
rect 11692 11398 11722 11450
rect 11722 11398 11734 11450
rect 11734 11398 11748 11450
rect 11772 11398 11786 11450
rect 11786 11398 11798 11450
rect 11798 11398 11828 11450
rect 11852 11398 11862 11450
rect 11862 11398 11908 11450
rect 11612 11396 11668 11398
rect 11692 11396 11748 11398
rect 11772 11396 11828 11398
rect 11852 11396 11908 11398
rect 13174 13096 13230 13152
rect 11612 10362 11668 10364
rect 11692 10362 11748 10364
rect 11772 10362 11828 10364
rect 11852 10362 11908 10364
rect 11612 10310 11658 10362
rect 11658 10310 11668 10362
rect 11692 10310 11722 10362
rect 11722 10310 11734 10362
rect 11734 10310 11748 10362
rect 11772 10310 11786 10362
rect 11786 10310 11798 10362
rect 11798 10310 11828 10362
rect 11852 10310 11862 10362
rect 11862 10310 11908 10362
rect 11612 10308 11668 10310
rect 11692 10308 11748 10310
rect 11772 10308 11828 10310
rect 11852 10308 11908 10310
rect 7350 6010 7406 6012
rect 7430 6010 7486 6012
rect 7510 6010 7566 6012
rect 7590 6010 7646 6012
rect 7350 5958 7396 6010
rect 7396 5958 7406 6010
rect 7430 5958 7460 6010
rect 7460 5958 7472 6010
rect 7472 5958 7486 6010
rect 7510 5958 7524 6010
rect 7524 5958 7536 6010
rect 7536 5958 7566 6010
rect 7590 5958 7600 6010
rect 7600 5958 7646 6010
rect 7350 5956 7406 5958
rect 7430 5956 7486 5958
rect 7510 5956 7566 5958
rect 7590 5956 7646 5958
rect 9481 9818 9537 9820
rect 9561 9818 9617 9820
rect 9641 9818 9697 9820
rect 9721 9818 9777 9820
rect 9481 9766 9527 9818
rect 9527 9766 9537 9818
rect 9561 9766 9591 9818
rect 9591 9766 9603 9818
rect 9603 9766 9617 9818
rect 9641 9766 9655 9818
rect 9655 9766 9667 9818
rect 9667 9766 9697 9818
rect 9721 9766 9731 9818
rect 9731 9766 9777 9818
rect 9481 9764 9537 9766
rect 9561 9764 9617 9766
rect 9641 9764 9697 9766
rect 9721 9764 9777 9766
rect 13174 9288 13230 9344
rect 11612 9274 11668 9276
rect 11692 9274 11748 9276
rect 11772 9274 11828 9276
rect 11852 9274 11908 9276
rect 11612 9222 11658 9274
rect 11658 9222 11668 9274
rect 11692 9222 11722 9274
rect 11722 9222 11734 9274
rect 11734 9222 11748 9274
rect 11772 9222 11786 9274
rect 11786 9222 11798 9274
rect 11798 9222 11828 9274
rect 11852 9222 11862 9274
rect 11862 9222 11908 9274
rect 11612 9220 11668 9222
rect 11692 9220 11748 9222
rect 11772 9220 11828 9222
rect 11852 9220 11908 9222
rect 9481 8730 9537 8732
rect 9561 8730 9617 8732
rect 9641 8730 9697 8732
rect 9721 8730 9777 8732
rect 9481 8678 9527 8730
rect 9527 8678 9537 8730
rect 9561 8678 9591 8730
rect 9591 8678 9603 8730
rect 9603 8678 9617 8730
rect 9641 8678 9655 8730
rect 9655 8678 9667 8730
rect 9667 8678 9697 8730
rect 9721 8678 9731 8730
rect 9731 8678 9777 8730
rect 9481 8676 9537 8678
rect 9561 8676 9617 8678
rect 9641 8676 9697 8678
rect 9721 8676 9777 8678
rect 9481 7642 9537 7644
rect 9561 7642 9617 7644
rect 9641 7642 9697 7644
rect 9721 7642 9777 7644
rect 9481 7590 9527 7642
rect 9527 7590 9537 7642
rect 9561 7590 9591 7642
rect 9591 7590 9603 7642
rect 9603 7590 9617 7642
rect 9641 7590 9655 7642
rect 9655 7590 9667 7642
rect 9667 7590 9697 7642
rect 9721 7590 9731 7642
rect 9731 7590 9777 7642
rect 9481 7588 9537 7590
rect 9561 7588 9617 7590
rect 9641 7588 9697 7590
rect 9721 7588 9777 7590
rect 11612 8186 11668 8188
rect 11692 8186 11748 8188
rect 11772 8186 11828 8188
rect 11852 8186 11908 8188
rect 11612 8134 11658 8186
rect 11658 8134 11668 8186
rect 11692 8134 11722 8186
rect 11722 8134 11734 8186
rect 11734 8134 11748 8186
rect 11772 8134 11786 8186
rect 11786 8134 11798 8186
rect 11798 8134 11828 8186
rect 11852 8134 11862 8186
rect 11862 8134 11908 8186
rect 11612 8132 11668 8134
rect 11692 8132 11748 8134
rect 11772 8132 11828 8134
rect 11852 8132 11908 8134
rect 11612 7098 11668 7100
rect 11692 7098 11748 7100
rect 11772 7098 11828 7100
rect 11852 7098 11908 7100
rect 11612 7046 11658 7098
rect 11658 7046 11668 7098
rect 11692 7046 11722 7098
rect 11722 7046 11734 7098
rect 11734 7046 11748 7098
rect 11772 7046 11786 7098
rect 11786 7046 11798 7098
rect 11798 7046 11828 7098
rect 11852 7046 11862 7098
rect 11862 7046 11908 7098
rect 11612 7044 11668 7046
rect 11692 7044 11748 7046
rect 11772 7044 11828 7046
rect 11852 7044 11908 7046
rect 9481 6554 9537 6556
rect 9561 6554 9617 6556
rect 9641 6554 9697 6556
rect 9721 6554 9777 6556
rect 9481 6502 9527 6554
rect 9527 6502 9537 6554
rect 9561 6502 9591 6554
rect 9591 6502 9603 6554
rect 9603 6502 9617 6554
rect 9641 6502 9655 6554
rect 9655 6502 9667 6554
rect 9667 6502 9697 6554
rect 9721 6502 9731 6554
rect 9731 6502 9777 6554
rect 9481 6500 9537 6502
rect 9561 6500 9617 6502
rect 9641 6500 9697 6502
rect 9721 6500 9777 6502
rect 7350 4922 7406 4924
rect 7430 4922 7486 4924
rect 7510 4922 7566 4924
rect 7590 4922 7646 4924
rect 7350 4870 7396 4922
rect 7396 4870 7406 4922
rect 7430 4870 7460 4922
rect 7460 4870 7472 4922
rect 7472 4870 7486 4922
rect 7510 4870 7524 4922
rect 7524 4870 7536 4922
rect 7536 4870 7566 4922
rect 7590 4870 7600 4922
rect 7600 4870 7646 4922
rect 7350 4868 7406 4870
rect 7430 4868 7486 4870
rect 7510 4868 7566 4870
rect 7590 4868 7646 4870
rect 7350 3834 7406 3836
rect 7430 3834 7486 3836
rect 7510 3834 7566 3836
rect 7590 3834 7646 3836
rect 7350 3782 7396 3834
rect 7396 3782 7406 3834
rect 7430 3782 7460 3834
rect 7460 3782 7472 3834
rect 7472 3782 7486 3834
rect 7510 3782 7524 3834
rect 7524 3782 7536 3834
rect 7536 3782 7566 3834
rect 7590 3782 7600 3834
rect 7600 3782 7646 3834
rect 7350 3780 7406 3782
rect 7430 3780 7486 3782
rect 7510 3780 7566 3782
rect 7590 3780 7646 3782
rect 7350 2746 7406 2748
rect 7430 2746 7486 2748
rect 7510 2746 7566 2748
rect 7590 2746 7646 2748
rect 7350 2694 7396 2746
rect 7396 2694 7406 2746
rect 7430 2694 7460 2746
rect 7460 2694 7472 2746
rect 7472 2694 7486 2746
rect 7510 2694 7524 2746
rect 7524 2694 7536 2746
rect 7536 2694 7566 2746
rect 7590 2694 7600 2746
rect 7600 2694 7646 2746
rect 7350 2692 7406 2694
rect 7430 2692 7486 2694
rect 7510 2692 7566 2694
rect 7590 2692 7646 2694
rect 11612 6010 11668 6012
rect 11692 6010 11748 6012
rect 11772 6010 11828 6012
rect 11852 6010 11908 6012
rect 11612 5958 11658 6010
rect 11658 5958 11668 6010
rect 11692 5958 11722 6010
rect 11722 5958 11734 6010
rect 11734 5958 11748 6010
rect 11772 5958 11786 6010
rect 11786 5958 11798 6010
rect 11798 5958 11828 6010
rect 11852 5958 11862 6010
rect 11862 5958 11908 6010
rect 11612 5956 11668 5958
rect 11692 5956 11748 5958
rect 11772 5956 11828 5958
rect 11852 5956 11908 5958
rect 9481 5466 9537 5468
rect 9561 5466 9617 5468
rect 9641 5466 9697 5468
rect 9721 5466 9777 5468
rect 9481 5414 9527 5466
rect 9527 5414 9537 5466
rect 9561 5414 9591 5466
rect 9591 5414 9603 5466
rect 9603 5414 9617 5466
rect 9641 5414 9655 5466
rect 9655 5414 9667 5466
rect 9667 5414 9697 5466
rect 9721 5414 9731 5466
rect 9731 5414 9777 5466
rect 9481 5412 9537 5414
rect 9561 5412 9617 5414
rect 9641 5412 9697 5414
rect 9721 5412 9777 5414
rect 9481 4378 9537 4380
rect 9561 4378 9617 4380
rect 9641 4378 9697 4380
rect 9721 4378 9777 4380
rect 9481 4326 9527 4378
rect 9527 4326 9537 4378
rect 9561 4326 9591 4378
rect 9591 4326 9603 4378
rect 9603 4326 9617 4378
rect 9641 4326 9655 4378
rect 9655 4326 9667 4378
rect 9667 4326 9697 4378
rect 9721 4326 9731 4378
rect 9731 4326 9777 4378
rect 9481 4324 9537 4326
rect 9561 4324 9617 4326
rect 9641 4324 9697 4326
rect 9721 4324 9777 4326
rect 9481 3290 9537 3292
rect 9561 3290 9617 3292
rect 9641 3290 9697 3292
rect 9721 3290 9777 3292
rect 9481 3238 9527 3290
rect 9527 3238 9537 3290
rect 9561 3238 9591 3290
rect 9591 3238 9603 3290
rect 9603 3238 9617 3290
rect 9641 3238 9655 3290
rect 9655 3238 9667 3290
rect 9667 3238 9697 3290
rect 9721 3238 9731 3290
rect 9731 3238 9777 3290
rect 9481 3236 9537 3238
rect 9561 3236 9617 3238
rect 9641 3236 9697 3238
rect 9721 3236 9777 3238
rect 13082 5208 13138 5264
rect 11612 4922 11668 4924
rect 11692 4922 11748 4924
rect 11772 4922 11828 4924
rect 11852 4922 11908 4924
rect 11612 4870 11658 4922
rect 11658 4870 11668 4922
rect 11692 4870 11722 4922
rect 11722 4870 11734 4922
rect 11734 4870 11748 4922
rect 11772 4870 11786 4922
rect 11786 4870 11798 4922
rect 11798 4870 11828 4922
rect 11852 4870 11862 4922
rect 11862 4870 11908 4922
rect 11612 4868 11668 4870
rect 11692 4868 11748 4870
rect 11772 4868 11828 4870
rect 11852 4868 11908 4870
rect 11612 3834 11668 3836
rect 11692 3834 11748 3836
rect 11772 3834 11828 3836
rect 11852 3834 11908 3836
rect 11612 3782 11658 3834
rect 11658 3782 11668 3834
rect 11692 3782 11722 3834
rect 11722 3782 11734 3834
rect 11734 3782 11748 3834
rect 11772 3782 11786 3834
rect 11786 3782 11798 3834
rect 11798 3782 11828 3834
rect 11852 3782 11862 3834
rect 11862 3782 11908 3834
rect 11612 3780 11668 3782
rect 11692 3780 11748 3782
rect 11772 3780 11828 3782
rect 11852 3780 11908 3782
rect 11612 2746 11668 2748
rect 11692 2746 11748 2748
rect 11772 2746 11828 2748
rect 11852 2746 11908 2748
rect 11612 2694 11658 2746
rect 11658 2694 11668 2746
rect 11692 2694 11722 2746
rect 11722 2694 11734 2746
rect 11734 2694 11748 2746
rect 11772 2694 11786 2746
rect 11786 2694 11798 2746
rect 11798 2694 11828 2746
rect 11852 2694 11862 2746
rect 11862 2694 11908 2746
rect 11612 2692 11668 2694
rect 11692 2692 11748 2694
rect 11772 2692 11828 2694
rect 11852 2692 11908 2694
rect 5218 2202 5274 2204
rect 5298 2202 5354 2204
rect 5378 2202 5434 2204
rect 5458 2202 5514 2204
rect 5218 2150 5264 2202
rect 5264 2150 5274 2202
rect 5298 2150 5328 2202
rect 5328 2150 5340 2202
rect 5340 2150 5354 2202
rect 5378 2150 5392 2202
rect 5392 2150 5404 2202
rect 5404 2150 5434 2202
rect 5458 2150 5468 2202
rect 5468 2150 5514 2202
rect 5218 2148 5274 2150
rect 5298 2148 5354 2150
rect 5378 2148 5434 2150
rect 5458 2148 5514 2150
rect 9481 2202 9537 2204
rect 9561 2202 9617 2204
rect 9641 2202 9697 2204
rect 9721 2202 9777 2204
rect 9481 2150 9527 2202
rect 9527 2150 9537 2202
rect 9561 2150 9591 2202
rect 9591 2150 9603 2202
rect 9603 2150 9617 2202
rect 9641 2150 9655 2202
rect 9655 2150 9667 2202
rect 9667 2150 9697 2202
rect 9721 2150 9731 2202
rect 9731 2150 9777 2202
rect 9481 2148 9537 2150
rect 9561 2148 9617 2150
rect 9641 2148 9697 2150
rect 9721 2148 9777 2150
<< metal3 >>
rect 0 15602 800 15632
rect 1485 15602 1551 15605
rect 0 15600 1551 15602
rect 0 15544 1490 15600
rect 1546 15544 1551 15600
rect 0 15542 1551 15544
rect 0 15512 800 15542
rect 1485 15539 1551 15542
rect 3075 14720 3395 14721
rect 3075 14656 3083 14720
rect 3147 14656 3163 14720
rect 3227 14656 3243 14720
rect 3307 14656 3323 14720
rect 3387 14656 3395 14720
rect 3075 14655 3395 14656
rect 7338 14720 7658 14721
rect 7338 14656 7346 14720
rect 7410 14656 7426 14720
rect 7490 14656 7506 14720
rect 7570 14656 7586 14720
rect 7650 14656 7658 14720
rect 7338 14655 7658 14656
rect 11600 14720 11920 14721
rect 11600 14656 11608 14720
rect 11672 14656 11688 14720
rect 11752 14656 11768 14720
rect 11832 14656 11848 14720
rect 11912 14656 11920 14720
rect 11600 14655 11920 14656
rect 5206 14176 5526 14177
rect 5206 14112 5214 14176
rect 5278 14112 5294 14176
rect 5358 14112 5374 14176
rect 5438 14112 5454 14176
rect 5518 14112 5526 14176
rect 5206 14111 5526 14112
rect 9469 14176 9789 14177
rect 9469 14112 9477 14176
rect 9541 14112 9557 14176
rect 9621 14112 9637 14176
rect 9701 14112 9717 14176
rect 9781 14112 9789 14176
rect 9469 14111 9789 14112
rect 3075 13632 3395 13633
rect 3075 13568 3083 13632
rect 3147 13568 3163 13632
rect 3227 13568 3243 13632
rect 3307 13568 3323 13632
rect 3387 13568 3395 13632
rect 3075 13567 3395 13568
rect 7338 13632 7658 13633
rect 7338 13568 7346 13632
rect 7410 13568 7426 13632
rect 7490 13568 7506 13632
rect 7570 13568 7586 13632
rect 7650 13568 7658 13632
rect 7338 13567 7658 13568
rect 11600 13632 11920 13633
rect 11600 13568 11608 13632
rect 11672 13568 11688 13632
rect 11752 13568 11768 13632
rect 11832 13568 11848 13632
rect 11912 13568 11920 13632
rect 11600 13567 11920 13568
rect 13169 13154 13235 13157
rect 14220 13154 15020 13184
rect 13169 13152 15020 13154
rect 13169 13096 13174 13152
rect 13230 13096 15020 13152
rect 13169 13094 15020 13096
rect 13169 13091 13235 13094
rect 5206 13088 5526 13089
rect 5206 13024 5214 13088
rect 5278 13024 5294 13088
rect 5358 13024 5374 13088
rect 5438 13024 5454 13088
rect 5518 13024 5526 13088
rect 5206 13023 5526 13024
rect 9469 13088 9789 13089
rect 9469 13024 9477 13088
rect 9541 13024 9557 13088
rect 9621 13024 9637 13088
rect 9701 13024 9717 13088
rect 9781 13024 9789 13088
rect 14220 13064 15020 13094
rect 9469 13023 9789 13024
rect 3075 12544 3395 12545
rect 3075 12480 3083 12544
rect 3147 12480 3163 12544
rect 3227 12480 3243 12544
rect 3307 12480 3323 12544
rect 3387 12480 3395 12544
rect 3075 12479 3395 12480
rect 7338 12544 7658 12545
rect 7338 12480 7346 12544
rect 7410 12480 7426 12544
rect 7490 12480 7506 12544
rect 7570 12480 7586 12544
rect 7650 12480 7658 12544
rect 7338 12479 7658 12480
rect 11600 12544 11920 12545
rect 11600 12480 11608 12544
rect 11672 12480 11688 12544
rect 11752 12480 11768 12544
rect 11832 12480 11848 12544
rect 11912 12480 11920 12544
rect 11600 12479 11920 12480
rect 5206 12000 5526 12001
rect 5206 11936 5214 12000
rect 5278 11936 5294 12000
rect 5358 11936 5374 12000
rect 5438 11936 5454 12000
rect 5518 11936 5526 12000
rect 5206 11935 5526 11936
rect 9469 12000 9789 12001
rect 9469 11936 9477 12000
rect 9541 11936 9557 12000
rect 9621 11936 9637 12000
rect 9701 11936 9717 12000
rect 9781 11936 9789 12000
rect 9469 11935 9789 11936
rect 0 11794 800 11824
rect 1485 11794 1551 11797
rect 0 11792 1551 11794
rect 0 11736 1490 11792
rect 1546 11736 1551 11792
rect 0 11734 1551 11736
rect 0 11704 800 11734
rect 1485 11731 1551 11734
rect 3075 11456 3395 11457
rect 3075 11392 3083 11456
rect 3147 11392 3163 11456
rect 3227 11392 3243 11456
rect 3307 11392 3323 11456
rect 3387 11392 3395 11456
rect 3075 11391 3395 11392
rect 7338 11456 7658 11457
rect 7338 11392 7346 11456
rect 7410 11392 7426 11456
rect 7490 11392 7506 11456
rect 7570 11392 7586 11456
rect 7650 11392 7658 11456
rect 7338 11391 7658 11392
rect 11600 11456 11920 11457
rect 11600 11392 11608 11456
rect 11672 11392 11688 11456
rect 11752 11392 11768 11456
rect 11832 11392 11848 11456
rect 11912 11392 11920 11456
rect 11600 11391 11920 11392
rect 5206 10912 5526 10913
rect 5206 10848 5214 10912
rect 5278 10848 5294 10912
rect 5358 10848 5374 10912
rect 5438 10848 5454 10912
rect 5518 10848 5526 10912
rect 5206 10847 5526 10848
rect 9469 10912 9789 10913
rect 9469 10848 9477 10912
rect 9541 10848 9557 10912
rect 9621 10848 9637 10912
rect 9701 10848 9717 10912
rect 9781 10848 9789 10912
rect 9469 10847 9789 10848
rect 3075 10368 3395 10369
rect 3075 10304 3083 10368
rect 3147 10304 3163 10368
rect 3227 10304 3243 10368
rect 3307 10304 3323 10368
rect 3387 10304 3395 10368
rect 3075 10303 3395 10304
rect 7338 10368 7658 10369
rect 7338 10304 7346 10368
rect 7410 10304 7426 10368
rect 7490 10304 7506 10368
rect 7570 10304 7586 10368
rect 7650 10304 7658 10368
rect 7338 10303 7658 10304
rect 11600 10368 11920 10369
rect 11600 10304 11608 10368
rect 11672 10304 11688 10368
rect 11752 10304 11768 10368
rect 11832 10304 11848 10368
rect 11912 10304 11920 10368
rect 11600 10303 11920 10304
rect 5206 9824 5526 9825
rect 5206 9760 5214 9824
rect 5278 9760 5294 9824
rect 5358 9760 5374 9824
rect 5438 9760 5454 9824
rect 5518 9760 5526 9824
rect 5206 9759 5526 9760
rect 9469 9824 9789 9825
rect 9469 9760 9477 9824
rect 9541 9760 9557 9824
rect 9621 9760 9637 9824
rect 9701 9760 9717 9824
rect 9781 9760 9789 9824
rect 9469 9759 9789 9760
rect 13169 9346 13235 9349
rect 14220 9346 15020 9376
rect 13169 9344 15020 9346
rect 13169 9288 13174 9344
rect 13230 9288 15020 9344
rect 13169 9286 15020 9288
rect 13169 9283 13235 9286
rect 3075 9280 3395 9281
rect 3075 9216 3083 9280
rect 3147 9216 3163 9280
rect 3227 9216 3243 9280
rect 3307 9216 3323 9280
rect 3387 9216 3395 9280
rect 3075 9215 3395 9216
rect 7338 9280 7658 9281
rect 7338 9216 7346 9280
rect 7410 9216 7426 9280
rect 7490 9216 7506 9280
rect 7570 9216 7586 9280
rect 7650 9216 7658 9280
rect 7338 9215 7658 9216
rect 11600 9280 11920 9281
rect 11600 9216 11608 9280
rect 11672 9216 11688 9280
rect 11752 9216 11768 9280
rect 11832 9216 11848 9280
rect 11912 9216 11920 9280
rect 14220 9256 15020 9286
rect 11600 9215 11920 9216
rect 5206 8736 5526 8737
rect 5206 8672 5214 8736
rect 5278 8672 5294 8736
rect 5358 8672 5374 8736
rect 5438 8672 5454 8736
rect 5518 8672 5526 8736
rect 5206 8671 5526 8672
rect 9469 8736 9789 8737
rect 9469 8672 9477 8736
rect 9541 8672 9557 8736
rect 9621 8672 9637 8736
rect 9701 8672 9717 8736
rect 9781 8672 9789 8736
rect 9469 8671 9789 8672
rect 3075 8192 3395 8193
rect 3075 8128 3083 8192
rect 3147 8128 3163 8192
rect 3227 8128 3243 8192
rect 3307 8128 3323 8192
rect 3387 8128 3395 8192
rect 3075 8127 3395 8128
rect 7338 8192 7658 8193
rect 7338 8128 7346 8192
rect 7410 8128 7426 8192
rect 7490 8128 7506 8192
rect 7570 8128 7586 8192
rect 7650 8128 7658 8192
rect 7338 8127 7658 8128
rect 11600 8192 11920 8193
rect 11600 8128 11608 8192
rect 11672 8128 11688 8192
rect 11752 8128 11768 8192
rect 11832 8128 11848 8192
rect 11912 8128 11920 8192
rect 11600 8127 11920 8128
rect 0 7714 800 7744
rect 1485 7714 1551 7717
rect 0 7712 1551 7714
rect 0 7656 1490 7712
rect 1546 7656 1551 7712
rect 0 7654 1551 7656
rect 0 7624 800 7654
rect 1485 7651 1551 7654
rect 5206 7648 5526 7649
rect 5206 7584 5214 7648
rect 5278 7584 5294 7648
rect 5358 7584 5374 7648
rect 5438 7584 5454 7648
rect 5518 7584 5526 7648
rect 5206 7583 5526 7584
rect 9469 7648 9789 7649
rect 9469 7584 9477 7648
rect 9541 7584 9557 7648
rect 9621 7584 9637 7648
rect 9701 7584 9717 7648
rect 9781 7584 9789 7648
rect 9469 7583 9789 7584
rect 3075 7104 3395 7105
rect 3075 7040 3083 7104
rect 3147 7040 3163 7104
rect 3227 7040 3243 7104
rect 3307 7040 3323 7104
rect 3387 7040 3395 7104
rect 3075 7039 3395 7040
rect 7338 7104 7658 7105
rect 7338 7040 7346 7104
rect 7410 7040 7426 7104
rect 7490 7040 7506 7104
rect 7570 7040 7586 7104
rect 7650 7040 7658 7104
rect 7338 7039 7658 7040
rect 11600 7104 11920 7105
rect 11600 7040 11608 7104
rect 11672 7040 11688 7104
rect 11752 7040 11768 7104
rect 11832 7040 11848 7104
rect 11912 7040 11920 7104
rect 11600 7039 11920 7040
rect 5206 6560 5526 6561
rect 5206 6496 5214 6560
rect 5278 6496 5294 6560
rect 5358 6496 5374 6560
rect 5438 6496 5454 6560
rect 5518 6496 5526 6560
rect 5206 6495 5526 6496
rect 9469 6560 9789 6561
rect 9469 6496 9477 6560
rect 9541 6496 9557 6560
rect 9621 6496 9637 6560
rect 9701 6496 9717 6560
rect 9781 6496 9789 6560
rect 9469 6495 9789 6496
rect 3075 6016 3395 6017
rect 3075 5952 3083 6016
rect 3147 5952 3163 6016
rect 3227 5952 3243 6016
rect 3307 5952 3323 6016
rect 3387 5952 3395 6016
rect 3075 5951 3395 5952
rect 7338 6016 7658 6017
rect 7338 5952 7346 6016
rect 7410 5952 7426 6016
rect 7490 5952 7506 6016
rect 7570 5952 7586 6016
rect 7650 5952 7658 6016
rect 7338 5951 7658 5952
rect 11600 6016 11920 6017
rect 11600 5952 11608 6016
rect 11672 5952 11688 6016
rect 11752 5952 11768 6016
rect 11832 5952 11848 6016
rect 11912 5952 11920 6016
rect 11600 5951 11920 5952
rect 5206 5472 5526 5473
rect 5206 5408 5214 5472
rect 5278 5408 5294 5472
rect 5358 5408 5374 5472
rect 5438 5408 5454 5472
rect 5518 5408 5526 5472
rect 5206 5407 5526 5408
rect 9469 5472 9789 5473
rect 9469 5408 9477 5472
rect 9541 5408 9557 5472
rect 9621 5408 9637 5472
rect 9701 5408 9717 5472
rect 9781 5408 9789 5472
rect 9469 5407 9789 5408
rect 13077 5266 13143 5269
rect 14220 5266 14794 5296
rect 13077 5264 14794 5266
rect 13077 5208 13082 5264
rect 13138 5208 14794 5264
rect 13077 5206 14794 5208
rect 13077 5203 13143 5206
rect 14220 5176 14794 5206
rect 3075 4928 3395 4929
rect 3075 4864 3083 4928
rect 3147 4864 3163 4928
rect 3227 4864 3243 4928
rect 3307 4864 3323 4928
rect 3387 4864 3395 4928
rect 3075 4863 3395 4864
rect 7338 4928 7658 4929
rect 7338 4864 7346 4928
rect 7410 4864 7426 4928
rect 7490 4864 7506 4928
rect 7570 4864 7586 4928
rect 7650 4864 7658 4928
rect 7338 4863 7658 4864
rect 11600 4928 11920 4929
rect 11600 4864 11608 4928
rect 11672 4864 11688 4928
rect 11752 4864 11768 4928
rect 11832 4864 11848 4928
rect 11912 4864 11920 4928
rect 11600 4863 11920 4864
rect 5206 4384 5526 4385
rect 5206 4320 5214 4384
rect 5278 4320 5294 4384
rect 5358 4320 5374 4384
rect 5438 4320 5454 4384
rect 5518 4320 5526 4384
rect 5206 4319 5526 4320
rect 9469 4384 9789 4385
rect 9469 4320 9477 4384
rect 9541 4320 9557 4384
rect 9621 4320 9637 4384
rect 9701 4320 9717 4384
rect 9781 4320 9789 4384
rect 9469 4319 9789 4320
rect 0 3906 800 3936
rect 1485 3906 1551 3909
rect 0 3904 1551 3906
rect 0 3848 1490 3904
rect 1546 3848 1551 3904
rect 0 3846 1551 3848
rect 0 3816 800 3846
rect 1485 3843 1551 3846
rect 3075 3840 3395 3841
rect 3075 3776 3083 3840
rect 3147 3776 3163 3840
rect 3227 3776 3243 3840
rect 3307 3776 3323 3840
rect 3387 3776 3395 3840
rect 3075 3775 3395 3776
rect 7338 3840 7658 3841
rect 7338 3776 7346 3840
rect 7410 3776 7426 3840
rect 7490 3776 7506 3840
rect 7570 3776 7586 3840
rect 7650 3776 7658 3840
rect 7338 3775 7658 3776
rect 11600 3840 11920 3841
rect 11600 3776 11608 3840
rect 11672 3776 11688 3840
rect 11752 3776 11768 3840
rect 11832 3776 11848 3840
rect 11912 3776 11920 3840
rect 11600 3775 11920 3776
rect 5206 3296 5526 3297
rect 5206 3232 5214 3296
rect 5278 3232 5294 3296
rect 5358 3232 5374 3296
rect 5438 3232 5454 3296
rect 5518 3232 5526 3296
rect 5206 3231 5526 3232
rect 9469 3296 9789 3297
rect 9469 3232 9477 3296
rect 9541 3232 9557 3296
rect 9621 3232 9637 3296
rect 9701 3232 9717 3296
rect 9781 3232 9789 3296
rect 9469 3231 9789 3232
rect 3075 2752 3395 2753
rect 3075 2688 3083 2752
rect 3147 2688 3163 2752
rect 3227 2688 3243 2752
rect 3307 2688 3323 2752
rect 3387 2688 3395 2752
rect 3075 2687 3395 2688
rect 7338 2752 7658 2753
rect 7338 2688 7346 2752
rect 7410 2688 7426 2752
rect 7490 2688 7506 2752
rect 7570 2688 7586 2752
rect 7650 2688 7658 2752
rect 7338 2687 7658 2688
rect 11600 2752 11920 2753
rect 11600 2688 11608 2752
rect 11672 2688 11688 2752
rect 11752 2688 11768 2752
rect 11832 2688 11848 2752
rect 11912 2688 11920 2752
rect 11600 2687 11920 2688
rect 5206 2208 5526 2209
rect 5206 2144 5214 2208
rect 5278 2144 5294 2208
rect 5358 2144 5374 2208
rect 5438 2144 5454 2208
rect 5518 2144 5526 2208
rect 5206 2143 5526 2144
rect 9469 2208 9789 2209
rect 9469 2144 9477 2208
rect 9541 2144 9557 2208
rect 9621 2144 9637 2208
rect 9701 2144 9717 2208
rect 9781 2144 9789 2208
rect 9469 2143 9789 2144
<< via3 >>
rect 3083 14716 3147 14720
rect 3083 14660 3087 14716
rect 3087 14660 3143 14716
rect 3143 14660 3147 14716
rect 3083 14656 3147 14660
rect 3163 14716 3227 14720
rect 3163 14660 3167 14716
rect 3167 14660 3223 14716
rect 3223 14660 3227 14716
rect 3163 14656 3227 14660
rect 3243 14716 3307 14720
rect 3243 14660 3247 14716
rect 3247 14660 3303 14716
rect 3303 14660 3307 14716
rect 3243 14656 3307 14660
rect 3323 14716 3387 14720
rect 3323 14660 3327 14716
rect 3327 14660 3383 14716
rect 3383 14660 3387 14716
rect 3323 14656 3387 14660
rect 7346 14716 7410 14720
rect 7346 14660 7350 14716
rect 7350 14660 7406 14716
rect 7406 14660 7410 14716
rect 7346 14656 7410 14660
rect 7426 14716 7490 14720
rect 7426 14660 7430 14716
rect 7430 14660 7486 14716
rect 7486 14660 7490 14716
rect 7426 14656 7490 14660
rect 7506 14716 7570 14720
rect 7506 14660 7510 14716
rect 7510 14660 7566 14716
rect 7566 14660 7570 14716
rect 7506 14656 7570 14660
rect 7586 14716 7650 14720
rect 7586 14660 7590 14716
rect 7590 14660 7646 14716
rect 7646 14660 7650 14716
rect 7586 14656 7650 14660
rect 11608 14716 11672 14720
rect 11608 14660 11612 14716
rect 11612 14660 11668 14716
rect 11668 14660 11672 14716
rect 11608 14656 11672 14660
rect 11688 14716 11752 14720
rect 11688 14660 11692 14716
rect 11692 14660 11748 14716
rect 11748 14660 11752 14716
rect 11688 14656 11752 14660
rect 11768 14716 11832 14720
rect 11768 14660 11772 14716
rect 11772 14660 11828 14716
rect 11828 14660 11832 14716
rect 11768 14656 11832 14660
rect 11848 14716 11912 14720
rect 11848 14660 11852 14716
rect 11852 14660 11908 14716
rect 11908 14660 11912 14716
rect 11848 14656 11912 14660
rect 5214 14172 5278 14176
rect 5214 14116 5218 14172
rect 5218 14116 5274 14172
rect 5274 14116 5278 14172
rect 5214 14112 5278 14116
rect 5294 14172 5358 14176
rect 5294 14116 5298 14172
rect 5298 14116 5354 14172
rect 5354 14116 5358 14172
rect 5294 14112 5358 14116
rect 5374 14172 5438 14176
rect 5374 14116 5378 14172
rect 5378 14116 5434 14172
rect 5434 14116 5438 14172
rect 5374 14112 5438 14116
rect 5454 14172 5518 14176
rect 5454 14116 5458 14172
rect 5458 14116 5514 14172
rect 5514 14116 5518 14172
rect 5454 14112 5518 14116
rect 9477 14172 9541 14176
rect 9477 14116 9481 14172
rect 9481 14116 9537 14172
rect 9537 14116 9541 14172
rect 9477 14112 9541 14116
rect 9557 14172 9621 14176
rect 9557 14116 9561 14172
rect 9561 14116 9617 14172
rect 9617 14116 9621 14172
rect 9557 14112 9621 14116
rect 9637 14172 9701 14176
rect 9637 14116 9641 14172
rect 9641 14116 9697 14172
rect 9697 14116 9701 14172
rect 9637 14112 9701 14116
rect 9717 14172 9781 14176
rect 9717 14116 9721 14172
rect 9721 14116 9777 14172
rect 9777 14116 9781 14172
rect 9717 14112 9781 14116
rect 3083 13628 3147 13632
rect 3083 13572 3087 13628
rect 3087 13572 3143 13628
rect 3143 13572 3147 13628
rect 3083 13568 3147 13572
rect 3163 13628 3227 13632
rect 3163 13572 3167 13628
rect 3167 13572 3223 13628
rect 3223 13572 3227 13628
rect 3163 13568 3227 13572
rect 3243 13628 3307 13632
rect 3243 13572 3247 13628
rect 3247 13572 3303 13628
rect 3303 13572 3307 13628
rect 3243 13568 3307 13572
rect 3323 13628 3387 13632
rect 3323 13572 3327 13628
rect 3327 13572 3383 13628
rect 3383 13572 3387 13628
rect 3323 13568 3387 13572
rect 7346 13628 7410 13632
rect 7346 13572 7350 13628
rect 7350 13572 7406 13628
rect 7406 13572 7410 13628
rect 7346 13568 7410 13572
rect 7426 13628 7490 13632
rect 7426 13572 7430 13628
rect 7430 13572 7486 13628
rect 7486 13572 7490 13628
rect 7426 13568 7490 13572
rect 7506 13628 7570 13632
rect 7506 13572 7510 13628
rect 7510 13572 7566 13628
rect 7566 13572 7570 13628
rect 7506 13568 7570 13572
rect 7586 13628 7650 13632
rect 7586 13572 7590 13628
rect 7590 13572 7646 13628
rect 7646 13572 7650 13628
rect 7586 13568 7650 13572
rect 11608 13628 11672 13632
rect 11608 13572 11612 13628
rect 11612 13572 11668 13628
rect 11668 13572 11672 13628
rect 11608 13568 11672 13572
rect 11688 13628 11752 13632
rect 11688 13572 11692 13628
rect 11692 13572 11748 13628
rect 11748 13572 11752 13628
rect 11688 13568 11752 13572
rect 11768 13628 11832 13632
rect 11768 13572 11772 13628
rect 11772 13572 11828 13628
rect 11828 13572 11832 13628
rect 11768 13568 11832 13572
rect 11848 13628 11912 13632
rect 11848 13572 11852 13628
rect 11852 13572 11908 13628
rect 11908 13572 11912 13628
rect 11848 13568 11912 13572
rect 5214 13084 5278 13088
rect 5214 13028 5218 13084
rect 5218 13028 5274 13084
rect 5274 13028 5278 13084
rect 5214 13024 5278 13028
rect 5294 13084 5358 13088
rect 5294 13028 5298 13084
rect 5298 13028 5354 13084
rect 5354 13028 5358 13084
rect 5294 13024 5358 13028
rect 5374 13084 5438 13088
rect 5374 13028 5378 13084
rect 5378 13028 5434 13084
rect 5434 13028 5438 13084
rect 5374 13024 5438 13028
rect 5454 13084 5518 13088
rect 5454 13028 5458 13084
rect 5458 13028 5514 13084
rect 5514 13028 5518 13084
rect 5454 13024 5518 13028
rect 9477 13084 9541 13088
rect 9477 13028 9481 13084
rect 9481 13028 9537 13084
rect 9537 13028 9541 13084
rect 9477 13024 9541 13028
rect 9557 13084 9621 13088
rect 9557 13028 9561 13084
rect 9561 13028 9617 13084
rect 9617 13028 9621 13084
rect 9557 13024 9621 13028
rect 9637 13084 9701 13088
rect 9637 13028 9641 13084
rect 9641 13028 9697 13084
rect 9697 13028 9701 13084
rect 9637 13024 9701 13028
rect 9717 13084 9781 13088
rect 9717 13028 9721 13084
rect 9721 13028 9777 13084
rect 9777 13028 9781 13084
rect 9717 13024 9781 13028
rect 3083 12540 3147 12544
rect 3083 12484 3087 12540
rect 3087 12484 3143 12540
rect 3143 12484 3147 12540
rect 3083 12480 3147 12484
rect 3163 12540 3227 12544
rect 3163 12484 3167 12540
rect 3167 12484 3223 12540
rect 3223 12484 3227 12540
rect 3163 12480 3227 12484
rect 3243 12540 3307 12544
rect 3243 12484 3247 12540
rect 3247 12484 3303 12540
rect 3303 12484 3307 12540
rect 3243 12480 3307 12484
rect 3323 12540 3387 12544
rect 3323 12484 3327 12540
rect 3327 12484 3383 12540
rect 3383 12484 3387 12540
rect 3323 12480 3387 12484
rect 7346 12540 7410 12544
rect 7346 12484 7350 12540
rect 7350 12484 7406 12540
rect 7406 12484 7410 12540
rect 7346 12480 7410 12484
rect 7426 12540 7490 12544
rect 7426 12484 7430 12540
rect 7430 12484 7486 12540
rect 7486 12484 7490 12540
rect 7426 12480 7490 12484
rect 7506 12540 7570 12544
rect 7506 12484 7510 12540
rect 7510 12484 7566 12540
rect 7566 12484 7570 12540
rect 7506 12480 7570 12484
rect 7586 12540 7650 12544
rect 7586 12484 7590 12540
rect 7590 12484 7646 12540
rect 7646 12484 7650 12540
rect 7586 12480 7650 12484
rect 11608 12540 11672 12544
rect 11608 12484 11612 12540
rect 11612 12484 11668 12540
rect 11668 12484 11672 12540
rect 11608 12480 11672 12484
rect 11688 12540 11752 12544
rect 11688 12484 11692 12540
rect 11692 12484 11748 12540
rect 11748 12484 11752 12540
rect 11688 12480 11752 12484
rect 11768 12540 11832 12544
rect 11768 12484 11772 12540
rect 11772 12484 11828 12540
rect 11828 12484 11832 12540
rect 11768 12480 11832 12484
rect 11848 12540 11912 12544
rect 11848 12484 11852 12540
rect 11852 12484 11908 12540
rect 11908 12484 11912 12540
rect 11848 12480 11912 12484
rect 5214 11996 5278 12000
rect 5214 11940 5218 11996
rect 5218 11940 5274 11996
rect 5274 11940 5278 11996
rect 5214 11936 5278 11940
rect 5294 11996 5358 12000
rect 5294 11940 5298 11996
rect 5298 11940 5354 11996
rect 5354 11940 5358 11996
rect 5294 11936 5358 11940
rect 5374 11996 5438 12000
rect 5374 11940 5378 11996
rect 5378 11940 5434 11996
rect 5434 11940 5438 11996
rect 5374 11936 5438 11940
rect 5454 11996 5518 12000
rect 5454 11940 5458 11996
rect 5458 11940 5514 11996
rect 5514 11940 5518 11996
rect 5454 11936 5518 11940
rect 9477 11996 9541 12000
rect 9477 11940 9481 11996
rect 9481 11940 9537 11996
rect 9537 11940 9541 11996
rect 9477 11936 9541 11940
rect 9557 11996 9621 12000
rect 9557 11940 9561 11996
rect 9561 11940 9617 11996
rect 9617 11940 9621 11996
rect 9557 11936 9621 11940
rect 9637 11996 9701 12000
rect 9637 11940 9641 11996
rect 9641 11940 9697 11996
rect 9697 11940 9701 11996
rect 9637 11936 9701 11940
rect 9717 11996 9781 12000
rect 9717 11940 9721 11996
rect 9721 11940 9777 11996
rect 9777 11940 9781 11996
rect 9717 11936 9781 11940
rect 3083 11452 3147 11456
rect 3083 11396 3087 11452
rect 3087 11396 3143 11452
rect 3143 11396 3147 11452
rect 3083 11392 3147 11396
rect 3163 11452 3227 11456
rect 3163 11396 3167 11452
rect 3167 11396 3223 11452
rect 3223 11396 3227 11452
rect 3163 11392 3227 11396
rect 3243 11452 3307 11456
rect 3243 11396 3247 11452
rect 3247 11396 3303 11452
rect 3303 11396 3307 11452
rect 3243 11392 3307 11396
rect 3323 11452 3387 11456
rect 3323 11396 3327 11452
rect 3327 11396 3383 11452
rect 3383 11396 3387 11452
rect 3323 11392 3387 11396
rect 7346 11452 7410 11456
rect 7346 11396 7350 11452
rect 7350 11396 7406 11452
rect 7406 11396 7410 11452
rect 7346 11392 7410 11396
rect 7426 11452 7490 11456
rect 7426 11396 7430 11452
rect 7430 11396 7486 11452
rect 7486 11396 7490 11452
rect 7426 11392 7490 11396
rect 7506 11452 7570 11456
rect 7506 11396 7510 11452
rect 7510 11396 7566 11452
rect 7566 11396 7570 11452
rect 7506 11392 7570 11396
rect 7586 11452 7650 11456
rect 7586 11396 7590 11452
rect 7590 11396 7646 11452
rect 7646 11396 7650 11452
rect 7586 11392 7650 11396
rect 11608 11452 11672 11456
rect 11608 11396 11612 11452
rect 11612 11396 11668 11452
rect 11668 11396 11672 11452
rect 11608 11392 11672 11396
rect 11688 11452 11752 11456
rect 11688 11396 11692 11452
rect 11692 11396 11748 11452
rect 11748 11396 11752 11452
rect 11688 11392 11752 11396
rect 11768 11452 11832 11456
rect 11768 11396 11772 11452
rect 11772 11396 11828 11452
rect 11828 11396 11832 11452
rect 11768 11392 11832 11396
rect 11848 11452 11912 11456
rect 11848 11396 11852 11452
rect 11852 11396 11908 11452
rect 11908 11396 11912 11452
rect 11848 11392 11912 11396
rect 5214 10908 5278 10912
rect 5214 10852 5218 10908
rect 5218 10852 5274 10908
rect 5274 10852 5278 10908
rect 5214 10848 5278 10852
rect 5294 10908 5358 10912
rect 5294 10852 5298 10908
rect 5298 10852 5354 10908
rect 5354 10852 5358 10908
rect 5294 10848 5358 10852
rect 5374 10908 5438 10912
rect 5374 10852 5378 10908
rect 5378 10852 5434 10908
rect 5434 10852 5438 10908
rect 5374 10848 5438 10852
rect 5454 10908 5518 10912
rect 5454 10852 5458 10908
rect 5458 10852 5514 10908
rect 5514 10852 5518 10908
rect 5454 10848 5518 10852
rect 9477 10908 9541 10912
rect 9477 10852 9481 10908
rect 9481 10852 9537 10908
rect 9537 10852 9541 10908
rect 9477 10848 9541 10852
rect 9557 10908 9621 10912
rect 9557 10852 9561 10908
rect 9561 10852 9617 10908
rect 9617 10852 9621 10908
rect 9557 10848 9621 10852
rect 9637 10908 9701 10912
rect 9637 10852 9641 10908
rect 9641 10852 9697 10908
rect 9697 10852 9701 10908
rect 9637 10848 9701 10852
rect 9717 10908 9781 10912
rect 9717 10852 9721 10908
rect 9721 10852 9777 10908
rect 9777 10852 9781 10908
rect 9717 10848 9781 10852
rect 3083 10364 3147 10368
rect 3083 10308 3087 10364
rect 3087 10308 3143 10364
rect 3143 10308 3147 10364
rect 3083 10304 3147 10308
rect 3163 10364 3227 10368
rect 3163 10308 3167 10364
rect 3167 10308 3223 10364
rect 3223 10308 3227 10364
rect 3163 10304 3227 10308
rect 3243 10364 3307 10368
rect 3243 10308 3247 10364
rect 3247 10308 3303 10364
rect 3303 10308 3307 10364
rect 3243 10304 3307 10308
rect 3323 10364 3387 10368
rect 3323 10308 3327 10364
rect 3327 10308 3383 10364
rect 3383 10308 3387 10364
rect 3323 10304 3387 10308
rect 7346 10364 7410 10368
rect 7346 10308 7350 10364
rect 7350 10308 7406 10364
rect 7406 10308 7410 10364
rect 7346 10304 7410 10308
rect 7426 10364 7490 10368
rect 7426 10308 7430 10364
rect 7430 10308 7486 10364
rect 7486 10308 7490 10364
rect 7426 10304 7490 10308
rect 7506 10364 7570 10368
rect 7506 10308 7510 10364
rect 7510 10308 7566 10364
rect 7566 10308 7570 10364
rect 7506 10304 7570 10308
rect 7586 10364 7650 10368
rect 7586 10308 7590 10364
rect 7590 10308 7646 10364
rect 7646 10308 7650 10364
rect 7586 10304 7650 10308
rect 11608 10364 11672 10368
rect 11608 10308 11612 10364
rect 11612 10308 11668 10364
rect 11668 10308 11672 10364
rect 11608 10304 11672 10308
rect 11688 10364 11752 10368
rect 11688 10308 11692 10364
rect 11692 10308 11748 10364
rect 11748 10308 11752 10364
rect 11688 10304 11752 10308
rect 11768 10364 11832 10368
rect 11768 10308 11772 10364
rect 11772 10308 11828 10364
rect 11828 10308 11832 10364
rect 11768 10304 11832 10308
rect 11848 10364 11912 10368
rect 11848 10308 11852 10364
rect 11852 10308 11908 10364
rect 11908 10308 11912 10364
rect 11848 10304 11912 10308
rect 5214 9820 5278 9824
rect 5214 9764 5218 9820
rect 5218 9764 5274 9820
rect 5274 9764 5278 9820
rect 5214 9760 5278 9764
rect 5294 9820 5358 9824
rect 5294 9764 5298 9820
rect 5298 9764 5354 9820
rect 5354 9764 5358 9820
rect 5294 9760 5358 9764
rect 5374 9820 5438 9824
rect 5374 9764 5378 9820
rect 5378 9764 5434 9820
rect 5434 9764 5438 9820
rect 5374 9760 5438 9764
rect 5454 9820 5518 9824
rect 5454 9764 5458 9820
rect 5458 9764 5514 9820
rect 5514 9764 5518 9820
rect 5454 9760 5518 9764
rect 9477 9820 9541 9824
rect 9477 9764 9481 9820
rect 9481 9764 9537 9820
rect 9537 9764 9541 9820
rect 9477 9760 9541 9764
rect 9557 9820 9621 9824
rect 9557 9764 9561 9820
rect 9561 9764 9617 9820
rect 9617 9764 9621 9820
rect 9557 9760 9621 9764
rect 9637 9820 9701 9824
rect 9637 9764 9641 9820
rect 9641 9764 9697 9820
rect 9697 9764 9701 9820
rect 9637 9760 9701 9764
rect 9717 9820 9781 9824
rect 9717 9764 9721 9820
rect 9721 9764 9777 9820
rect 9777 9764 9781 9820
rect 9717 9760 9781 9764
rect 3083 9276 3147 9280
rect 3083 9220 3087 9276
rect 3087 9220 3143 9276
rect 3143 9220 3147 9276
rect 3083 9216 3147 9220
rect 3163 9276 3227 9280
rect 3163 9220 3167 9276
rect 3167 9220 3223 9276
rect 3223 9220 3227 9276
rect 3163 9216 3227 9220
rect 3243 9276 3307 9280
rect 3243 9220 3247 9276
rect 3247 9220 3303 9276
rect 3303 9220 3307 9276
rect 3243 9216 3307 9220
rect 3323 9276 3387 9280
rect 3323 9220 3327 9276
rect 3327 9220 3383 9276
rect 3383 9220 3387 9276
rect 3323 9216 3387 9220
rect 7346 9276 7410 9280
rect 7346 9220 7350 9276
rect 7350 9220 7406 9276
rect 7406 9220 7410 9276
rect 7346 9216 7410 9220
rect 7426 9276 7490 9280
rect 7426 9220 7430 9276
rect 7430 9220 7486 9276
rect 7486 9220 7490 9276
rect 7426 9216 7490 9220
rect 7506 9276 7570 9280
rect 7506 9220 7510 9276
rect 7510 9220 7566 9276
rect 7566 9220 7570 9276
rect 7506 9216 7570 9220
rect 7586 9276 7650 9280
rect 7586 9220 7590 9276
rect 7590 9220 7646 9276
rect 7646 9220 7650 9276
rect 7586 9216 7650 9220
rect 11608 9276 11672 9280
rect 11608 9220 11612 9276
rect 11612 9220 11668 9276
rect 11668 9220 11672 9276
rect 11608 9216 11672 9220
rect 11688 9276 11752 9280
rect 11688 9220 11692 9276
rect 11692 9220 11748 9276
rect 11748 9220 11752 9276
rect 11688 9216 11752 9220
rect 11768 9276 11832 9280
rect 11768 9220 11772 9276
rect 11772 9220 11828 9276
rect 11828 9220 11832 9276
rect 11768 9216 11832 9220
rect 11848 9276 11912 9280
rect 11848 9220 11852 9276
rect 11852 9220 11908 9276
rect 11908 9220 11912 9276
rect 11848 9216 11912 9220
rect 5214 8732 5278 8736
rect 5214 8676 5218 8732
rect 5218 8676 5274 8732
rect 5274 8676 5278 8732
rect 5214 8672 5278 8676
rect 5294 8732 5358 8736
rect 5294 8676 5298 8732
rect 5298 8676 5354 8732
rect 5354 8676 5358 8732
rect 5294 8672 5358 8676
rect 5374 8732 5438 8736
rect 5374 8676 5378 8732
rect 5378 8676 5434 8732
rect 5434 8676 5438 8732
rect 5374 8672 5438 8676
rect 5454 8732 5518 8736
rect 5454 8676 5458 8732
rect 5458 8676 5514 8732
rect 5514 8676 5518 8732
rect 5454 8672 5518 8676
rect 9477 8732 9541 8736
rect 9477 8676 9481 8732
rect 9481 8676 9537 8732
rect 9537 8676 9541 8732
rect 9477 8672 9541 8676
rect 9557 8732 9621 8736
rect 9557 8676 9561 8732
rect 9561 8676 9617 8732
rect 9617 8676 9621 8732
rect 9557 8672 9621 8676
rect 9637 8732 9701 8736
rect 9637 8676 9641 8732
rect 9641 8676 9697 8732
rect 9697 8676 9701 8732
rect 9637 8672 9701 8676
rect 9717 8732 9781 8736
rect 9717 8676 9721 8732
rect 9721 8676 9777 8732
rect 9777 8676 9781 8732
rect 9717 8672 9781 8676
rect 3083 8188 3147 8192
rect 3083 8132 3087 8188
rect 3087 8132 3143 8188
rect 3143 8132 3147 8188
rect 3083 8128 3147 8132
rect 3163 8188 3227 8192
rect 3163 8132 3167 8188
rect 3167 8132 3223 8188
rect 3223 8132 3227 8188
rect 3163 8128 3227 8132
rect 3243 8188 3307 8192
rect 3243 8132 3247 8188
rect 3247 8132 3303 8188
rect 3303 8132 3307 8188
rect 3243 8128 3307 8132
rect 3323 8188 3387 8192
rect 3323 8132 3327 8188
rect 3327 8132 3383 8188
rect 3383 8132 3387 8188
rect 3323 8128 3387 8132
rect 7346 8188 7410 8192
rect 7346 8132 7350 8188
rect 7350 8132 7406 8188
rect 7406 8132 7410 8188
rect 7346 8128 7410 8132
rect 7426 8188 7490 8192
rect 7426 8132 7430 8188
rect 7430 8132 7486 8188
rect 7486 8132 7490 8188
rect 7426 8128 7490 8132
rect 7506 8188 7570 8192
rect 7506 8132 7510 8188
rect 7510 8132 7566 8188
rect 7566 8132 7570 8188
rect 7506 8128 7570 8132
rect 7586 8188 7650 8192
rect 7586 8132 7590 8188
rect 7590 8132 7646 8188
rect 7646 8132 7650 8188
rect 7586 8128 7650 8132
rect 11608 8188 11672 8192
rect 11608 8132 11612 8188
rect 11612 8132 11668 8188
rect 11668 8132 11672 8188
rect 11608 8128 11672 8132
rect 11688 8188 11752 8192
rect 11688 8132 11692 8188
rect 11692 8132 11748 8188
rect 11748 8132 11752 8188
rect 11688 8128 11752 8132
rect 11768 8188 11832 8192
rect 11768 8132 11772 8188
rect 11772 8132 11828 8188
rect 11828 8132 11832 8188
rect 11768 8128 11832 8132
rect 11848 8188 11912 8192
rect 11848 8132 11852 8188
rect 11852 8132 11908 8188
rect 11908 8132 11912 8188
rect 11848 8128 11912 8132
rect 5214 7644 5278 7648
rect 5214 7588 5218 7644
rect 5218 7588 5274 7644
rect 5274 7588 5278 7644
rect 5214 7584 5278 7588
rect 5294 7644 5358 7648
rect 5294 7588 5298 7644
rect 5298 7588 5354 7644
rect 5354 7588 5358 7644
rect 5294 7584 5358 7588
rect 5374 7644 5438 7648
rect 5374 7588 5378 7644
rect 5378 7588 5434 7644
rect 5434 7588 5438 7644
rect 5374 7584 5438 7588
rect 5454 7644 5518 7648
rect 5454 7588 5458 7644
rect 5458 7588 5514 7644
rect 5514 7588 5518 7644
rect 5454 7584 5518 7588
rect 9477 7644 9541 7648
rect 9477 7588 9481 7644
rect 9481 7588 9537 7644
rect 9537 7588 9541 7644
rect 9477 7584 9541 7588
rect 9557 7644 9621 7648
rect 9557 7588 9561 7644
rect 9561 7588 9617 7644
rect 9617 7588 9621 7644
rect 9557 7584 9621 7588
rect 9637 7644 9701 7648
rect 9637 7588 9641 7644
rect 9641 7588 9697 7644
rect 9697 7588 9701 7644
rect 9637 7584 9701 7588
rect 9717 7644 9781 7648
rect 9717 7588 9721 7644
rect 9721 7588 9777 7644
rect 9777 7588 9781 7644
rect 9717 7584 9781 7588
rect 3083 7100 3147 7104
rect 3083 7044 3087 7100
rect 3087 7044 3143 7100
rect 3143 7044 3147 7100
rect 3083 7040 3147 7044
rect 3163 7100 3227 7104
rect 3163 7044 3167 7100
rect 3167 7044 3223 7100
rect 3223 7044 3227 7100
rect 3163 7040 3227 7044
rect 3243 7100 3307 7104
rect 3243 7044 3247 7100
rect 3247 7044 3303 7100
rect 3303 7044 3307 7100
rect 3243 7040 3307 7044
rect 3323 7100 3387 7104
rect 3323 7044 3327 7100
rect 3327 7044 3383 7100
rect 3383 7044 3387 7100
rect 3323 7040 3387 7044
rect 7346 7100 7410 7104
rect 7346 7044 7350 7100
rect 7350 7044 7406 7100
rect 7406 7044 7410 7100
rect 7346 7040 7410 7044
rect 7426 7100 7490 7104
rect 7426 7044 7430 7100
rect 7430 7044 7486 7100
rect 7486 7044 7490 7100
rect 7426 7040 7490 7044
rect 7506 7100 7570 7104
rect 7506 7044 7510 7100
rect 7510 7044 7566 7100
rect 7566 7044 7570 7100
rect 7506 7040 7570 7044
rect 7586 7100 7650 7104
rect 7586 7044 7590 7100
rect 7590 7044 7646 7100
rect 7646 7044 7650 7100
rect 7586 7040 7650 7044
rect 11608 7100 11672 7104
rect 11608 7044 11612 7100
rect 11612 7044 11668 7100
rect 11668 7044 11672 7100
rect 11608 7040 11672 7044
rect 11688 7100 11752 7104
rect 11688 7044 11692 7100
rect 11692 7044 11748 7100
rect 11748 7044 11752 7100
rect 11688 7040 11752 7044
rect 11768 7100 11832 7104
rect 11768 7044 11772 7100
rect 11772 7044 11828 7100
rect 11828 7044 11832 7100
rect 11768 7040 11832 7044
rect 11848 7100 11912 7104
rect 11848 7044 11852 7100
rect 11852 7044 11908 7100
rect 11908 7044 11912 7100
rect 11848 7040 11912 7044
rect 5214 6556 5278 6560
rect 5214 6500 5218 6556
rect 5218 6500 5274 6556
rect 5274 6500 5278 6556
rect 5214 6496 5278 6500
rect 5294 6556 5358 6560
rect 5294 6500 5298 6556
rect 5298 6500 5354 6556
rect 5354 6500 5358 6556
rect 5294 6496 5358 6500
rect 5374 6556 5438 6560
rect 5374 6500 5378 6556
rect 5378 6500 5434 6556
rect 5434 6500 5438 6556
rect 5374 6496 5438 6500
rect 5454 6556 5518 6560
rect 5454 6500 5458 6556
rect 5458 6500 5514 6556
rect 5514 6500 5518 6556
rect 5454 6496 5518 6500
rect 9477 6556 9541 6560
rect 9477 6500 9481 6556
rect 9481 6500 9537 6556
rect 9537 6500 9541 6556
rect 9477 6496 9541 6500
rect 9557 6556 9621 6560
rect 9557 6500 9561 6556
rect 9561 6500 9617 6556
rect 9617 6500 9621 6556
rect 9557 6496 9621 6500
rect 9637 6556 9701 6560
rect 9637 6500 9641 6556
rect 9641 6500 9697 6556
rect 9697 6500 9701 6556
rect 9637 6496 9701 6500
rect 9717 6556 9781 6560
rect 9717 6500 9721 6556
rect 9721 6500 9777 6556
rect 9777 6500 9781 6556
rect 9717 6496 9781 6500
rect 3083 6012 3147 6016
rect 3083 5956 3087 6012
rect 3087 5956 3143 6012
rect 3143 5956 3147 6012
rect 3083 5952 3147 5956
rect 3163 6012 3227 6016
rect 3163 5956 3167 6012
rect 3167 5956 3223 6012
rect 3223 5956 3227 6012
rect 3163 5952 3227 5956
rect 3243 6012 3307 6016
rect 3243 5956 3247 6012
rect 3247 5956 3303 6012
rect 3303 5956 3307 6012
rect 3243 5952 3307 5956
rect 3323 6012 3387 6016
rect 3323 5956 3327 6012
rect 3327 5956 3383 6012
rect 3383 5956 3387 6012
rect 3323 5952 3387 5956
rect 7346 6012 7410 6016
rect 7346 5956 7350 6012
rect 7350 5956 7406 6012
rect 7406 5956 7410 6012
rect 7346 5952 7410 5956
rect 7426 6012 7490 6016
rect 7426 5956 7430 6012
rect 7430 5956 7486 6012
rect 7486 5956 7490 6012
rect 7426 5952 7490 5956
rect 7506 6012 7570 6016
rect 7506 5956 7510 6012
rect 7510 5956 7566 6012
rect 7566 5956 7570 6012
rect 7506 5952 7570 5956
rect 7586 6012 7650 6016
rect 7586 5956 7590 6012
rect 7590 5956 7646 6012
rect 7646 5956 7650 6012
rect 7586 5952 7650 5956
rect 11608 6012 11672 6016
rect 11608 5956 11612 6012
rect 11612 5956 11668 6012
rect 11668 5956 11672 6012
rect 11608 5952 11672 5956
rect 11688 6012 11752 6016
rect 11688 5956 11692 6012
rect 11692 5956 11748 6012
rect 11748 5956 11752 6012
rect 11688 5952 11752 5956
rect 11768 6012 11832 6016
rect 11768 5956 11772 6012
rect 11772 5956 11828 6012
rect 11828 5956 11832 6012
rect 11768 5952 11832 5956
rect 11848 6012 11912 6016
rect 11848 5956 11852 6012
rect 11852 5956 11908 6012
rect 11908 5956 11912 6012
rect 11848 5952 11912 5956
rect 5214 5468 5278 5472
rect 5214 5412 5218 5468
rect 5218 5412 5274 5468
rect 5274 5412 5278 5468
rect 5214 5408 5278 5412
rect 5294 5468 5358 5472
rect 5294 5412 5298 5468
rect 5298 5412 5354 5468
rect 5354 5412 5358 5468
rect 5294 5408 5358 5412
rect 5374 5468 5438 5472
rect 5374 5412 5378 5468
rect 5378 5412 5434 5468
rect 5434 5412 5438 5468
rect 5374 5408 5438 5412
rect 5454 5468 5518 5472
rect 5454 5412 5458 5468
rect 5458 5412 5514 5468
rect 5514 5412 5518 5468
rect 5454 5408 5518 5412
rect 9477 5468 9541 5472
rect 9477 5412 9481 5468
rect 9481 5412 9537 5468
rect 9537 5412 9541 5468
rect 9477 5408 9541 5412
rect 9557 5468 9621 5472
rect 9557 5412 9561 5468
rect 9561 5412 9617 5468
rect 9617 5412 9621 5468
rect 9557 5408 9621 5412
rect 9637 5468 9701 5472
rect 9637 5412 9641 5468
rect 9641 5412 9697 5468
rect 9697 5412 9701 5468
rect 9637 5408 9701 5412
rect 9717 5468 9781 5472
rect 9717 5412 9721 5468
rect 9721 5412 9777 5468
rect 9777 5412 9781 5468
rect 9717 5408 9781 5412
rect 3083 4924 3147 4928
rect 3083 4868 3087 4924
rect 3087 4868 3143 4924
rect 3143 4868 3147 4924
rect 3083 4864 3147 4868
rect 3163 4924 3227 4928
rect 3163 4868 3167 4924
rect 3167 4868 3223 4924
rect 3223 4868 3227 4924
rect 3163 4864 3227 4868
rect 3243 4924 3307 4928
rect 3243 4868 3247 4924
rect 3247 4868 3303 4924
rect 3303 4868 3307 4924
rect 3243 4864 3307 4868
rect 3323 4924 3387 4928
rect 3323 4868 3327 4924
rect 3327 4868 3383 4924
rect 3383 4868 3387 4924
rect 3323 4864 3387 4868
rect 7346 4924 7410 4928
rect 7346 4868 7350 4924
rect 7350 4868 7406 4924
rect 7406 4868 7410 4924
rect 7346 4864 7410 4868
rect 7426 4924 7490 4928
rect 7426 4868 7430 4924
rect 7430 4868 7486 4924
rect 7486 4868 7490 4924
rect 7426 4864 7490 4868
rect 7506 4924 7570 4928
rect 7506 4868 7510 4924
rect 7510 4868 7566 4924
rect 7566 4868 7570 4924
rect 7506 4864 7570 4868
rect 7586 4924 7650 4928
rect 7586 4868 7590 4924
rect 7590 4868 7646 4924
rect 7646 4868 7650 4924
rect 7586 4864 7650 4868
rect 11608 4924 11672 4928
rect 11608 4868 11612 4924
rect 11612 4868 11668 4924
rect 11668 4868 11672 4924
rect 11608 4864 11672 4868
rect 11688 4924 11752 4928
rect 11688 4868 11692 4924
rect 11692 4868 11748 4924
rect 11748 4868 11752 4924
rect 11688 4864 11752 4868
rect 11768 4924 11832 4928
rect 11768 4868 11772 4924
rect 11772 4868 11828 4924
rect 11828 4868 11832 4924
rect 11768 4864 11832 4868
rect 11848 4924 11912 4928
rect 11848 4868 11852 4924
rect 11852 4868 11908 4924
rect 11908 4868 11912 4924
rect 11848 4864 11912 4868
rect 5214 4380 5278 4384
rect 5214 4324 5218 4380
rect 5218 4324 5274 4380
rect 5274 4324 5278 4380
rect 5214 4320 5278 4324
rect 5294 4380 5358 4384
rect 5294 4324 5298 4380
rect 5298 4324 5354 4380
rect 5354 4324 5358 4380
rect 5294 4320 5358 4324
rect 5374 4380 5438 4384
rect 5374 4324 5378 4380
rect 5378 4324 5434 4380
rect 5434 4324 5438 4380
rect 5374 4320 5438 4324
rect 5454 4380 5518 4384
rect 5454 4324 5458 4380
rect 5458 4324 5514 4380
rect 5514 4324 5518 4380
rect 5454 4320 5518 4324
rect 9477 4380 9541 4384
rect 9477 4324 9481 4380
rect 9481 4324 9537 4380
rect 9537 4324 9541 4380
rect 9477 4320 9541 4324
rect 9557 4380 9621 4384
rect 9557 4324 9561 4380
rect 9561 4324 9617 4380
rect 9617 4324 9621 4380
rect 9557 4320 9621 4324
rect 9637 4380 9701 4384
rect 9637 4324 9641 4380
rect 9641 4324 9697 4380
rect 9697 4324 9701 4380
rect 9637 4320 9701 4324
rect 9717 4380 9781 4384
rect 9717 4324 9721 4380
rect 9721 4324 9777 4380
rect 9777 4324 9781 4380
rect 9717 4320 9781 4324
rect 3083 3836 3147 3840
rect 3083 3780 3087 3836
rect 3087 3780 3143 3836
rect 3143 3780 3147 3836
rect 3083 3776 3147 3780
rect 3163 3836 3227 3840
rect 3163 3780 3167 3836
rect 3167 3780 3223 3836
rect 3223 3780 3227 3836
rect 3163 3776 3227 3780
rect 3243 3836 3307 3840
rect 3243 3780 3247 3836
rect 3247 3780 3303 3836
rect 3303 3780 3307 3836
rect 3243 3776 3307 3780
rect 3323 3836 3387 3840
rect 3323 3780 3327 3836
rect 3327 3780 3383 3836
rect 3383 3780 3387 3836
rect 3323 3776 3387 3780
rect 7346 3836 7410 3840
rect 7346 3780 7350 3836
rect 7350 3780 7406 3836
rect 7406 3780 7410 3836
rect 7346 3776 7410 3780
rect 7426 3836 7490 3840
rect 7426 3780 7430 3836
rect 7430 3780 7486 3836
rect 7486 3780 7490 3836
rect 7426 3776 7490 3780
rect 7506 3836 7570 3840
rect 7506 3780 7510 3836
rect 7510 3780 7566 3836
rect 7566 3780 7570 3836
rect 7506 3776 7570 3780
rect 7586 3836 7650 3840
rect 7586 3780 7590 3836
rect 7590 3780 7646 3836
rect 7646 3780 7650 3836
rect 7586 3776 7650 3780
rect 11608 3836 11672 3840
rect 11608 3780 11612 3836
rect 11612 3780 11668 3836
rect 11668 3780 11672 3836
rect 11608 3776 11672 3780
rect 11688 3836 11752 3840
rect 11688 3780 11692 3836
rect 11692 3780 11748 3836
rect 11748 3780 11752 3836
rect 11688 3776 11752 3780
rect 11768 3836 11832 3840
rect 11768 3780 11772 3836
rect 11772 3780 11828 3836
rect 11828 3780 11832 3836
rect 11768 3776 11832 3780
rect 11848 3836 11912 3840
rect 11848 3780 11852 3836
rect 11852 3780 11908 3836
rect 11908 3780 11912 3836
rect 11848 3776 11912 3780
rect 5214 3292 5278 3296
rect 5214 3236 5218 3292
rect 5218 3236 5274 3292
rect 5274 3236 5278 3292
rect 5214 3232 5278 3236
rect 5294 3292 5358 3296
rect 5294 3236 5298 3292
rect 5298 3236 5354 3292
rect 5354 3236 5358 3292
rect 5294 3232 5358 3236
rect 5374 3292 5438 3296
rect 5374 3236 5378 3292
rect 5378 3236 5434 3292
rect 5434 3236 5438 3292
rect 5374 3232 5438 3236
rect 5454 3292 5518 3296
rect 5454 3236 5458 3292
rect 5458 3236 5514 3292
rect 5514 3236 5518 3292
rect 5454 3232 5518 3236
rect 9477 3292 9541 3296
rect 9477 3236 9481 3292
rect 9481 3236 9537 3292
rect 9537 3236 9541 3292
rect 9477 3232 9541 3236
rect 9557 3292 9621 3296
rect 9557 3236 9561 3292
rect 9561 3236 9617 3292
rect 9617 3236 9621 3292
rect 9557 3232 9621 3236
rect 9637 3292 9701 3296
rect 9637 3236 9641 3292
rect 9641 3236 9697 3292
rect 9697 3236 9701 3292
rect 9637 3232 9701 3236
rect 9717 3292 9781 3296
rect 9717 3236 9721 3292
rect 9721 3236 9777 3292
rect 9777 3236 9781 3292
rect 9717 3232 9781 3236
rect 3083 2748 3147 2752
rect 3083 2692 3087 2748
rect 3087 2692 3143 2748
rect 3143 2692 3147 2748
rect 3083 2688 3147 2692
rect 3163 2748 3227 2752
rect 3163 2692 3167 2748
rect 3167 2692 3223 2748
rect 3223 2692 3227 2748
rect 3163 2688 3227 2692
rect 3243 2748 3307 2752
rect 3243 2692 3247 2748
rect 3247 2692 3303 2748
rect 3303 2692 3307 2748
rect 3243 2688 3307 2692
rect 3323 2748 3387 2752
rect 3323 2692 3327 2748
rect 3327 2692 3383 2748
rect 3383 2692 3387 2748
rect 3323 2688 3387 2692
rect 7346 2748 7410 2752
rect 7346 2692 7350 2748
rect 7350 2692 7406 2748
rect 7406 2692 7410 2748
rect 7346 2688 7410 2692
rect 7426 2748 7490 2752
rect 7426 2692 7430 2748
rect 7430 2692 7486 2748
rect 7486 2692 7490 2748
rect 7426 2688 7490 2692
rect 7506 2748 7570 2752
rect 7506 2692 7510 2748
rect 7510 2692 7566 2748
rect 7566 2692 7570 2748
rect 7506 2688 7570 2692
rect 7586 2748 7650 2752
rect 7586 2692 7590 2748
rect 7590 2692 7646 2748
rect 7646 2692 7650 2748
rect 7586 2688 7650 2692
rect 11608 2748 11672 2752
rect 11608 2692 11612 2748
rect 11612 2692 11668 2748
rect 11668 2692 11672 2748
rect 11608 2688 11672 2692
rect 11688 2748 11752 2752
rect 11688 2692 11692 2748
rect 11692 2692 11748 2748
rect 11748 2692 11752 2748
rect 11688 2688 11752 2692
rect 11768 2748 11832 2752
rect 11768 2692 11772 2748
rect 11772 2692 11828 2748
rect 11828 2692 11832 2748
rect 11768 2688 11832 2692
rect 11848 2748 11912 2752
rect 11848 2692 11852 2748
rect 11852 2692 11908 2748
rect 11908 2692 11912 2748
rect 11848 2688 11912 2692
rect 5214 2204 5278 2208
rect 5214 2148 5218 2204
rect 5218 2148 5274 2204
rect 5274 2148 5278 2204
rect 5214 2144 5278 2148
rect 5294 2204 5358 2208
rect 5294 2148 5298 2204
rect 5298 2148 5354 2204
rect 5354 2148 5358 2204
rect 5294 2144 5358 2148
rect 5374 2204 5438 2208
rect 5374 2148 5378 2204
rect 5378 2148 5434 2204
rect 5434 2148 5438 2204
rect 5374 2144 5438 2148
rect 5454 2204 5518 2208
rect 5454 2148 5458 2204
rect 5458 2148 5514 2204
rect 5514 2148 5518 2204
rect 5454 2144 5518 2148
rect 9477 2204 9541 2208
rect 9477 2148 9481 2204
rect 9481 2148 9537 2204
rect 9537 2148 9541 2204
rect 9477 2144 9541 2148
rect 9557 2204 9621 2208
rect 9557 2148 9561 2204
rect 9561 2148 9617 2204
rect 9617 2148 9621 2204
rect 9557 2144 9621 2148
rect 9637 2204 9701 2208
rect 9637 2148 9641 2204
rect 9641 2148 9697 2204
rect 9697 2148 9701 2204
rect 9637 2144 9701 2148
rect 9717 2204 9781 2208
rect 9717 2148 9721 2204
rect 9721 2148 9777 2204
rect 9777 2148 9781 2204
rect 9717 2144 9781 2148
<< metal4 >>
rect 3075 14720 3395 14736
rect 3075 14656 3083 14720
rect 3147 14656 3163 14720
rect 3227 14656 3243 14720
rect 3307 14656 3323 14720
rect 3387 14656 3395 14720
rect 3075 13632 3395 14656
rect 3075 13568 3083 13632
rect 3147 13568 3163 13632
rect 3227 13568 3243 13632
rect 3307 13568 3323 13632
rect 3387 13568 3395 13632
rect 3075 12672 3395 13568
rect 3075 12544 3117 12672
rect 3353 12544 3395 12672
rect 3075 12480 3083 12544
rect 3387 12480 3395 12544
rect 3075 12436 3117 12480
rect 3353 12436 3395 12480
rect 3075 11456 3395 12436
rect 3075 11392 3083 11456
rect 3147 11392 3163 11456
rect 3227 11392 3243 11456
rect 3307 11392 3323 11456
rect 3387 11392 3395 11456
rect 3075 10368 3395 11392
rect 3075 10304 3083 10368
rect 3147 10304 3163 10368
rect 3227 10304 3243 10368
rect 3307 10304 3323 10368
rect 3387 10304 3395 10368
rect 3075 9280 3395 10304
rect 3075 9216 3083 9280
rect 3147 9216 3163 9280
rect 3227 9216 3243 9280
rect 3307 9216 3323 9280
rect 3387 9216 3395 9280
rect 3075 8502 3395 9216
rect 3075 8266 3117 8502
rect 3353 8266 3395 8502
rect 3075 8192 3395 8266
rect 3075 8128 3083 8192
rect 3147 8128 3163 8192
rect 3227 8128 3243 8192
rect 3307 8128 3323 8192
rect 3387 8128 3395 8192
rect 3075 7104 3395 8128
rect 3075 7040 3083 7104
rect 3147 7040 3163 7104
rect 3227 7040 3243 7104
rect 3307 7040 3323 7104
rect 3387 7040 3395 7104
rect 3075 6016 3395 7040
rect 3075 5952 3083 6016
rect 3147 5952 3163 6016
rect 3227 5952 3243 6016
rect 3307 5952 3323 6016
rect 3387 5952 3395 6016
rect 3075 4928 3395 5952
rect 3075 4864 3083 4928
rect 3147 4864 3163 4928
rect 3227 4864 3243 4928
rect 3307 4864 3323 4928
rect 3387 4864 3395 4928
rect 3075 4331 3395 4864
rect 3075 4095 3117 4331
rect 3353 4095 3395 4331
rect 3075 3840 3395 4095
rect 3075 3776 3083 3840
rect 3147 3776 3163 3840
rect 3227 3776 3243 3840
rect 3307 3776 3323 3840
rect 3387 3776 3395 3840
rect 3075 2752 3395 3776
rect 3075 2688 3083 2752
rect 3147 2688 3163 2752
rect 3227 2688 3243 2752
rect 3307 2688 3323 2752
rect 3387 2688 3395 2752
rect 3075 2128 3395 2688
rect 5206 14176 5526 14736
rect 5206 14112 5214 14176
rect 5278 14112 5294 14176
rect 5358 14112 5374 14176
rect 5438 14112 5454 14176
rect 5518 14112 5526 14176
rect 5206 13088 5526 14112
rect 5206 13024 5214 13088
rect 5278 13024 5294 13088
rect 5358 13024 5374 13088
rect 5438 13024 5454 13088
rect 5518 13024 5526 13088
rect 5206 12000 5526 13024
rect 5206 11936 5214 12000
rect 5278 11936 5294 12000
rect 5358 11936 5374 12000
rect 5438 11936 5454 12000
rect 5518 11936 5526 12000
rect 5206 10912 5526 11936
rect 5206 10848 5214 10912
rect 5278 10848 5294 10912
rect 5358 10848 5374 10912
rect 5438 10848 5454 10912
rect 5518 10848 5526 10912
rect 5206 10587 5526 10848
rect 5206 10351 5248 10587
rect 5484 10351 5526 10587
rect 5206 9824 5526 10351
rect 5206 9760 5214 9824
rect 5278 9760 5294 9824
rect 5358 9760 5374 9824
rect 5438 9760 5454 9824
rect 5518 9760 5526 9824
rect 5206 8736 5526 9760
rect 5206 8672 5214 8736
rect 5278 8672 5294 8736
rect 5358 8672 5374 8736
rect 5438 8672 5454 8736
rect 5518 8672 5526 8736
rect 5206 7648 5526 8672
rect 5206 7584 5214 7648
rect 5278 7584 5294 7648
rect 5358 7584 5374 7648
rect 5438 7584 5454 7648
rect 5518 7584 5526 7648
rect 5206 6560 5526 7584
rect 5206 6496 5214 6560
rect 5278 6496 5294 6560
rect 5358 6496 5374 6560
rect 5438 6496 5454 6560
rect 5518 6496 5526 6560
rect 5206 6416 5526 6496
rect 5206 6180 5248 6416
rect 5484 6180 5526 6416
rect 5206 5472 5526 6180
rect 5206 5408 5214 5472
rect 5278 5408 5294 5472
rect 5358 5408 5374 5472
rect 5438 5408 5454 5472
rect 5518 5408 5526 5472
rect 5206 4384 5526 5408
rect 5206 4320 5214 4384
rect 5278 4320 5294 4384
rect 5358 4320 5374 4384
rect 5438 4320 5454 4384
rect 5518 4320 5526 4384
rect 5206 3296 5526 4320
rect 5206 3232 5214 3296
rect 5278 3232 5294 3296
rect 5358 3232 5374 3296
rect 5438 3232 5454 3296
rect 5518 3232 5526 3296
rect 5206 2208 5526 3232
rect 5206 2144 5214 2208
rect 5278 2144 5294 2208
rect 5358 2144 5374 2208
rect 5438 2144 5454 2208
rect 5518 2144 5526 2208
rect 5206 2128 5526 2144
rect 7338 14720 7658 14736
rect 7338 14656 7346 14720
rect 7410 14656 7426 14720
rect 7490 14656 7506 14720
rect 7570 14656 7586 14720
rect 7650 14656 7658 14720
rect 7338 13632 7658 14656
rect 7338 13568 7346 13632
rect 7410 13568 7426 13632
rect 7490 13568 7506 13632
rect 7570 13568 7586 13632
rect 7650 13568 7658 13632
rect 7338 12672 7658 13568
rect 7338 12544 7380 12672
rect 7616 12544 7658 12672
rect 7338 12480 7346 12544
rect 7650 12480 7658 12544
rect 7338 12436 7380 12480
rect 7616 12436 7658 12480
rect 7338 11456 7658 12436
rect 7338 11392 7346 11456
rect 7410 11392 7426 11456
rect 7490 11392 7506 11456
rect 7570 11392 7586 11456
rect 7650 11392 7658 11456
rect 7338 10368 7658 11392
rect 7338 10304 7346 10368
rect 7410 10304 7426 10368
rect 7490 10304 7506 10368
rect 7570 10304 7586 10368
rect 7650 10304 7658 10368
rect 7338 9280 7658 10304
rect 7338 9216 7346 9280
rect 7410 9216 7426 9280
rect 7490 9216 7506 9280
rect 7570 9216 7586 9280
rect 7650 9216 7658 9280
rect 7338 8502 7658 9216
rect 7338 8266 7380 8502
rect 7616 8266 7658 8502
rect 7338 8192 7658 8266
rect 7338 8128 7346 8192
rect 7410 8128 7426 8192
rect 7490 8128 7506 8192
rect 7570 8128 7586 8192
rect 7650 8128 7658 8192
rect 7338 7104 7658 8128
rect 7338 7040 7346 7104
rect 7410 7040 7426 7104
rect 7490 7040 7506 7104
rect 7570 7040 7586 7104
rect 7650 7040 7658 7104
rect 7338 6016 7658 7040
rect 7338 5952 7346 6016
rect 7410 5952 7426 6016
rect 7490 5952 7506 6016
rect 7570 5952 7586 6016
rect 7650 5952 7658 6016
rect 7338 4928 7658 5952
rect 7338 4864 7346 4928
rect 7410 4864 7426 4928
rect 7490 4864 7506 4928
rect 7570 4864 7586 4928
rect 7650 4864 7658 4928
rect 7338 4331 7658 4864
rect 7338 4095 7380 4331
rect 7616 4095 7658 4331
rect 7338 3840 7658 4095
rect 7338 3776 7346 3840
rect 7410 3776 7426 3840
rect 7490 3776 7506 3840
rect 7570 3776 7586 3840
rect 7650 3776 7658 3840
rect 7338 2752 7658 3776
rect 7338 2688 7346 2752
rect 7410 2688 7426 2752
rect 7490 2688 7506 2752
rect 7570 2688 7586 2752
rect 7650 2688 7658 2752
rect 7338 2128 7658 2688
rect 9469 14176 9789 14736
rect 9469 14112 9477 14176
rect 9541 14112 9557 14176
rect 9621 14112 9637 14176
rect 9701 14112 9717 14176
rect 9781 14112 9789 14176
rect 9469 13088 9789 14112
rect 9469 13024 9477 13088
rect 9541 13024 9557 13088
rect 9621 13024 9637 13088
rect 9701 13024 9717 13088
rect 9781 13024 9789 13088
rect 9469 12000 9789 13024
rect 9469 11936 9477 12000
rect 9541 11936 9557 12000
rect 9621 11936 9637 12000
rect 9701 11936 9717 12000
rect 9781 11936 9789 12000
rect 9469 10912 9789 11936
rect 9469 10848 9477 10912
rect 9541 10848 9557 10912
rect 9621 10848 9637 10912
rect 9701 10848 9717 10912
rect 9781 10848 9789 10912
rect 9469 10587 9789 10848
rect 9469 10351 9511 10587
rect 9747 10351 9789 10587
rect 9469 9824 9789 10351
rect 9469 9760 9477 9824
rect 9541 9760 9557 9824
rect 9621 9760 9637 9824
rect 9701 9760 9717 9824
rect 9781 9760 9789 9824
rect 9469 8736 9789 9760
rect 9469 8672 9477 8736
rect 9541 8672 9557 8736
rect 9621 8672 9637 8736
rect 9701 8672 9717 8736
rect 9781 8672 9789 8736
rect 9469 7648 9789 8672
rect 9469 7584 9477 7648
rect 9541 7584 9557 7648
rect 9621 7584 9637 7648
rect 9701 7584 9717 7648
rect 9781 7584 9789 7648
rect 9469 6560 9789 7584
rect 9469 6496 9477 6560
rect 9541 6496 9557 6560
rect 9621 6496 9637 6560
rect 9701 6496 9717 6560
rect 9781 6496 9789 6560
rect 9469 6416 9789 6496
rect 9469 6180 9511 6416
rect 9747 6180 9789 6416
rect 9469 5472 9789 6180
rect 9469 5408 9477 5472
rect 9541 5408 9557 5472
rect 9621 5408 9637 5472
rect 9701 5408 9717 5472
rect 9781 5408 9789 5472
rect 9469 4384 9789 5408
rect 9469 4320 9477 4384
rect 9541 4320 9557 4384
rect 9621 4320 9637 4384
rect 9701 4320 9717 4384
rect 9781 4320 9789 4384
rect 9469 3296 9789 4320
rect 9469 3232 9477 3296
rect 9541 3232 9557 3296
rect 9621 3232 9637 3296
rect 9701 3232 9717 3296
rect 9781 3232 9789 3296
rect 9469 2208 9789 3232
rect 9469 2144 9477 2208
rect 9541 2144 9557 2208
rect 9621 2144 9637 2208
rect 9701 2144 9717 2208
rect 9781 2144 9789 2208
rect 9469 2128 9789 2144
rect 11600 14720 11920 14736
rect 11600 14656 11608 14720
rect 11672 14656 11688 14720
rect 11752 14656 11768 14720
rect 11832 14656 11848 14720
rect 11912 14656 11920 14720
rect 11600 13632 11920 14656
rect 11600 13568 11608 13632
rect 11672 13568 11688 13632
rect 11752 13568 11768 13632
rect 11832 13568 11848 13632
rect 11912 13568 11920 13632
rect 11600 12672 11920 13568
rect 11600 12544 11642 12672
rect 11878 12544 11920 12672
rect 11600 12480 11608 12544
rect 11912 12480 11920 12544
rect 11600 12436 11642 12480
rect 11878 12436 11920 12480
rect 11600 11456 11920 12436
rect 11600 11392 11608 11456
rect 11672 11392 11688 11456
rect 11752 11392 11768 11456
rect 11832 11392 11848 11456
rect 11912 11392 11920 11456
rect 11600 10368 11920 11392
rect 11600 10304 11608 10368
rect 11672 10304 11688 10368
rect 11752 10304 11768 10368
rect 11832 10304 11848 10368
rect 11912 10304 11920 10368
rect 11600 9280 11920 10304
rect 11600 9216 11608 9280
rect 11672 9216 11688 9280
rect 11752 9216 11768 9280
rect 11832 9216 11848 9280
rect 11912 9216 11920 9280
rect 11600 8502 11920 9216
rect 11600 8266 11642 8502
rect 11878 8266 11920 8502
rect 11600 8192 11920 8266
rect 11600 8128 11608 8192
rect 11672 8128 11688 8192
rect 11752 8128 11768 8192
rect 11832 8128 11848 8192
rect 11912 8128 11920 8192
rect 11600 7104 11920 8128
rect 11600 7040 11608 7104
rect 11672 7040 11688 7104
rect 11752 7040 11768 7104
rect 11832 7040 11848 7104
rect 11912 7040 11920 7104
rect 11600 6016 11920 7040
rect 11600 5952 11608 6016
rect 11672 5952 11688 6016
rect 11752 5952 11768 6016
rect 11832 5952 11848 6016
rect 11912 5952 11920 6016
rect 11600 4928 11920 5952
rect 11600 4864 11608 4928
rect 11672 4864 11688 4928
rect 11752 4864 11768 4928
rect 11832 4864 11848 4928
rect 11912 4864 11920 4928
rect 11600 4331 11920 4864
rect 11600 4095 11642 4331
rect 11878 4095 11920 4331
rect 11600 3840 11920 4095
rect 11600 3776 11608 3840
rect 11672 3776 11688 3840
rect 11752 3776 11768 3840
rect 11832 3776 11848 3840
rect 11912 3776 11920 3840
rect 11600 2752 11920 3776
rect 11600 2688 11608 2752
rect 11672 2688 11688 2752
rect 11752 2688 11768 2752
rect 11832 2688 11848 2752
rect 11912 2688 11920 2752
rect 11600 2128 11920 2688
<< via4 >>
rect 3117 12544 3353 12672
rect 3117 12480 3147 12544
rect 3147 12480 3163 12544
rect 3163 12480 3227 12544
rect 3227 12480 3243 12544
rect 3243 12480 3307 12544
rect 3307 12480 3323 12544
rect 3323 12480 3353 12544
rect 3117 12436 3353 12480
rect 3117 8266 3353 8502
rect 3117 4095 3353 4331
rect 5248 10351 5484 10587
rect 5248 6180 5484 6416
rect 7380 12544 7616 12672
rect 7380 12480 7410 12544
rect 7410 12480 7426 12544
rect 7426 12480 7490 12544
rect 7490 12480 7506 12544
rect 7506 12480 7570 12544
rect 7570 12480 7586 12544
rect 7586 12480 7616 12544
rect 7380 12436 7616 12480
rect 7380 8266 7616 8502
rect 7380 4095 7616 4331
rect 9511 10351 9747 10587
rect 9511 6180 9747 6416
rect 11642 12544 11878 12672
rect 11642 12480 11672 12544
rect 11672 12480 11688 12544
rect 11688 12480 11752 12544
rect 11752 12480 11768 12544
rect 11768 12480 11832 12544
rect 11832 12480 11848 12544
rect 11848 12480 11878 12544
rect 11642 12436 11878 12480
rect 11642 8266 11878 8502
rect 11642 4095 11878 4331
<< metal5 >>
rect 1104 12672 13892 12714
rect 1104 12436 3117 12672
rect 3353 12436 7380 12672
rect 7616 12436 11642 12672
rect 11878 12436 13892 12672
rect 1104 12394 13892 12436
rect 1104 10587 13892 10629
rect 1104 10351 5248 10587
rect 5484 10351 9511 10587
rect 9747 10351 13892 10587
rect 1104 10309 13892 10351
rect 1104 8502 13892 8544
rect 1104 8266 3117 8502
rect 3353 8266 7380 8502
rect 7616 8266 11642 8502
rect 11878 8266 13892 8502
rect 1104 8224 13892 8266
rect 1104 6416 13892 6458
rect 1104 6180 5248 6416
rect 5484 6180 9511 6416
rect 9747 6180 13892 6416
rect 1104 6138 13892 6180
rect 1104 4331 13892 4373
rect 1104 4095 3117 4331
rect 3353 4095 7380 4331
rect 7616 4095 11642 4331
rect 11878 4095 13892 4331
rect 1104 4053 13892 4095
use sky130_fd_sc_hd__decap_8  FILLER_0_7 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 1748 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output9 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform -1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1632082664
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 2484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1632082664
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output12
timestamp 1632082664
transform -1 0 3036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1632082664
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1632082664
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41
timestamp 1632082664
transform 1 0 4876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1632082664
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1632082664
transform 1 0 5428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1632082664
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1632082664
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1632082664
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1632082664
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1632082664
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1632082664
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1632082664
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69
timestamp 1632082664
transform 1 0 7452 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1632082664
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output17
timestamp 1632082664
transform -1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1632082664
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_81
timestamp 1632082664
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1632082664
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1632082664
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79
timestamp 1632082664
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_97
timestamp 1632082664
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1632082664
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1632082664
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1632082664
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1632082664
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1632082664
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output11
timestamp 1632082664
transform -1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1632082664
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1632082664
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_117
timestamp 1632082664
transform 1 0 11868 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1632082664
transform -1 0 13248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output6
timestamp 1632082664
transform 1 0 12880 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_125
timestamp 1632082664
transform 1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_125
timestamp 1632082664
transform 1 0 12604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_132
timestamp 1632082664
transform 1 0 13248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_132
timestamp 1632082664
transform 1 0 13248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1632082664
transform -1 0 13892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1632082664
transform -1 0 13892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1632082664
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1632082664
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1632082664
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1632082664
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1632082664
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1632082664
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1632082664
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1632082664
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1632082664
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1632082664
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1632082664
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1632082664
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1632082664
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 1632082664
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_109
timestamp 1632082664
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_121
timestamp 1632082664
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_133
timestamp 1632082664
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1632082664
transform -1 0 13892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_7
timestamp 1632082664
transform 1 0 1748 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output13
timestamp 1632082664
transform -1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1632082664
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_19
timestamp 1632082664
transform 1 0 2852 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_31
timestamp 1632082664
transform 1 0 3956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_43
timestamp 1632082664
transform 1 0 5060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1632082664
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1632082664
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1632082664
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1632082664
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1632082664
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1632082664
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1632082664
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1632082664
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1632082664
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1632082664
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_125
timestamp 1632082664
transform 1 0 12604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_133
timestamp 1632082664
transform 1 0 13340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1632082664
transform -1 0 13892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1632082664
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1632082664
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1632082664
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1632082664
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1632082664
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1632082664
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1632082664
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1632082664
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1632082664
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1632082664
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1632082664
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1632082664
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1632082664
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1632082664
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1632082664
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1632082664
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_133
timestamp 1632082664
transform 1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1632082664
transform -1 0 13892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1632082664
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1632082664
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1632082664
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1632082664
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1632082664
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1632082664
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1632082664
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1632082664
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1632082664
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1632082664
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1632082664
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1632082664
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1632082664
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1632082664
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1632082664
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1632082664
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_125
timestamp 1632082664
transform 1 0 12604 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_133
timestamp 1632082664
transform 1 0 13340 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1632082664
transform -1 0 13892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1632082664
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1632082664
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1632082664
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1632082664
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1632082664
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1632082664
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1632082664
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1632082664
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1632082664
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1632082664
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_48
timestamp 1632082664
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_39
timestamp 1632082664
transform 1 0 4692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1632082664
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _37_ sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform -1 0 5520 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1632082664
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1632082664
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_64
timestamp 1632082664
transform 1 0 6992 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _21_
timestamp 1632082664
transform -1 0 6992 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1632082664
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_75
timestamp 1632082664
transform 1 0 8004 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1632082664
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _29_
timestamp 1632082664
transform 1 0 7360 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_7_89
timestamp 1632082664
transform 1 0 9292 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1632082664
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1632082664
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_81
timestamp 1632082664
transform 1 0 8556 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__and4_1  _34_
timestamp 1632082664
transform 1 0 8648 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _39_
timestamp 1632082664
transform 1 0 8924 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_7_101
timestamp 1632082664
transform 1 0 10396 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_92
timestamp 1632082664
transform 1 0 9568 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_104
timestamp 1632082664
transform 1 0 10672 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1632082664
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1632082664
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 1632082664
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_125
timestamp 1632082664
transform 1 0 12604 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_116
timestamp 1632082664
transform 1 0 11776 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output20
timestamp 1632082664
transform 1 0 12880 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_132
timestamp 1632082664
transform 1 0 13248 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_133
timestamp 1632082664
transform 1 0 13340 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1632082664
transform -1 0 13892 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1632082664
transform -1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1632082664
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1632082664
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1632082664
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1632082664
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1632082664
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1632082664
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1632082664
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1632082664
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1632082664
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1632082664
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1632082664
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1632082664
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1632082664
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1632082664
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1632082664
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1632082664
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_133
timestamp 1632082664
transform 1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1632082664
transform -1 0 13892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1632082664
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1632082664
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1632082664
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1632082664
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_39
timestamp 1632082664
transform 1 0 4692 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _22_
timestamp 1632082664
transform -1 0 5888 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_9_57
timestamp 1632082664
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1632082664
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_63
timestamp 1632082664
transform 1 0 6900 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1632082664
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _31_ sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 6992 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_75
timestamp 1632082664
transform 1 0 8004 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_71
timestamp 1632082664
transform 1 0 7636 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_67
timestamp 1632082664
transform 1 0 7268 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _26_
timestamp 1632082664
transform 1 0 7728 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_83
timestamp 1632082664
transform 1 0 8740 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__and4_1  _33_
timestamp 1632082664
transform 1 0 8924 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_9_92
timestamp 1632082664
transform 1 0 9568 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_104
timestamp 1632082664
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1632082664
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1632082664
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_125
timestamp 1632082664
transform 1 0 12604 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_133
timestamp 1632082664
transform 1 0 13340 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1632082664
transform -1 0 13892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_7
timestamp 1632082664
transform 1 0 1748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output15
timestamp 1632082664
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1632082664
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1632082664
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1632082664
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1632082664
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1632082664
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1632082664
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_53
timestamp 1632082664
transform 1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_61
timestamp 1632082664
transform 1 0 6716 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _16_ sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 6992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_75
timestamp 1632082664
transform 1 0 8004 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_71
timestamp 1632082664
transform 1 0 7636 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_67
timestamp 1632082664
transform 1 0 7268 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _14_
timestamp 1632082664
transform -1 0 8004 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1632082664
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1632082664
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1632082664
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1632082664
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1632082664
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1632082664
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_133
timestamp 1632082664
transform 1 0 13340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1632082664
transform -1 0 13892 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1632082664
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1632082664
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1632082664
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1632082664
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_49
timestamp 1632082664
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_39
timestamp 1632082664
transform 1 0 4692 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _25_
timestamp 1632082664
transform -1 0 5612 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_11_57
timestamp 1632082664
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1632082664
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1632082664
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _13_
timestamp 1632082664
transform 1 0 6900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_66
timestamp 1632082664
transform 1 0 7176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_73
timestamp 1632082664
transform 1 0 7820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _15_
timestamp 1632082664
transform 1 0 7544 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _17_
timestamp 1632082664
transform 1 0 8188 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_87
timestamp 1632082664
transform 1 0 9108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_80
timestamp 1632082664
transform 1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _19_
timestamp 1632082664
transform 1 0 8832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_99
timestamp 1632082664
transform 1 0 10212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1632082664
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1632082664
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1632082664
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_125
timestamp 1632082664
transform 1 0 12604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_133
timestamp 1632082664
transform 1 0 13340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1632082664
transform -1 0 13892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1632082664
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1632082664
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1632082664
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1632082664
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1632082664
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1632082664
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1632082664
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_53
timestamp 1632082664
transform 1 0 5980 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_61
timestamp 1632082664
transform 1 0 6716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _18_
timestamp 1632082664
transform 1 0 6992 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_74
timestamp 1632082664
transform 1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_67
timestamp 1632082664
transform 1 0 7268 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _12_
timestamp 1632082664
transform -1 0 7912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1632082664
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1632082664
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1632082664
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_98
timestamp 1632082664
transform 1 0 10120 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _23_
timestamp 1632082664
transform 1 0 9476 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_12_110
timestamp 1632082664
transform 1 0 11224 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_122
timestamp 1632082664
transform 1 0 12328 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_134
timestamp 1632082664
transform 1 0 13432 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1632082664
transform -1 0 13892 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1632082664
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1632082664
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1632082664
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1632082664
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1632082664
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1632082664
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1632082664
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1632082664
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1632082664
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1632082664
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_49
timestamp 1632082664
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_41
timestamp 1632082664
transform 1 0 4876 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_49
timestamp 1632082664
transform 1 0 5612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_39
timestamp 1632082664
transform 1 0 4692 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _30_
timestamp 1632082664
transform -1 0 5612 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _35_
timestamp 1632082664
transform -1 0 5612 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1632082664
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_60
timestamp 1632082664
transform 1 0 6624 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1632082664
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1632082664
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__and4_1  _38_
timestamp 1632082664
transform -1 0 6624 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_14_72
timestamp 1632082664
transform 1 0 7728 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_72
timestamp 1632082664
transform 1 0 7728 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _24_
timestamp 1632082664
transform 1 0 7452 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _28_
timestamp 1632082664
transform 1 0 8096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_79
timestamp 1632082664
transform 1 0 8372 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1632082664
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__and4_1  _20_
timestamp 1632082664
transform 1 0 8924 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_13_91
timestamp 1632082664
transform 1 0 9476 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_92
timestamp 1632082664
transform 1 0 9568 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_103
timestamp 1632082664
transform 1 0 10580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1632082664
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_104
timestamp 1632082664
transform 1 0 10672 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1632082664
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1632082664
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_128
timestamp 1632082664
transform 1 0 12880 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_116
timestamp 1632082664
transform 1 0 11776 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output14
timestamp 1632082664
transform 1 0 12880 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_125
timestamp 1632082664
transform 1 0 12604 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_132
timestamp 1632082664
transform 1 0 13248 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1632082664
transform -1 0 13892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1632082664
transform -1 0 13892 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1632082664
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1632082664
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1632082664
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1632082664
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_39
timestamp 1632082664
transform 1 0 4692 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _32_
timestamp 1632082664
transform -1 0 5888 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1632082664
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_61
timestamp 1632082664
transform 1 0 6716 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1632082664
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1632082664
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _36_
timestamp 1632082664
transform 1 0 6808 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_15_69
timestamp 1632082664
transform 1 0 7452 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_77
timestamp 1632082664
transform 1 0 8188 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1632082664
transform 1 0 9016 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _27_
timestamp 1632082664
transform 1 0 8372 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 1632082664
transform 1 0 10120 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1632082664
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1632082664
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1632082664
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_125
timestamp 1632082664
transform 1 0 12604 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_133
timestamp 1632082664
transform 1 0 13340 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1632082664
transform -1 0 13892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1632082664
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1632082664
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1632082664
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1632082664
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1632082664
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1632082664
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1632082664
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1632082664
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1632082664
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1632082664
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1632082664
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1632082664
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1632082664
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1632082664
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1632082664
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1632082664
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_133
timestamp 1632082664
transform 1 0 13340 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1632082664
transform -1 0 13892 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1632082664
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1632082664
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1632082664
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1632082664
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1632082664
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1632082664
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1632082664
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1632082664
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1632082664
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1632082664
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1632082664
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1632082664
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1632082664
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1632082664
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1632082664
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1632082664
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_125
timestamp 1632082664
transform 1 0 12604 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_133
timestamp 1632082664
transform 1 0 13340 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1632082664
transform -1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_7
timestamp 1632082664
transform 1 0 1748 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output18
timestamp 1632082664
transform -1 0 1748 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1632082664
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_19
timestamp 1632082664
transform 1 0 2852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1632082664
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1632082664
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1632082664
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1632082664
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1632082664
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1632082664
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1632082664
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1632082664
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1632082664
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1632082664
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1632082664
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1632082664
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1632082664
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_133
timestamp 1632082664
transform 1 0 13340 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1632082664
transform -1 0 13892 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1632082664
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1632082664
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1632082664
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1632082664
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1632082664
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1632082664
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1632082664
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1632082664
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1632082664
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1632082664
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1632082664
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1632082664
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1632082664
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1632082664
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1632082664
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1632082664
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1632082664
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1632082664
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1632082664
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1632082664
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1632082664
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1632082664
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1632082664
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1632082664
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1632082664
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1632082664
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1632082664
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1632082664
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1632082664
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1632082664
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1632082664
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_125
timestamp 1632082664
transform 1 0 12604 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_121
timestamp 1632082664
transform 1 0 12236 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output5
timestamp 1632082664
transform 1 0 12880 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_127
timestamp 1632082664
transform 1 0 12788 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_132
timestamp 1632082664
transform 1 0 13248 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_133
timestamp 1632082664
transform 1 0 13340 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1632082664
transform -1 0 13892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1632082664
transform -1 0 13892 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1632082664
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1632082664
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1632082664
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1632082664
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1632082664
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1632082664
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1632082664
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1632082664
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1632082664
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1632082664
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1632082664
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1632082664
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1632082664
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1632082664
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1632082664
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1632082664
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_125
timestamp 1632082664
transform 1 0 12604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_133
timestamp 1632082664
transform 1 0 13340 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1632082664
transform -1 0 13892 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output19
timestamp 1632082664
transform -1 0 2484 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output7
timestamp 1632082664
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_7
timestamp 1632082664
transform 1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1632082664
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1632082664
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_29
timestamp 1632082664
transform 1 0 3772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1632082664
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output10
timestamp 1632082664
transform -1 0 4692 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1632082664
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_39
timestamp 1632082664
transform 1 0 4692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_51
timestamp 1632082664
transform 1 0 5796 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_57
timestamp 1632082664
transform 1 0 6348 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1632082664
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_55
timestamp 1632082664
transform 1 0 6164 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_69
timestamp 1632082664
transform 1 0 7452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output8
timestamp 1632082664
transform -1 0 7452 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1632082664
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1632082664
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1632082664
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1632082664
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1632082664
transform -1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_113
timestamp 1632082664
transform 1 0 11500 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1632082664
transform 1 0 11408 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_109
timestamp 1632082664
transform 1 0 11132 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1632082664
transform -1 0 13248 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output16
timestamp 1632082664
transform 1 0 12144 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_119
timestamp 1632082664
transform 1 0 12052 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1632082664
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_132
timestamp 1632082664
transform 1 0 13248 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1632082664
transform -1 0 13892 0 1 14144
box -38 -48 314 592
<< labels >>
rlabel metal5 s 1104 6138 13892 6458 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 4053 13892 4373 6 VPWR
port 1 nsew power input
rlabel metal2 s 14922 16364 14978 17164 6 addr[1]
port 3 nsew signal input
rlabel metal2 s 9586 16364 9642 17164 6 addr[2]
port 4 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 addr[3]
port 5 nsew signal input
rlabel metal3 s 14220 13064 15020 13184 6 fet_on[0]
port 6 nsew signal tristate
rlabel metal2 s 13266 0 13322 800 6 fet_on[10]
port 7 nsew signal tristate
rlabel metal3 s 0 15512 800 15632 6 fet_on[11]
port 8 nsew signal tristate
rlabel metal2 s 7010 16364 7066 17164 6 fet_on[12]
port 9 nsew signal tristate
rlabel metal2 s 18 0 74 800 6 fet_on[13]
port 10 nsew signal tristate
rlabel metal2 s 4250 16364 4306 17164 6 fet_on[14]
port 11 nsew signal tristate
rlabel metal2 s 10690 0 10746 800 6 fet_on[15]
port 12 nsew signal tristate
rlabel metal2 s 2594 0 2650 800 6 fet_on[1]
port 13 nsew signal tristate
rlabel metal3 s 0 3816 800 3936 6 fet_on[2]
port 14 nsew signal tristate
rlabel metal3 s 14220 9256 15020 9376 6 fet_on[3]
port 15 nsew signal tristate
rlabel metal3 s 0 7624 800 7744 6 fet_on[4]
port 16 nsew signal tristate
rlabel metal2 s 12346 16364 12402 17164 6 fet_on[5]
port 17 nsew signal tristate
rlabel metal2 s 7930 0 7986 800 6 fet_on[6]
port 18 nsew signal tristate
rlabel metal3 s 0 11704 800 11824 6 fet_on[7]
port 19 nsew signal tristate
rlabel metal2 s 1674 16364 1730 17164 6 fet_on[8]
port 20 nsew signal tristate
rlabel metal3 s 14220 5176 15020 5296 6 fet_on[9]
port 21 nsew signal tristate
rlabel space 13076 1392 13136 1462 1 'addr_0'
<< properties >>
string FIXED_BBOX 0 0 15020 17164
<< end >>
