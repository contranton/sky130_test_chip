* NGSPICE file created from shift_reg.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

.subckt shift_reg VGND VPWR clk din out_window[0] out_window[1] out_window[2] out_window[3]
XFILLER_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0367_ _1088_/CLK _0367_/D VGND VGND VPWR VPWR _0368_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_39_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0298_ _0316_/CLK _0298_/D VGND VGND VPWR VPWR _0299_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_54_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1270_ _1302_/CLK _1270_/D VGND VGND VPWR VPWR _1271_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0221_ _0316_/CLK _0221_/D VGND VGND VPWR VPWR _0222_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0152_ _1162_/CLK _0152_/D VGND VGND VPWR VPWR _0153_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0083_ _1229_/CLK _0083_/D VGND VGND VPWR VPWR _0084_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_32_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0985_ _1017_/CLK _0985_/D VGND VGND VPWR VPWR _0986_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_8_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1606_ _1611_/CLK _1606_/D VGND VGND VPWR VPWR _1607_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1537_ _1578_/CLK _1537_/D VGND VGND VPWR VPWR _1538_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_59_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1468_ _1687_/CLK _1468_/D VGND VGND VPWR VPWR _1469_/D sky130_fd_sc_hd__dfxtp_1
X_0419_ _1077_/CLK _0419_/D VGND VGND VPWR VPWR _0420_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_86_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1399_ _1754_/CLK _1399_/D VGND VGND VPWR VPWR _1400_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0770_ _1827_/CLK _0770_/D VGND VGND VPWR VPWR _0781_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1322_ _1788_/CLK _1322_/D VGND VGND VPWR VPWR _1323_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1253_ _1272_/CLK _1253_/D VGND VGND VPWR VPWR _1254_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0204_ _1178_/CLK _0204_/D VGND VGND VPWR VPWR _0205_/D sky130_fd_sc_hd__dfxtp_1
X_1184_ _1185_/CLK _1184_/D VGND VGND VPWR VPWR _1185_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_37_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0135_ _1162_/CLK _0135_/D VGND VGND VPWR VPWR _0136_/D sky130_fd_sc_hd__dfxtp_1
X_0066_ _1635_/CLK _0066_/D VGND VGND VPWR VPWR _0077_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0968_ _1826_/CLK _0968_/D VGND VGND VPWR VPWR _0979_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_12_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_4_12_0_clk/X sky130_fd_sc_hd__clkbuf_1
X_0899_ _0908_/CLK _0899_/D VGND VGND VPWR VPWR _0900_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1940_ _1956_/CLK _1940_/D VGND VGND VPWR VPWR _1941_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_61_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1871_ _1995_/CLK _1871_/D VGND VGND VPWR VPWR _1872_/D sky130_fd_sc_hd__dfxtp_1
X_0822_ _0831_/CLK _0822_/D VGND VGND VPWR VPWR _0823_/D sky130_fd_sc_hd__dfxtp_1
X_0753_ _0761_/CLK _0753_/D VGND VGND VPWR VPWR _0754_/D sky130_fd_sc_hd__dfxtp_1
X_0684_ _0898_/CLK _0684_/D VGND VGND VPWR VPWR _0685_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_6_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1305_ _1320_/CLK _1305_/D VGND VGND VPWR VPWR _1306_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_84_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1236_ _1244_/CLK _1236_/D VGND VGND VPWR VPWR _1237_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1167_ _1170_/CLK _1167_/D VGND VGND VPWR VPWR _1168_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0118_ _1138_/CLK _0118_/D VGND VGND VPWR VPWR _0119_/D sky130_fd_sc_hd__dfxtp_1
X_1098_ _1103_/CLK _1098_/D VGND VGND VPWR VPWR _1099_/D sky130_fd_sc_hd__dfxtp_1
X_0049_ _1841_/CLK _0049_/D VGND VGND VPWR VPWR _0050_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1021_ _1033_/CLK _1021_/D VGND VGND VPWR VPWR _1022_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1923_ _1936_/CLK _1923_/D VGND VGND VPWR VPWR _1924_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1854_ _1862_/CLK _1854_/D VGND VGND VPWR VPWR _1856_/D sky130_fd_sc_hd__dfxtp_1
X_0805_ _0906_/CLK _0805_/D VGND VGND VPWR VPWR _0806_/D sky130_fd_sc_hd__dfxtp_1
X_1785_ _1788_/CLK _1785_/D VGND VGND VPWR VPWR _1786_/D sky130_fd_sc_hd__dfxtp_1
X_0736_ _1147_/CLK _0736_/D VGND VGND VPWR VPWR _0738_/D sky130_fd_sc_hd__dfxtp_1
X_0667_ _0916_/CLK _0667_/D VGND VGND VPWR VPWR _0668_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0598_ _0632_/CLK _0598_/D VGND VGND VPWR VPWR _0599_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_69_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1219_ _1228_/CLK _1219_/D VGND VGND VPWR VPWR _1220_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1570_ _1592_/CLK _1570_/D VGND VGND VPWR VPWR _1571_/D sky130_fd_sc_hd__dfxtp_1
X_0521_ _0529_/CLK _0521_/D VGND VGND VPWR VPWR _0522_/D sky130_fd_sc_hd__dfxtp_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0452_ _0585_/CLK _0452_/D VGND VGND VPWR VPWR _0453_/D sky130_fd_sc_hd__dfxtp_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0383_ _1103_/CLK _0383_/D VGND VGND VPWR VPWR _0384_/D sky130_fd_sc_hd__dfxtp_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1004_ _1010_/CLK _1004_/D VGND VGND VPWR VPWR _1005_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_22_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1906_ _1936_/CLK _1906_/D VGND VGND VPWR VPWR _1907_/D sky130_fd_sc_hd__dfxtp_1
X_1837_ _1846_/CLK _1837_/D VGND VGND VPWR VPWR _1838_/D sky130_fd_sc_hd__dfxtp_1
X_1768_ _1772_/CLK _1768_/D VGND VGND VPWR VPWR _1769_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_104_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1699_ _1710_/CLK _1699_/D VGND VGND VPWR VPWR _1700_/D sky130_fd_sc_hd__dfxtp_1
X_0719_ _0793_/CLK _0719_/D VGND VGND VPWR VPWR _0720_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_106_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_114_clk clkbuf_4_1_0_clk/X VGND VGND VPWR VPWR _1747_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_105_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _1862_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1622_ _1673_/CLK _1622_/D VGND VGND VPWR VPWR _1623_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1553_ _1592_/CLK _1553_/D VGND VGND VPWR VPWR _1554_/D sky130_fd_sc_hd__dfxtp_1
X_0504_ _0508_/CLK _0504_/D VGND VGND VPWR VPWR _0505_/D sky130_fd_sc_hd__dfxtp_1
X_1484_ _1965_/CLK _1484_/D VGND VGND VPWR VPWR _1485_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0435_ _0973_/CLK _0435_/D VGND VGND VPWR VPWR _0436_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_86_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0366_ _1112_/CLK _0366_/D VGND VGND VPWR VPWR _0367_/D sky130_fd_sc_hd__dfxtp_1
X_0297_ _0539_/CLK _0297_/D VGND VGND VPWR VPWR _0308_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0220_ _1594_/CLK _0220_/D VGND VGND VPWR VPWR _0231_/D sky130_fd_sc_hd__dfxtp_1
X_0151_ _1170_/CLK _0151_/D VGND VGND VPWR VPWR _0152_/D sky130_fd_sc_hd__dfxtp_1
X_0082_ _1229_/CLK _0082_/D VGND VGND VPWR VPWR _0083_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0984_ _1039_/CLK _0984_/D VGND VGND VPWR VPWR _0985_/D sky130_fd_sc_hd__dfxtp_1
X_1605_ _1611_/CLK _1605_/D VGND VGND VPWR VPWR _1606_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1536_ _1578_/CLK _1536_/D VGND VGND VPWR VPWR _1537_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1467_ _1726_/CLK _1467_/D VGND VGND VPWR VPWR _1468_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1398_ _1754_/CLK _1398_/D VGND VGND VPWR VPWR _1399_/D sky130_fd_sc_hd__dfxtp_1
X_0418_ _0539_/CLK _0418_/D VGND VGND VPWR VPWR _0429_/D sky130_fd_sc_hd__dfxtp_1
X_0349_ _1181_/CLK _0349_/D VGND VGND VPWR VPWR _0350_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_82_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1321_ _1788_/CLK _1321_/D VGND VGND VPWR VPWR _1322_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1252_ _1272_/CLK _1252_/D VGND VGND VPWR VPWR _1253_/D sky130_fd_sc_hd__dfxtp_1
X_0203_ _1178_/CLK _0203_/D VGND VGND VPWR VPWR _0204_/D sky130_fd_sc_hd__dfxtp_1
X_1183_ _1578_/CLK _1183_/D VGND VGND VPWR VPWR _1183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0134_ _1228_/CLK _0134_/D VGND VGND VPWR VPWR _0135_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0065_ _1185_/CLK _0065_/D VGND VGND VPWR VPWR _0067_/D sky130_fd_sc_hd__dfxtp_1
X_0967_ _1039_/CLK _0967_/D VGND VGND VPWR VPWR _0969_/D sky130_fd_sc_hd__dfxtp_1
X_0898_ _0898_/CLK _0898_/D VGND VGND VPWR VPWR _0899_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1519_ _1587_/CLK _1519_/D VGND VGND VPWR VPWR _1520_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_94_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _1600_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_85_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _1936_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1870_ _1997_/CLK _1870_/D VGND VGND VPWR VPWR _1871_/D sky130_fd_sc_hd__dfxtp_1
X_0821_ _0831_/CLK _0821_/D VGND VGND VPWR VPWR _0822_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0752_ _0761_/CLK _0752_/D VGND VGND VPWR VPWR _0753_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_6_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0683_ _0898_/CLK _0683_/D VGND VGND VPWR VPWR _0684_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1304_ _1320_/CLK _1304_/D VGND VGND VPWR VPWR _1305_/D sky130_fd_sc_hd__dfxtp_1
X_1235_ _1302_/CLK _1235_/D VGND VGND VPWR VPWR _1236_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_76_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _1858_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1166_ _1841_/CLK _1166_/D VGND VGND VPWR VPWR _1177_/D sky130_fd_sc_hd__dfxtp_1
X_0117_ _0743_/CLK _0117_/D VGND VGND VPWR VPWR _0118_/D sky130_fd_sc_hd__dfxtp_1
X_1097_ _1104_/CLK _1097_/D VGND VGND VPWR VPWR _1098_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0048_ _0169_/CLK _0048_/D VGND VGND VPWR VPWR _0049_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_69_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_67_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _0280_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_58_clk clkbuf_4_15_0_clk/X VGND VGND VPWR VPWR _0573_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_11_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_4_11_0_clk/X sky130_fd_sc_hd__clkbuf_1
X_1020_ _1039_/CLK _1020_/D VGND VGND VPWR VPWR _1021_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_34_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1922_ _1936_/CLK _1922_/D VGND VGND VPWR VPWR _1923_/D sky130_fd_sc_hd__dfxtp_1
X_1853_ _1997_/CLK _1853_/D VGND VGND VPWR VPWR _1854_/D sky130_fd_sc_hd__dfxtp_1
X_0804_ _0906_/CLK _0804_/D VGND VGND VPWR VPWR _0805_/D sky130_fd_sc_hd__dfxtp_1
X_1784_ _1788_/CLK _1784_/D VGND VGND VPWR VPWR _1785_/D sky130_fd_sc_hd__dfxtp_1
X_0735_ _0743_/CLK _0735_/D VGND VGND VPWR VPWR _0736_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_103_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0666_ _0908_/CLK _0666_/D VGND VGND VPWR VPWR _0667_/D sky130_fd_sc_hd__dfxtp_1
X_0597_ _0610_/CLK _0597_/D VGND VGND VPWR VPWR _0598_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_49_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _0966_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1218_ _1228_/CLK _1218_/D VGND VGND VPWR VPWR _1219_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1149_ _1162_/CLK _1149_/D VGND VGND VPWR VPWR _1150_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_21_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0520_ _0529_/CLK _0520_/D VGND VGND VPWR VPWR _0521_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_6_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0451_ _1985_/CLK _0451_/D VGND VGND VPWR VPWR _0462_/D sky130_fd_sc_hd__dfxtp_1
X_0382_ _1104_/CLK _0382_/D VGND VGND VPWR VPWR _0383_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1003_ _1010_/CLK _1003_/D VGND VGND VPWR VPWR _1004_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_50_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1905_ _1907_/CLK _1905_/D VGND VGND VPWR VPWR _1906_/D sky130_fd_sc_hd__dfxtp_1
X_1836_ _1846_/CLK _1836_/D VGND VGND VPWR VPWR _1837_/D sky130_fd_sc_hd__dfxtp_1
X_1767_ _1833_/CLK _1767_/D VGND VGND VPWR VPWR _1778_/D sky130_fd_sc_hd__dfxtp_1
X_0718_ _0793_/CLK _0718_/D VGND VGND VPWR VPWR _0719_/D sky130_fd_sc_hd__dfxtp_1
X_1698_ _1710_/CLK _1698_/D VGND VGND VPWR VPWR _1699_/D sky130_fd_sc_hd__dfxtp_1
X_0649_ _1649_/CLK _0649_/D VGND VGND VPWR VPWR _0660_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_97_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1621_ _1673_/CLK _1621_/D VGND VGND VPWR VPWR _1622_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1552_ _1918_/CLK _1552_/D VGND VGND VPWR VPWR _1553_/D sky130_fd_sc_hd__dfxtp_1
X_0503_ _0529_/CLK _0503_/D VGND VGND VPWR VPWR _0504_/D sky130_fd_sc_hd__dfxtp_1
X_1483_ _1987_/CLK _1483_/D VGND VGND VPWR VPWR _1484_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0434_ _0973_/CLK _0434_/D VGND VGND VPWR VPWR _0435_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_100_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0365_ _1088_/CLK _0365_/D VGND VGND VPWR VPWR _0366_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0296_ _0316_/CLK _0296_/D VGND VGND VPWR VPWR _0298_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_82_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1819_ _1826_/CLK _1819_/D VGND VGND VPWR VPWR _1820_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0150_ _1170_/CLK _0150_/D VGND VGND VPWR VPWR _0151_/D sky130_fd_sc_hd__dfxtp_1
X_0081_ _1228_/CLK _0081_/D VGND VGND VPWR VPWR _0082_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_17_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0983_ _1039_/CLK _0983_/D VGND VGND VPWR VPWR _0984_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1604_ _1604_/CLK _1604_/D VGND VGND VPWR VPWR _1605_/D sky130_fd_sc_hd__dfxtp_1
X_1535_ _1578_/CLK _1535_/D VGND VGND VPWR VPWR _1536_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1466_ _1687_/CLK _1466_/D VGND VGND VPWR VPWR _1467_/D sky130_fd_sc_hd__dfxtp_1
X_0417_ _1077_/CLK _0417_/D VGND VGND VPWR VPWR _0419_/D sky130_fd_sc_hd__dfxtp_1
X_1397_ _1754_/CLK _1397_/D VGND VGND VPWR VPWR _1398_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0348_ _1181_/CLK _0348_/D VGND VGND VPWR VPWR _0349_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_94_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0279_ _1980_/CLK _0279_/D VGND VGND VPWR VPWR _0280_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_70_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1320_ _1320_/CLK _1320_/D VGND VGND VPWR VPWR _1321_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1251_ _1272_/CLK _1251_/D VGND VGND VPWR VPWR _1252_/D sky130_fd_sc_hd__dfxtp_1
X_1182_ _1182_/CLK _1182_/D VGND VGND VPWR VPWR _1183_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0202_ _1178_/CLK _0202_/D VGND VGND VPWR VPWR _0203_/D sky130_fd_sc_hd__dfxtp_1
X_0133_ _1138_/CLK _0133_/D VGND VGND VPWR VPWR _0134_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_91_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0064_ _1185_/CLK _0064_/D VGND VGND VPWR VPWR _0065_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0966_ _0966_/CLK _0966_/D VGND VGND VPWR VPWR _0967_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_9_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0897_ _0908_/CLK _0897_/D VGND VGND VPWR VPWR _0898_/D sky130_fd_sc_hd__dfxtp_1
X_1518_ _1604_/CLK _1518_/D VGND VGND VPWR VPWR _1519_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1449_ _1695_/CLK _1449_/D VGND VGND VPWR VPWR _1450_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_59_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0820_ _0831_/CLK _0820_/D VGND VGND VPWR VPWR _0821_/D sky130_fd_sc_hd__dfxtp_1
X_0751_ _0761_/CLK _0751_/D VGND VGND VPWR VPWR _0752_/D sky130_fd_sc_hd__dfxtp_1
X_0682_ _1862_/CLK _0682_/D VGND VGND VPWR VPWR _0693_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1303_ _1336_/CLK _1303_/D VGND VGND VPWR VPWR _1304_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_96_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1234_ _1302_/CLK _1234_/D VGND VGND VPWR VPWR _1235_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_77_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1165_ _1170_/CLK _1165_/D VGND VGND VPWR VPWR _1167_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1096_ _1104_/CLK _1096_/D VGND VGND VPWR VPWR _1097_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_18_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0116_ _0743_/CLK _0116_/D VGND VGND VPWR VPWR _0117_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0047_ _1841_/CLK _0047_/D VGND VGND VPWR VPWR _0048_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0949_ _0953_/CLK _0949_/D VGND VGND VPWR VPWR _0950_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1921_ _1965_/CLK _1921_/D VGND VGND VPWR VPWR _1932_/D sky130_fd_sc_hd__dfxtp_1
X_1852_ _1862_/CLK _1852_/D VGND VGND VPWR VPWR _1853_/D sky130_fd_sc_hd__dfxtp_1
X_0803_ _1827_/CLK _0803_/D VGND VGND VPWR VPWR _0814_/D sky130_fd_sc_hd__dfxtp_1
X_1783_ _1783_/CLK _1783_/D VGND VGND VPWR VPWR _1784_/D sky130_fd_sc_hd__dfxtp_1
X_0734_ _1147_/CLK _0734_/D VGND VGND VPWR VPWR _0735_/D sky130_fd_sc_hd__dfxtp_1
X_0665_ _0908_/CLK _0665_/D VGND VGND VPWR VPWR _0666_/D sky130_fd_sc_hd__dfxtp_1
X_0596_ _0610_/CLK _0596_/D VGND VGND VPWR VPWR _0597_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_97_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1217_ _1816_/CLK _1217_/D VGND VGND VPWR VPWR _1218_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_65_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1148_ _1162_/CLK _1148_/D VGND VGND VPWR VPWR _1149_/D sky130_fd_sc_hd__dfxtp_1
X_1079_ _1104_/CLK _1079_/D VGND VGND VPWR VPWR _1080_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0450_ _0585_/CLK _0450_/D VGND VGND VPWR VPWR _0452_/D sky130_fd_sc_hd__dfxtp_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0381_ _0906_/CLK _0381_/D VGND VGND VPWR VPWR _0382_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_79_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1002_ _1010_/CLK _1002_/D VGND VGND VPWR VPWR _1003_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_19_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1904_ _1985_/CLK _1904_/D VGND VGND VPWR VPWR _1905_/D sky130_fd_sc_hd__dfxtp_1
X_1835_ _1846_/CLK _1835_/D VGND VGND VPWR VPWR _1836_/D sky130_fd_sc_hd__dfxtp_1
X_1766_ _1772_/CLK _1766_/D VGND VGND VPWR VPWR _1768_/D sky130_fd_sc_hd__dfxtp_1
X_0717_ _0793_/CLK _0717_/D VGND VGND VPWR VPWR _0718_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_104_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1697_ _1710_/CLK _1697_/D VGND VGND VPWR VPWR _1698_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_106_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0648_ _0919_/CLK _0648_/D VGND VGND VPWR VPWR _0650_/D sky130_fd_sc_hd__dfxtp_1
X_0579_ _0585_/CLK _0579_/D VGND VGND VPWR VPWR _0580_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_85_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_10_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_4_10_0_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1620_ _1965_/CLK _1620_/D VGND VGND VPWR VPWR _1621_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1551_ _1918_/CLK _1551_/D VGND VGND VPWR VPWR _1552_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0502_ _0508_/CLK _0502_/D VGND VGND VPWR VPWR _0503_/D sky130_fd_sc_hd__dfxtp_1
X_1482_ _1965_/CLK _1482_/D VGND VGND VPWR VPWR _1483_/D sky130_fd_sc_hd__dfxtp_1
X_0433_ _0973_/CLK _0433_/D VGND VGND VPWR VPWR _0434_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0364_ _1112_/CLK _0364_/D VGND VGND VPWR VPWR _0365_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_54_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0295_ _0295_/CLK _0295_/D VGND VGND VPWR VPWR _0296_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_82_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1818_ _1841_/CLK _1818_/D VGND VGND VPWR VPWR _1819_/D sky130_fd_sc_hd__dfxtp_1
X_1749_ _1783_/CLK _1749_/D VGND VGND VPWR VPWR _1750_/D sky130_fd_sc_hd__dfxtp_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0080_ _1228_/CLK _0080_/D VGND VGND VPWR VPWR _0081_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0982_ _1017_/CLK _0982_/D VGND VGND VPWR VPWR _0983_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1603_ _1604_/CLK _1603_/D VGND VGND VPWR VPWR _1604_/D sky130_fd_sc_hd__dfxtp_1
X_1534_ _1578_/CLK _1534_/D VGND VGND VPWR VPWR _1535_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_87_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1465_ _1687_/CLK _1465_/D VGND VGND VPWR VPWR _1466_/D sky130_fd_sc_hd__dfxtp_1
X_0416_ _1077_/CLK _0416_/D VGND VGND VPWR VPWR _0417_/D sky130_fd_sc_hd__dfxtp_1
X_1396_ _1754_/CLK _1396_/D VGND VGND VPWR VPWR _1397_/D sky130_fd_sc_hd__dfxtp_1
X_0347_ _1181_/CLK _0347_/D VGND VGND VPWR VPWR _0348_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_103_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0278_ _1980_/CLK _0278_/D VGND VGND VPWR VPWR _0279_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_23_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1250_ _1272_/CLK _1250_/D VGND VGND VPWR VPWR _1251_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0201_ _1178_/CLK _0201_/D VGND VGND VPWR VPWR _0202_/D sky130_fd_sc_hd__dfxtp_1
X_1181_ _1181_/CLK _1181_/D VGND VGND VPWR VPWR _1182_/D sky130_fd_sc_hd__dfxtp_2
X_0132_ _1635_/CLK _0132_/D VGND VGND VPWR VPWR _0143_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_94_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0063_ _1162_/CLK _0063_/D VGND VGND VPWR VPWR _0064_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0965_ _0973_/CLK _0965_/D VGND VGND VPWR VPWR _0966_/D sky130_fd_sc_hd__dfxtp_1
X_0896_ _0898_/CLK _0896_/D VGND VGND VPWR VPWR _0897_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1517_ _1587_/CLK _1517_/D VGND VGND VPWR VPWR _1518_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1448_ _1695_/CLK _1448_/D VGND VGND VPWR VPWR _1449_/D sky130_fd_sc_hd__dfxtp_1
X_1379_ _1764_/CLK _1379_/D VGND VGND VPWR VPWR _1380_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_82_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0750_ _0750_/CLK _0750_/D VGND VGND VPWR VPWR _0751_/D sky130_fd_sc_hd__dfxtp_1
X_0681_ _0898_/CLK _0681_/D VGND VGND VPWR VPWR _0683_/D sky130_fd_sc_hd__dfxtp_1
X_1302_ _1302_/CLK _1302_/D VGND VGND VPWR VPWR _1303_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1233_ _1233_/CLK _1233_/D VGND VGND VPWR VPWR _1234_/D sky130_fd_sc_hd__dfxtp_1
X_1164_ _1170_/CLK _1164_/D VGND VGND VPWR VPWR _1165_/D sky130_fd_sc_hd__dfxtp_1
X_1095_ _1104_/CLK _1095_/D VGND VGND VPWR VPWR _1096_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0115_ _1138_/CLK _0115_/D VGND VGND VPWR VPWR _0116_/D sky130_fd_sc_hd__dfxtp_1
X_0046_ _0169_/CLK _0046_/D VGND VGND VPWR VPWR _0047_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_33_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1997_ _1997_/CLK _1997_/D VGND VGND VPWR VPWR _1997_/Q sky130_fd_sc_hd__dfxtp_1
X_0948_ _0953_/CLK _0948_/D VGND VGND VPWR VPWR _0949_/D sky130_fd_sc_hd__dfxtp_1
X_0879_ _0894_/CLK _0879_/D VGND VGND VPWR VPWR _0881_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_87_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1920_ _1936_/CLK _1920_/D VGND VGND VPWR VPWR _1922_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_42_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1851_ _1862_/CLK _1851_/D VGND VGND VPWR VPWR _1852_/D sky130_fd_sc_hd__dfxtp_1
X_0802_ _0906_/CLK _0802_/D VGND VGND VPWR VPWR _0804_/D sky130_fd_sc_hd__dfxtp_1
X_1782_ _1783_/CLK _1782_/D VGND VGND VPWR VPWR _1783_/D sky130_fd_sc_hd__dfxtp_1
X_0733_ _0793_/CLK _0733_/D VGND VGND VPWR VPWR _0734_/D sky130_fd_sc_hd__dfxtp_1
X_0664_ _0916_/CLK _0664_/D VGND VGND VPWR VPWR _0665_/D sky130_fd_sc_hd__dfxtp_1
X_0595_ _0595_/CLK _0595_/D VGND VGND VPWR VPWR _0596_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_84_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1216_ _1228_/CLK _1216_/D VGND VGND VPWR VPWR _1217_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1147_ _1147_/CLK _1147_/D VGND VGND VPWR VPWR _1148_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1078_ _1826_/CLK _1078_/D VGND VGND VPWR VPWR _1089_/D sky130_fd_sc_hd__dfxtp_1
X_0029_ _1846_/CLK _0029_/D VGND VGND VPWR VPWR _0030_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_117_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _1788_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0380_ _1103_/CLK _0380_/D VGND VGND VPWR VPWR _0381_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1001_ _1686_/CLK _1001_/D VGND VGND VPWR VPWR _1012_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_35_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_108_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _1686_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1903_ _1907_/CLK _1903_/D VGND VGND VPWR VPWR _1904_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1834_ _1862_/CLK _1834_/D VGND VGND VPWR VPWR _1835_/D sky130_fd_sc_hd__dfxtp_1
X_1765_ _1772_/CLK _1765_/D VGND VGND VPWR VPWR _1766_/D sky130_fd_sc_hd__dfxtp_1
X_0716_ _0793_/CLK _0716_/D VGND VGND VPWR VPWR _0717_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1696_ _1710_/CLK _1696_/D VGND VGND VPWR VPWR _1697_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0647_ _0919_/CLK _0647_/D VGND VGND VPWR VPWR _0648_/D sky130_fd_sc_hd__dfxtp_1
X_0578_ _0585_/CLK _0578_/D VGND VGND VPWR VPWR _0579_/D sky130_fd_sc_hd__dfxtp_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1550_ _1918_/CLK _1550_/D VGND VGND VPWR VPWR _1551_/D sky130_fd_sc_hd__dfxtp_1
X_0501_ _0508_/CLK _0501_/D VGND VGND VPWR VPWR _0502_/D sky130_fd_sc_hd__dfxtp_1
X_1481_ _1833_/CLK _1481_/D VGND VGND VPWR VPWR _1482_/D sky130_fd_sc_hd__dfxtp_1
X_0432_ _0966_/CLK _0432_/D VGND VGND VPWR VPWR _0433_/D sky130_fd_sc_hd__dfxtp_1
X_0363_ _1907_/CLK _0363_/D VGND VGND VPWR VPWR _0374_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0294_ _0295_/CLK _0294_/D VGND VGND VPWR VPWR _0295_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_54_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1817_ _1841_/CLK _1817_/D VGND VGND VPWR VPWR _1818_/D sky130_fd_sc_hd__dfxtp_1
X_1748_ _1783_/CLK _1748_/D VGND VGND VPWR VPWR _1749_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_2_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1679_ _1687_/CLK _1679_/D VGND VGND VPWR VPWR _1680_/D sky130_fd_sc_hd__dfxtp_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0981_ _1039_/CLK _0981_/D VGND VGND VPWR VPWR _0982_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_12_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1602_ _1611_/CLK _1602_/D VGND VGND VPWR VPWR _1603_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1533_ _1578_/CLK _1533_/D VGND VGND VPWR VPWR _1534_/D sky130_fd_sc_hd__dfxtp_1
X_1464_ _1687_/CLK _1464_/D VGND VGND VPWR VPWR _1465_/D sky130_fd_sc_hd__dfxtp_1
X_0415_ _1077_/CLK _0415_/D VGND VGND VPWR VPWR _0416_/D sky130_fd_sc_hd__dfxtp_1
X_1395_ _1754_/CLK _1395_/D VGND VGND VPWR VPWR _1396_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0346_ _1181_/CLK _0346_/D VGND VGND VPWR VPWR _0347_/D sky130_fd_sc_hd__dfxtp_1
X_0277_ _1010_/CLK _0277_/D VGND VGND VPWR VPWR _0278_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_35_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_30_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _0874_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_97_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _1987_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_85_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_21_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _0743_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_88_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _1594_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_49_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0200_ _1178_/CLK _0200_/D VGND VGND VPWR VPWR _0201_/D sky130_fd_sc_hd__dfxtp_1
X_1180_ _1180_/CLK _1180_/D VGND VGND VPWR VPWR _1181_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_76_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0131_ _1147_/CLK _0131_/D VGND VGND VPWR VPWR _0133_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0062_ _1185_/CLK _0062_/D VGND VGND VPWR VPWR _0063_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_60_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0964_ _0966_/CLK _0964_/D VGND VGND VPWR VPWR _0965_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_12_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _1185_/CLK sky130_fd_sc_hd__clkbuf_16
X_0895_ _0908_/CLK _0895_/D VGND VGND VPWR VPWR _0896_/D sky130_fd_sc_hd__dfxtp_1
X_1516_ _1604_/CLK _1516_/D VGND VGND VPWR VPWR _1517_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1447_ _1695_/CLK _1447_/D VGND VGND VPWR VPWR _1448_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_79_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _1649_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1378_ _1764_/CLK _1378_/D VGND VGND VPWR VPWR _1379_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_28_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0329_ _1070_/CLK _0329_/D VGND VGND VPWR VPWR _0331_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0680_ _0898_/CLK _0680_/D VGND VGND VPWR VPWR _0681_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_10_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1301_ _1320_/CLK _1301_/D VGND VGND VPWR VPWR _1302_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_1_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _1336_/CLK sky130_fd_sc_hd__clkbuf_16
X_1232_ _1233_/CLK _1232_/D VGND VGND VPWR VPWR _1233_/D sky130_fd_sc_hd__dfxtp_1
X_1163_ _1163_/CLK _1163_/D VGND VGND VPWR VPWR _1164_/D sky130_fd_sc_hd__dfxtp_1
X_1094_ _1104_/CLK _1094_/D VGND VGND VPWR VPWR _1095_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_18_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0114_ _0743_/CLK _0114_/D VGND VGND VPWR VPWR _0115_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0045_ _0169_/CLK _0045_/D VGND VGND VPWR VPWR _0046_/D sky130_fd_sc_hd__dfxtp_1
X_1996_ _1996_/CLK _1996_/D VGND VGND VPWR VPWR _1997_/D sky130_fd_sc_hd__dfxtp_1
X_0947_ _0953_/CLK _0947_/D VGND VGND VPWR VPWR _0948_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0878_ _0894_/CLK _0878_/D VGND VGND VPWR VPWR _0879_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_0_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1850_ _1862_/CLK _1850_/D VGND VGND VPWR VPWR _1851_/D sky130_fd_sc_hd__dfxtp_1
X_0801_ _0813_/CLK _0801_/D VGND VGND VPWR VPWR _0802_/D sky130_fd_sc_hd__dfxtp_1
X_1781_ _1783_/CLK _1781_/D VGND VGND VPWR VPWR _1782_/D sky130_fd_sc_hd__dfxtp_1
X_0732_ _0793_/CLK _0732_/D VGND VGND VPWR VPWR _0733_/D sky130_fd_sc_hd__dfxtp_1
X_0663_ _0908_/CLK _0663_/D VGND VGND VPWR VPWR _0664_/D sky130_fd_sc_hd__dfxtp_1
X_0594_ _1649_/CLK _0594_/D VGND VGND VPWR VPWR _0605_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1215_ _1228_/CLK _1215_/D VGND VGND VPWR VPWR _1216_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1146_ _1162_/CLK _1146_/D VGND VGND VPWR VPWR _1147_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1077_ _1077_/CLK _1077_/D VGND VGND VPWR VPWR _1079_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0028_ _1858_/CLK _0028_/D VGND VGND VPWR VPWR _0029_/D sky130_fd_sc_hd__dfxtp_1
X_1979_ _1991_/CLK _1979_/D VGND VGND VPWR VPWR _1980_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1000_ _1010_/CLK _1000_/D VGND VGND VPWR VPWR _1002_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_19_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1902_ _1985_/CLK _1902_/D VGND VGND VPWR VPWR _1903_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1833_ _1833_/CLK _1833_/D VGND VGND VPWR VPWR _1844_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1764_ _1764_/CLK _1764_/D VGND VGND VPWR VPWR _1765_/D sky130_fd_sc_hd__dfxtp_1
X_0715_ _1665_/CLK _0715_/D VGND VGND VPWR VPWR _0726_/D sky130_fd_sc_hd__dfxtp_1
X_1695_ _1695_/CLK _1695_/D VGND VGND VPWR VPWR _1696_/D sky130_fd_sc_hd__dfxtp_1
X_0646_ _0919_/CLK _0646_/D VGND VGND VPWR VPWR _0647_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_103_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0577_ _0585_/CLK _0577_/D VGND VGND VPWR VPWR _0578_/D sky130_fd_sc_hd__dfxtp_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1129_ _1147_/CLK _1129_/D VGND VGND VPWR VPWR _1130_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0500_ _0508_/CLK _0500_/D VGND VGND VPWR VPWR _0501_/D sky130_fd_sc_hd__dfxtp_1
X_1480_ _1965_/CLK _1480_/D VGND VGND VPWR VPWR _1481_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_97_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0431_ _0973_/CLK _0431_/D VGND VGND VPWR VPWR _0432_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0362_ _1112_/CLK _0362_/D VGND VGND VPWR VPWR _0364_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0293_ _0295_/CLK _0293_/D VGND VGND VPWR VPWR _0294_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_94_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1816_ _1816_/CLK _1816_/D VGND VGND VPWR VPWR _1817_/D sky130_fd_sc_hd__dfxtp_1
X_1747_ _1747_/CLK _1747_/D VGND VGND VPWR VPWR _1748_/D sky130_fd_sc_hd__dfxtp_1
X_1678_ _1687_/CLK _1678_/D VGND VGND VPWR VPWR _1679_/D sky130_fd_sc_hd__dfxtp_1
X_0629_ _0632_/CLK _0629_/D VGND VGND VPWR VPWR _0630_/D sky130_fd_sc_hd__dfxtp_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0980_ _1039_/CLK _0980_/D VGND VGND VPWR VPWR _0981_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1601_ _1611_/CLK _1601_/D VGND VGND VPWR VPWR _1602_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1532_ _1578_/CLK _1532_/D VGND VGND VPWR VPWR _1533_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1463_ _1687_/CLK _1463_/D VGND VGND VPWR VPWR _1464_/D sky130_fd_sc_hd__dfxtp_1
X_0414_ _0622_/CLK _0414_/D VGND VGND VPWR VPWR _0415_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_86_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1394_ _1754_/CLK _1394_/D VGND VGND VPWR VPWR _1395_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0345_ _1181_/CLK _0345_/D VGND VGND VPWR VPWR _0346_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_82_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0276_ _0280_/CLK _0276_/D VGND VGND VPWR VPWR _0277_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0130_ _1138_/CLK _0130_/D VGND VGND VPWR VPWR _0131_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0061_ _1185_/CLK _0061_/D VGND VGND VPWR VPWR _0062_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_17_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0963_ _0966_/CLK _0963_/D VGND VGND VPWR VPWR _0964_/D sky130_fd_sc_hd__dfxtp_1
X_0894_ _0894_/CLK _0894_/D VGND VGND VPWR VPWR _0895_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1515_ _1604_/CLK _1515_/D VGND VGND VPWR VPWR _1516_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1446_ _1695_/CLK _1446_/D VGND VGND VPWR VPWR _1447_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1377_ _1764_/CLK _1377_/D VGND VGND VPWR VPWR _1378_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0328_ _1070_/CLK _0328_/D VGND VGND VPWR VPWR _0329_/D sky130_fd_sc_hd__dfxtp_1
X_0259_ _1973_/CLK _0259_/D VGND VGND VPWR VPWR _0260_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_70_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1300_ _1348_/CLK _1300_/D VGND VGND VPWR VPWR _1301_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_96_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1231_ _1233_/CLK _1231_/D VGND VGND VPWR VPWR _1232_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_77_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1162_ _1162_/CLK _1162_/D VGND VGND VPWR VPWR _1163_/D sky130_fd_sc_hd__dfxtp_1
X_1093_ _1104_/CLK _1093_/D VGND VGND VPWR VPWR _1094_/D sky130_fd_sc_hd__dfxtp_1
X_0113_ _0743_/CLK _0113_/D VGND VGND VPWR VPWR _0114_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0044_ _1635_/CLK _0044_/D VGND VGND VPWR VPWR _0055_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_33_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1995_ _1995_/CLK _1995_/D VGND VGND VPWR VPWR _1996_/D sky130_fd_sc_hd__dfxtp_1
X_0946_ _1686_/CLK _0946_/D VGND VGND VPWR VPWR _0957_/D sky130_fd_sc_hd__dfxtp_1
X_0877_ _0894_/CLK _0877_/D VGND VGND VPWR VPWR _0878_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1429_ _1695_/CLK _1429_/D VGND VGND VPWR VPWR _1430_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0800_ _0906_/CLK _0800_/D VGND VGND VPWR VPWR _0801_/D sky130_fd_sc_hd__dfxtp_1
X_1780_ _1783_/CLK _1780_/D VGND VGND VPWR VPWR _1781_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0731_ _0761_/CLK _0731_/D VGND VGND VPWR VPWR _0732_/D sky130_fd_sc_hd__dfxtp_1
X_0662_ _0908_/CLK _0662_/D VGND VGND VPWR VPWR _0663_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_6_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0593_ _0595_/CLK _0593_/D VGND VGND VPWR VPWR _0595_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1214_ _1228_/CLK _1214_/D VGND VGND VPWR VPWR _1215_/D sky130_fd_sc_hd__dfxtp_1
X_1145_ _1147_/CLK _1145_/D VGND VGND VPWR VPWR _1146_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1076_ _1181_/CLK _1076_/D VGND VGND VPWR VPWR _1077_/D sky130_fd_sc_hd__dfxtp_1
X_0027_ _1862_/CLK _0027_/D VGND VGND VPWR VPWR _0028_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_21_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1978_ _1991_/CLK _1978_/D VGND VGND VPWR VPWR _1979_/D sky130_fd_sc_hd__dfxtp_1
X_0929_ _0932_/CLK _0929_/D VGND VGND VPWR VPWR _0930_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_88_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1901_ _1985_/CLK _1901_/D VGND VGND VPWR VPWR _1902_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1832_ _1862_/CLK _1832_/D VGND VGND VPWR VPWR _1834_/D sky130_fd_sc_hd__dfxtp_1
X_1763_ _1772_/CLK _1763_/D VGND VGND VPWR VPWR _1764_/D sky130_fd_sc_hd__dfxtp_1
X_1694_ _1710_/CLK _1694_/D VGND VGND VPWR VPWR _1695_/D sky130_fd_sc_hd__dfxtp_1
X_0714_ _1127_/CLK _0714_/D VGND VGND VPWR VPWR _0716_/D sky130_fd_sc_hd__dfxtp_1
X_0645_ _0919_/CLK _0645_/D VGND VGND VPWR VPWR _0646_/D sky130_fd_sc_hd__dfxtp_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0576_ _0585_/CLK _0576_/D VGND VGND VPWR VPWR _0577_/D sky130_fd_sc_hd__dfxtp_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1128_ _1147_/CLK _1128_/D VGND VGND VPWR VPWR _1129_/D sky130_fd_sc_hd__dfxtp_1
X_1059_ _1071_/CLK _1059_/D VGND VGND VPWR VPWR _1060_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0430_ _0953_/CLK _0430_/D VGND VGND VPWR VPWR _0431_/D sky130_fd_sc_hd__dfxtp_1
X_0361_ _1112_/CLK _0361_/D VGND VGND VPWR VPWR _0362_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0292_ _0316_/CLK _0292_/D VGND VGND VPWR VPWR _0293_/D sky130_fd_sc_hd__dfxtp_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1815_ _1816_/CLK _1815_/D VGND VGND VPWR VPWR _1816_/D sky130_fd_sc_hd__dfxtp_1
X_1746_ _1747_/CLK _1746_/D VGND VGND VPWR VPWR _1747_/D sky130_fd_sc_hd__dfxtp_1
X_1677_ _1687_/CLK _1677_/D VGND VGND VPWR VPWR _1678_/D sky130_fd_sc_hd__dfxtp_1
X_0628_ _0632_/CLK _0628_/D VGND VGND VPWR VPWR _0629_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_89_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0559_ _0610_/CLK _0559_/D VGND VGND VPWR VPWR _0560_/D sky130_fd_sc_hd__dfxtp_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1600_ _1600_/CLK _1600_/D VGND VGND VPWR VPWR _1601_/D sky130_fd_sc_hd__dfxtp_1
X_1531_ _1578_/CLK _1531_/D VGND VGND VPWR VPWR _1532_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_4_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1462_ _1687_/CLK _1462_/D VGND VGND VPWR VPWR _1463_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_4_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0413_ _0622_/CLK _0413_/D VGND VGND VPWR VPWR _0414_/D sky130_fd_sc_hd__dfxtp_1
X_1393_ _1754_/CLK _1393_/D VGND VGND VPWR VPWR _1394_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_94_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0344_ _1181_/CLK _0344_/D VGND VGND VPWR VPWR _0345_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_82_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0275_ _0539_/CLK _0275_/D VGND VGND VPWR VPWR _0286_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1729_ _1747_/CLK _1729_/D VGND VGND VPWR VPWR _1730_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0060_ _1170_/CLK _0060_/D VGND VGND VPWR VPWR _0061_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_45_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0962_ _0966_/CLK _0962_/D VGND VGND VPWR VPWR _0963_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0893_ _0898_/CLK _0893_/D VGND VGND VPWR VPWR _0894_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1514_ _1604_/CLK _1514_/D VGND VGND VPWR VPWR _1515_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1445_ _1686_/CLK _1445_/D VGND VGND VPWR VPWR _1446_/D sky130_fd_sc_hd__dfxtp_1
X_1376_ _1764_/CLK _1376_/D VGND VGND VPWR VPWR _1377_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0327_ _1070_/CLK _0327_/D VGND VGND VPWR VPWR _0328_/D sky130_fd_sc_hd__dfxtp_1
X_0258_ _1973_/CLK _0258_/D VGND VGND VPWR VPWR _0259_/D sky130_fd_sc_hd__dfxtp_1
X_0189_ _0214_/CLK _0189_/D VGND VGND VPWR VPWR _0190_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_11_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1230_ _1233_/CLK _1230_/D VGND VGND VPWR VPWR _1231_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_49_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1161_ _1162_/CLK _1161_/D VGND VGND VPWR VPWR _1162_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0112_ _0743_/CLK _0112_/D VGND VGND VPWR VPWR _0113_/D sky130_fd_sc_hd__dfxtp_1
X_1092_ _1104_/CLK _1092_/D VGND VGND VPWR VPWR _1093_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0043_ _0169_/CLK _0043_/D VGND VGND VPWR VPWR _0045_/D sky130_fd_sc_hd__dfxtp_1
X_1994_ _1995_/CLK _1994_/D VGND VGND VPWR VPWR _1995_/D sky130_fd_sc_hd__dfxtp_1
X_0945_ _0953_/CLK _0945_/D VGND VGND VPWR VPWR _0947_/D sky130_fd_sc_hd__dfxtp_1
X_0876_ _0894_/CLK _0876_/D VGND VGND VPWR VPWR _0877_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1428_ _1794_/CLK _1428_/D VGND VGND VPWR VPWR _1429_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1359_ _1364_/CLK _1359_/D VGND VGND VPWR VPWR _1360_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0730_ _0793_/CLK _0730_/D VGND VGND VPWR VPWR _0731_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_6_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0661_ _0916_/CLK _0661_/D VGND VGND VPWR VPWR _0662_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_97_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0592_ _0595_/CLK _0592_/D VGND VGND VPWR VPWR _0593_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_97_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1213_ _1228_/CLK _1213_/D VGND VGND VPWR VPWR _1214_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1144_ _1841_/CLK _1144_/D VGND VGND VPWR VPWR _1155_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_53_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1075_ _1181_/CLK _1075_/D VGND VGND VPWR VPWR _1076_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_18_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0026_ _1858_/CLK _0026_/D VGND VGND VPWR VPWR _0027_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1977_ _1991_/CLK _1977_/D VGND VGND VPWR VPWR _1978_/D sky130_fd_sc_hd__dfxtp_1
X_0928_ _0932_/CLK _0928_/D VGND VGND VPWR VPWR _0929_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0859_ _0864_/CLK _0859_/D VGND VGND VPWR VPWR _0860_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_88_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1900_ _1985_/CLK _1900_/D VGND VGND VPWR VPWR _1901_/D sky130_fd_sc_hd__dfxtp_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1831_ _1846_/CLK _1831_/D VGND VGND VPWR VPWR _1832_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1762_ _1772_/CLK _1762_/D VGND VGND VPWR VPWR _1763_/D sky130_fd_sc_hd__dfxtp_1
X_1693_ _1695_/CLK _1693_/D VGND VGND VPWR VPWR _1694_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_7_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0713_ _0793_/CLK _0713_/D VGND VGND VPWR VPWR _0714_/D sky130_fd_sc_hd__dfxtp_1
X_0644_ _0919_/CLK _0644_/D VGND VGND VPWR VPWR _0645_/D sky130_fd_sc_hd__dfxtp_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0575_ _0585_/CLK _0575_/D VGND VGND VPWR VPWR _0576_/D sky130_fd_sc_hd__dfxtp_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1127_ _1127_/CLK _1127_/D VGND VGND VPWR VPWR _1128_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1058_ _1071_/CLK _1058_/D VGND VGND VPWR VPWR _1059_/D sky130_fd_sc_hd__dfxtp_1
X_0009_ _1996_/CLK _0009_/D VGND VGND VPWR VPWR _0010_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_60_clk clkbuf_4_15_0_clk/X VGND VGND VPWR VPWR _0529_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_21_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _1077_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0360_ _1112_/CLK _0360_/D VGND VGND VPWR VPWR _0361_/D sky130_fd_sc_hd__dfxtp_1
X_0291_ _0295_/CLK _0291_/D VGND VGND VPWR VPWR _0292_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_42_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _1088_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1814_ _1814_/CLK _1814_/D VGND VGND VPWR VPWR _1815_/D sky130_fd_sc_hd__dfxtp_1
X_1745_ _1747_/CLK _1745_/D VGND VGND VPWR VPWR _1746_/D sky130_fd_sc_hd__dfxtp_1
X_1676_ _1687_/CLK _1676_/D VGND VGND VPWR VPWR _1677_/D sky130_fd_sc_hd__dfxtp_1
X_0627_ _1665_/CLK _0627_/D VGND VGND VPWR VPWR _0638_/D sky130_fd_sc_hd__dfxtp_1
X_0558_ _0610_/CLK _0558_/D VGND VGND VPWR VPWR _0559_/D sky130_fd_sc_hd__dfxtp_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0489_ _0998_/CLK _0489_/D VGND VGND VPWR VPWR _0490_/D sky130_fd_sc_hd__dfxtp_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_33_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _0906_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_1_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _0791_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1530_ _1578_/CLK _1530_/D VGND VGND VPWR VPWR _1531_/D sky130_fd_sc_hd__dfxtp_1
X_1461_ _1710_/CLK _1461_/D VGND VGND VPWR VPWR _1462_/D sky130_fd_sc_hd__dfxtp_1
X_0412_ _1077_/CLK _0412_/D VGND VGND VPWR VPWR _0413_/D sky130_fd_sc_hd__dfxtp_1
X_1392_ _1754_/CLK _1392_/D VGND VGND VPWR VPWR _1393_/D sky130_fd_sc_hd__dfxtp_1
X_0343_ _1181_/CLK _0343_/D VGND VGND VPWR VPWR _0344_/D sky130_fd_sc_hd__dfxtp_1
X_0274_ _1010_/CLK _0274_/D VGND VGND VPWR VPWR _0276_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_48_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_15_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _1170_/CLK sky130_fd_sc_hd__clkbuf_16
X_1728_ _1736_/CLK _1728_/D VGND VGND VPWR VPWR _1729_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1659_ _1659_/CLK _1659_/D VGND VGND VPWR VPWR _1660_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_104_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0961_ _0966_/CLK _0961_/D VGND VGND VPWR VPWR _0962_/D sky130_fd_sc_hd__dfxtp_1
X_0892_ _0894_/CLK _0892_/D VGND VGND VPWR VPWR _0893_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1513_ _1587_/CLK _1513_/D VGND VGND VPWR VPWR _1514_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1444_ _1686_/CLK _1444_/D VGND VGND VPWR VPWR _1445_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_4_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _1272_/CLK sky130_fd_sc_hd__clkbuf_16
X_1375_ _1764_/CLK _1375_/D VGND VGND VPWR VPWR _1376_/D sky130_fd_sc_hd__dfxtp_1
X_0326_ _1071_/CLK _0326_/D VGND VGND VPWR VPWR _0327_/D sky130_fd_sc_hd__dfxtp_1
X_0257_ _1973_/CLK _0257_/D VGND VGND VPWR VPWR _0258_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_23_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0188_ _1858_/CLK _0188_/D VGND VGND VPWR VPWR _0189_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_63_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1160_ _1163_/CLK _1160_/D VGND VGND VPWR VPWR _1161_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0111_ _0743_/CLK _0111_/D VGND VGND VPWR VPWR _0112_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1091_ _1104_/CLK _1091_/D VGND VGND VPWR VPWR _1092_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0042_ _1841_/CLK _0042_/D VGND VGND VPWR VPWR _0043_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1993_ _1997_/CLK _1993_/D VGND VGND VPWR VPWR _1994_/D sky130_fd_sc_hd__dfxtp_1
X_0944_ _0953_/CLK _0944_/D VGND VGND VPWR VPWR _0945_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0875_ _0894_/CLK _0875_/D VGND VGND VPWR VPWR _0876_/D sky130_fd_sc_hd__dfxtp_1
X_1427_ _1794_/CLK _1427_/D VGND VGND VPWR VPWR _1428_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1358_ _1364_/CLK _1358_/D VGND VGND VPWR VPWR _1359_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1289_ _1348_/CLK _1289_/D VGND VGND VPWR VPWR _1290_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_55_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0309_ _1046_/CLK _0309_/D VGND VGND VPWR VPWR _0310_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0660_ _1649_/CLK _0660_/D VGND VGND VPWR VPWR _0671_/D sky130_fd_sc_hd__dfxtp_1
X_0591_ _0595_/CLK _0591_/D VGND VGND VPWR VPWR _0592_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_97_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1212_ _1233_/CLK _1212_/D VGND VGND VPWR VPWR _1213_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1143_ _1162_/CLK _1143_/D VGND VGND VPWR VPWR _1145_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_65_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1074_ _1181_/CLK _1074_/D VGND VGND VPWR VPWR _1075_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0025_ _1858_/CLK _0025_/D VGND VGND VPWR VPWR _0026_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_60_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1976_ _1987_/CLK _1976_/D VGND VGND VPWR VPWR _1987_/D sky130_fd_sc_hd__dfxtp_1
X_0927_ _1077_/CLK _0927_/D VGND VGND VPWR VPWR _0928_/D sky130_fd_sc_hd__dfxtp_1
X_0858_ _1665_/CLK _0858_/D VGND VGND VPWR VPWR _0869_/D sky130_fd_sc_hd__dfxtp_1
X_0789_ _0791_/CLK _0789_/D VGND VGND VPWR VPWR _0790_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1830_ _1862_/CLK _1830_/D VGND VGND VPWR VPWR _1831_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1761_ _1772_/CLK _1761_/D VGND VGND VPWR VPWR _1762_/D sky130_fd_sc_hd__dfxtp_1
X_0712_ _0793_/CLK _0712_/D VGND VGND VPWR VPWR _0713_/D sky130_fd_sc_hd__dfxtp_1
X_1692_ _1695_/CLK _1692_/D VGND VGND VPWR VPWR _1693_/D sky130_fd_sc_hd__dfxtp_1
X_0643_ _0919_/CLK _0643_/D VGND VGND VPWR VPWR _0644_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_7_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0574_ _0585_/CLK _0574_/D VGND VGND VPWR VPWR _0575_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_97_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1126_ _1127_/CLK _1126_/D VGND VGND VPWR VPWR _1127_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_38_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1057_ _1071_/CLK _1057_/D VGND VGND VPWR VPWR _1058_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0008_ _1997_/CLK _0008_/D VGND VGND VPWR VPWR _0009_/D sky130_fd_sc_hd__dfxtp_1
X_1959_ _1973_/CLK _1959_/D VGND VGND VPWR VPWR _1960_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_102_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0290_ _0295_/CLK _0290_/D VGND VGND VPWR VPWR _0291_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1813_ _1814_/CLK _1813_/D VGND VGND VPWR VPWR _1814_/D sky130_fd_sc_hd__dfxtp_1
X_1744_ _1754_/CLK _1744_/D VGND VGND VPWR VPWR _1745_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1675_ _1687_/CLK _1675_/D VGND VGND VPWR VPWR _1676_/D sky130_fd_sc_hd__dfxtp_1
X_0626_ _0632_/CLK _0626_/D VGND VGND VPWR VPWR _0628_/D sky130_fd_sc_hd__dfxtp_1
X_0557_ _0595_/CLK _0557_/D VGND VGND VPWR VPWR _0558_/D sky130_fd_sc_hd__dfxtp_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0488_ _0998_/CLK _0488_/D VGND VGND VPWR VPWR _0489_/D sky130_fd_sc_hd__dfxtp_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1109_ _1112_/CLK _1109_/D VGND VGND VPWR VPWR _1110_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_22_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1460_ _1687_/CLK _1460_/D VGND VGND VPWR VPWR _1461_/D sky130_fd_sc_hd__dfxtp_1
X_0411_ _0622_/CLK _0411_/D VGND VGND VPWR VPWR _0412_/D sky130_fd_sc_hd__dfxtp_1
X_1391_ _1754_/CLK _1391_/D VGND VGND VPWR VPWR _1392_/D sky130_fd_sc_hd__dfxtp_1
X_0342_ _1181_/CLK _0342_/D VGND VGND VPWR VPWR _0343_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_94_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0273_ _0280_/CLK _0273_/D VGND VGND VPWR VPWR _0274_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1727_ _1736_/CLK _1727_/D VGND VGND VPWR VPWR _1728_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_104_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1658_ _1659_/CLK _1658_/D VGND VGND VPWR VPWR _1659_/D sky130_fd_sc_hd__dfxtp_1
X_0609_ _0610_/CLK _0609_/D VGND VGND VPWR VPWR _0610_/D sky130_fd_sc_hd__dfxtp_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1589_ _1592_/CLK _1589_/D VGND VGND VPWR VPWR _1590_/D sky130_fd_sc_hd__dfxtp_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0960_ _0966_/CLK _0960_/D VGND VGND VPWR VPWR _0961_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_32_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0891_ _1665_/CLK _0891_/D VGND VGND VPWR VPWR _0902_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1512_ _1604_/CLK _1512_/D VGND VGND VPWR VPWR _1513_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1443_ _1686_/CLK _1443_/D VGND VGND VPWR VPWR _1444_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1374_ _1764_/CLK _1374_/D VGND VGND VPWR VPWR _1375_/D sky130_fd_sc_hd__dfxtp_1
X_0325_ _1070_/CLK _0325_/D VGND VGND VPWR VPWR _0326_/D sky130_fd_sc_hd__dfxtp_1
X_0256_ _1980_/CLK _0256_/D VGND VGND VPWR VPWR _0257_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0187_ _1635_/CLK _0187_/D VGND VGND VPWR VPWR _0198_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0110_ _1635_/CLK _0110_/D VGND VGND VPWR VPWR _0121_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1090_ _1104_/CLK _1090_/D VGND VGND VPWR VPWR _1091_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0041_ _1841_/CLK _0041_/D VGND VGND VPWR VPWR _0042_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1992_ _1995_/CLK _1992_/D VGND VGND VPWR VPWR _1993_/D sky130_fd_sc_hd__dfxtp_1
X_0943_ _1077_/CLK _0943_/D VGND VGND VPWR VPWR _0944_/D sky130_fd_sc_hd__dfxtp_1
X_0874_ _0874_/CLK _0874_/D VGND VGND VPWR VPWR _0875_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_102_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1426_ _1794_/CLK _1426_/D VGND VGND VPWR VPWR _1427_/D sky130_fd_sc_hd__dfxtp_1
X_1357_ _1364_/CLK _1357_/D VGND VGND VPWR VPWR _1358_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0308_ _1907_/CLK _0308_/D VGND VGND VPWR VPWR _0319_/D sky130_fd_sc_hd__dfxtp_1
X_1288_ _1348_/CLK _1288_/D VGND VGND VPWR VPWR _1289_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_43_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0239_ _0295_/CLK _0239_/D VGND VGND VPWR VPWR _0240_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_71_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0590_ _0595_/CLK _0590_/D VGND VGND VPWR VPWR _0591_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_97_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1211_ _1233_/CLK _1211_/D VGND VGND VPWR VPWR _1212_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1142_ _1147_/CLK _1142_/D VGND VGND VPWR VPWR _1143_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1073_ _1181_/CLK _1073_/D VGND VGND VPWR VPWR _1074_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_25_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0024_ _1858_/CLK _0024_/D VGND VGND VPWR VPWR _0025_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1975_ _1975_/CLK _1975_/D VGND VGND VPWR VPWR _1977_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0926_ _0932_/CLK _0926_/D VGND VGND VPWR VPWR _0927_/D sky130_fd_sc_hd__dfxtp_1
X_0857_ _0864_/CLK _0857_/D VGND VGND VPWR VPWR _0859_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0788_ _0793_/CLK _0788_/D VGND VGND VPWR VPWR _0789_/D sky130_fd_sc_hd__dfxtp_1
X_1409_ _1747_/CLK _1409_/D VGND VGND VPWR VPWR _1410_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1760_ _1772_/CLK _1760_/D VGND VGND VPWR VPWR _1761_/D sky130_fd_sc_hd__dfxtp_1
X_0711_ _1127_/CLK _0711_/D VGND VGND VPWR VPWR _0712_/D sky130_fd_sc_hd__dfxtp_1
X_1691_ _1695_/CLK _1691_/D VGND VGND VPWR VPWR _1692_/D sky130_fd_sc_hd__dfxtp_1
X_0642_ _0642_/CLK _0642_/D VGND VGND VPWR VPWR _0643_/D sky130_fd_sc_hd__dfxtp_1
X_0573_ _0573_/CLK _0573_/D VGND VGND VPWR VPWR _0574_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_97_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1125_ _1127_/CLK _1125_/D VGND VGND VPWR VPWR _1126_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_93_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1056_ _1826_/CLK _1056_/D VGND VGND VPWR VPWR _1067_/D sky130_fd_sc_hd__dfxtp_1
X_0007_ _1997_/CLK _0007_/D VGND VGND VPWR VPWR _0008_/D sky130_fd_sc_hd__dfxtp_1
X_1958_ _1973_/CLK _1958_/D VGND VGND VPWR VPWR _1959_/D sky130_fd_sc_hd__dfxtp_1
X_0909_ _0919_/CLK _0909_/D VGND VGND VPWR VPWR _0910_/D sky130_fd_sc_hd__dfxtp_1
X_1889_ _1991_/CLK _1889_/D VGND VGND VPWR VPWR _1890_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_103_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1812_ _1816_/CLK _1812_/D VGND VGND VPWR VPWR _1813_/D sky130_fd_sc_hd__dfxtp_1
X_1743_ _1747_/CLK _1743_/D VGND VGND VPWR VPWR _1744_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1674_ _1687_/CLK _1674_/D VGND VGND VPWR VPWR _1675_/D sky130_fd_sc_hd__dfxtp_1
X_0625_ _0632_/CLK _0625_/D VGND VGND VPWR VPWR _0626_/D sky130_fd_sc_hd__dfxtp_1
X_0556_ _0573_/CLK _0556_/D VGND VGND VPWR VPWR _0557_/D sky130_fd_sc_hd__dfxtp_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0487_ _0998_/CLK _0487_/D VGND VGND VPWR VPWR _0488_/D sky130_fd_sc_hd__dfxtp_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1108_ _1112_/CLK _1108_/D VGND VGND VPWR VPWR _1109_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_53_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1039_ _1039_/CLK _1039_/D VGND VGND VPWR VPWR _1040_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_41_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_110_clk clkbuf_4_1_0_clk/X VGND VGND VPWR VPWR _1794_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_89_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_101_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _1673_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0410_ _0622_/CLK _0410_/D VGND VGND VPWR VPWR _0411_/D sky130_fd_sc_hd__dfxtp_1
X_1390_ _1754_/CLK _1390_/D VGND VGND VPWR VPWR _1391_/D sky130_fd_sc_hd__dfxtp_1
X_0341_ _0539_/CLK _0341_/D VGND VGND VPWR VPWR _0352_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_79_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0272_ _0280_/CLK _0272_/D VGND VGND VPWR VPWR _0273_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1726_ _1726_/CLK _1726_/D VGND VGND VPWR VPWR _1727_/D sky130_fd_sc_hd__dfxtp_1
X_1657_ _1659_/CLK _1657_/D VGND VGND VPWR VPWR _1658_/D sky130_fd_sc_hd__dfxtp_1
X_0608_ _0610_/CLK _0608_/D VGND VGND VPWR VPWR _0609_/D sky130_fd_sc_hd__dfxtp_1
X_1588_ _1592_/CLK _1588_/D VGND VGND VPWR VPWR _1589_/D sky130_fd_sc_hd__dfxtp_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0539_ _0539_/CLK _0539_/D VGND VGND VPWR VPWR _0550_/D sky130_fd_sc_hd__dfxtp_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0890_ _0894_/CLK _0890_/D VGND VGND VPWR VPWR _0892_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_9_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1511_ _1604_/CLK _1511_/D VGND VGND VPWR VPWR _1512_/D sky130_fd_sc_hd__dfxtp_1
X_1442_ _1686_/CLK _1442_/D VGND VGND VPWR VPWR _1443_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1373_ _1373_/CLK _1373_/D VGND VGND VPWR VPWR _1374_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0324_ _1071_/CLK _0324_/D VGND VGND VPWR VPWR _0325_/D sky130_fd_sc_hd__dfxtp_1
X_0255_ _1973_/CLK _0255_/D VGND VGND VPWR VPWR _0256_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0186_ _0214_/CLK _0186_/D VGND VGND VPWR VPWR _0188_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1709_ _1726_/CLK _1709_/D VGND VGND VPWR VPWR _1710_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0040_ _0169_/CLK _0040_/D VGND VGND VPWR VPWR _0041_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1991_ _1991_/CLK _1991_/D VGND VGND VPWR VPWR _1992_/D sky130_fd_sc_hd__dfxtp_1
X_0942_ _0953_/CLK _0942_/D VGND VGND VPWR VPWR _0943_/D sky130_fd_sc_hd__dfxtp_1
X_0873_ _0874_/CLK _0873_/D VGND VGND VPWR VPWR _0874_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_9_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1425_ _1794_/CLK _1425_/D VGND VGND VPWR VPWR _1426_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1356_ _1364_/CLK _1356_/D VGND VGND VPWR VPWR _1357_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_56_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0307_ _1046_/CLK _0307_/D VGND VGND VPWR VPWR _0309_/D sky130_fd_sc_hd__dfxtp_1
X_1287_ _1348_/CLK _1287_/D VGND VGND VPWR VPWR _1288_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_55_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0238_ _1996_/CLK _0238_/D VGND VGND VPWR VPWR _0239_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_90_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _1578_/CLK sky130_fd_sc_hd__clkbuf_16
X_0169_ _0169_/CLK _0169_/D VGND VGND VPWR VPWR _0170_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_51_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _1985_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1210_ _1233_/CLK _1210_/D VGND VGND VPWR VPWR _1211_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_37_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1141_ _1147_/CLK _1141_/D VGND VGND VPWR VPWR _1142_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1072_ _1077_/CLK _1072_/D VGND VGND VPWR VPWR _1073_/D sky130_fd_sc_hd__dfxtp_1
X_0023_ _1858_/CLK _0023_/D VGND VGND VPWR VPWR _0024_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_33_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_72_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _1046_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1974_ _1980_/CLK _1974_/D VGND VGND VPWR VPWR _1975_/D sky130_fd_sc_hd__dfxtp_1
X_0925_ _0932_/CLK _0925_/D VGND VGND VPWR VPWR _0926_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_106_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0856_ _0864_/CLK _0856_/D VGND VGND VPWR VPWR _0857_/D sky130_fd_sc_hd__dfxtp_1
X_0787_ _0813_/CLK _0787_/D VGND VGND VPWR VPWR _0788_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_0_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1408_ _1710_/CLK _1408_/D VGND VGND VPWR VPWR _1409_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_56_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1339_ _1772_/CLK _1339_/D VGND VGND VPWR VPWR _1340_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_63_clk clkbuf_4_15_0_clk/X VGND VGND VPWR VPWR _0977_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _0610_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0710_ _0793_/CLK _0710_/D VGND VGND VPWR VPWR _0711_/D sky130_fd_sc_hd__dfxtp_1
X_1690_ _1695_/CLK _1690_/D VGND VGND VPWR VPWR _1691_/D sky130_fd_sc_hd__dfxtp_1
X_0641_ _0642_/CLK _0641_/D VGND VGND VPWR VPWR _0642_/D sky130_fd_sc_hd__dfxtp_1
X_0572_ _1649_/CLK _0572_/D VGND VGND VPWR VPWR _0583_/D sky130_fd_sc_hd__dfxtp_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1124_ _1127_/CLK _1124_/D VGND VGND VPWR VPWR _1125_/D sky130_fd_sc_hd__dfxtp_1
X_1055_ _1055_/CLK _1055_/D VGND VGND VPWR VPWR _1057_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0006_ _1997_/CLK _0006_/D VGND VGND VPWR VPWR _0007_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_45_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _1178_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1957_ _1973_/CLK _1957_/D VGND VGND VPWR VPWR _1958_/D sky130_fd_sc_hd__dfxtp_1
X_0908_ _0908_/CLK _0908_/D VGND VGND VPWR VPWR _0909_/D sky130_fd_sc_hd__dfxtp_1
X_1888_ _1987_/CLK _1888_/D VGND VGND VPWR VPWR _1899_/D sky130_fd_sc_hd__dfxtp_1
X_0839_ _0845_/CLK _0839_/D VGND VGND VPWR VPWR _0840_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_102_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_36_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _0919_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _0831_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1811_ _1833_/CLK _1811_/D VGND VGND VPWR VPWR _1822_/D sky130_fd_sc_hd__dfxtp_1
X_1742_ _1747_/CLK _1742_/D VGND VGND VPWR VPWR _1743_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1673_ _1673_/CLK _1673_/D VGND VGND VPWR VPWR _1674_/D sky130_fd_sc_hd__dfxtp_1
X_0624_ _0632_/CLK _0624_/D VGND VGND VPWR VPWR _0625_/D sky130_fd_sc_hd__dfxtp_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0555_ _0573_/CLK _0555_/D VGND VGND VPWR VPWR _0556_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_97_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0486_ _0977_/CLK _0486_/D VGND VGND VPWR VPWR _0487_/D sky130_fd_sc_hd__dfxtp_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1107_ _1112_/CLK _1107_/D VGND VGND VPWR VPWR _1108_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_18_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _1127_/CLK sky130_fd_sc_hd__clkbuf_16
X_1038_ _1039_/CLK _1038_/D VGND VGND VPWR VPWR _1039_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0340_ _1181_/CLK _0340_/D VGND VGND VPWR VPWR _0342_/D sky130_fd_sc_hd__dfxtp_1
X_0271_ _0280_/CLK _0271_/D VGND VGND VPWR VPWR _0272_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_63_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1725_ _1736_/CLK _1725_/D VGND VGND VPWR VPWR _1726_/D sky130_fd_sc_hd__dfxtp_1
X_1656_ _1665_/CLK _1656_/D VGND VGND VPWR VPWR _1657_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_7_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _1229_/CLK sky130_fd_sc_hd__clkbuf_16
X_0607_ _0610_/CLK _0607_/D VGND VGND VPWR VPWR _0608_/D sky130_fd_sc_hd__dfxtp_1
X_1587_ _1587_/CLK _1587_/D VGND VGND VPWR VPWR _1588_/D sky130_fd_sc_hd__dfxtp_1
X_0538_ _0573_/CLK _0538_/D VGND VGND VPWR VPWR _0540_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0469_ _0508_/CLK _0469_/D VGND VGND VPWR VPWR _0470_/D sky130_fd_sc_hd__dfxtp_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1510_ _1604_/CLK _1510_/D VGND VGND VPWR VPWR _1511_/D sky130_fd_sc_hd__dfxtp_1
X_1441_ _1686_/CLK _1441_/D VGND VGND VPWR VPWR _1442_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1372_ _1764_/CLK _1372_/D VGND VGND VPWR VPWR _1373_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0323_ _1071_/CLK _0323_/D VGND VGND VPWR VPWR _0324_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0254_ _1973_/CLK _0254_/D VGND VGND VPWR VPWR _0255_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0185_ _1858_/CLK _0185_/D VGND VGND VPWR VPWR _0186_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_51_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1708_ _1736_/CLK _1708_/D VGND VGND VPWR VPWR _1709_/D sky130_fd_sc_hd__dfxtp_1
X_1639_ _1659_/CLK _1639_/D VGND VGND VPWR VPWR _1640_/D sky130_fd_sc_hd__dfxtp_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1990_ _1991_/CLK _1990_/D VGND VGND VPWR VPWR _1991_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_54_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0941_ _1077_/CLK _0941_/D VGND VGND VPWR VPWR _0942_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0872_ _0874_/CLK _0872_/D VGND VGND VPWR VPWR _0873_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_9_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1424_ _1794_/CLK _1424_/D VGND VGND VPWR VPWR _1425_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1355_ _1364_/CLK _1355_/D VGND VGND VPWR VPWR _1356_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0306_ _1033_/CLK _0306_/D VGND VGND VPWR VPWR _0307_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1286_ _1336_/CLK _1286_/D VGND VGND VPWR VPWR _1287_/D sky130_fd_sc_hd__dfxtp_1
X_0237_ _0295_/CLK _0237_/D VGND VGND VPWR VPWR _0238_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_70_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0168_ _0169_/CLK _0168_/D VGND VGND VPWR VPWR _0169_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_24_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0099_ _1635_/CLK _0099_/D VGND VGND VPWR VPWR _0110_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_3_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1140_ _1147_/CLK _1140_/D VGND VGND VPWR VPWR _1141_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1071_ _1071_/CLK _1071_/D VGND VGND VPWR VPWR _1072_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0022_ _1965_/CLK _0022_/D VGND VGND VPWR VPWR _0033_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_21_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1973_ _1973_/CLK _1973_/D VGND VGND VPWR VPWR _1974_/D sky130_fd_sc_hd__dfxtp_1
X_0924_ _1826_/CLK _0924_/D VGND VGND VPWR VPWR _0935_/D sky130_fd_sc_hd__dfxtp_1
X_0855_ _0864_/CLK _0855_/D VGND VGND VPWR VPWR _0856_/D sky130_fd_sc_hd__dfxtp_1
X_0786_ _0791_/CLK _0786_/D VGND VGND VPWR VPWR _0787_/D sky130_fd_sc_hd__dfxtp_1
X_1407_ _1710_/CLK _1407_/D VGND VGND VPWR VPWR _1408_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1338_ _1772_/CLK _1338_/D VGND VGND VPWR VPWR _1339_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_56_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1269_ _1272_/CLK _1269_/D VGND VGND VPWR VPWR _1270_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_43_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0640_ _0642_/CLK _0640_/D VGND VGND VPWR VPWR _0641_/D sky130_fd_sc_hd__dfxtp_1
X_0571_ _0573_/CLK _0571_/D VGND VGND VPWR VPWR _0573_/D sky130_fd_sc_hd__dfxtp_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1123_ _1127_/CLK _1123_/D VGND VGND VPWR VPWR _1124_/D sky130_fd_sc_hd__dfxtp_1
X_1054_ _1055_/CLK _1054_/D VGND VGND VPWR VPWR _1055_/D sky130_fd_sc_hd__dfxtp_1
X_0005_ _1997_/CLK _0005_/D VGND VGND VPWR VPWR _0006_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_33_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1956_ _1956_/CLK _1956_/D VGND VGND VPWR VPWR _1957_/D sky130_fd_sc_hd__dfxtp_1
X_0907_ _0919_/CLK _0907_/D VGND VGND VPWR VPWR _0908_/D sky130_fd_sc_hd__dfxtp_1
X_1887_ _1991_/CLK _1887_/D VGND VGND VPWR VPWR _1889_/D sky130_fd_sc_hd__dfxtp_1
X_0838_ _0845_/CLK _0838_/D VGND VGND VPWR VPWR _0839_/D sky130_fd_sc_hd__dfxtp_1
X_0769_ _0791_/CLK _0769_/D VGND VGND VPWR VPWR _0771_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_88_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1810_ _1816_/CLK _1810_/D VGND VGND VPWR VPWR _1812_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1741_ _1747_/CLK _1741_/D VGND VGND VPWR VPWR _1742_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1672_ _1687_/CLK _1672_/D VGND VGND VPWR VPWR _1673_/D sky130_fd_sc_hd__dfxtp_1
X_0623_ _0632_/CLK _0623_/D VGND VGND VPWR VPWR _0624_/D sky130_fd_sc_hd__dfxtp_1
X_0554_ _0595_/CLK _0554_/D VGND VGND VPWR VPWR _0555_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0485_ _0998_/CLK _0485_/D VGND VGND VPWR VPWR _0486_/D sky130_fd_sc_hd__dfxtp_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1106_ _1112_/CLK _1106_/D VGND VGND VPWR VPWR _1107_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1037_ _1039_/CLK _1037_/D VGND VGND VPWR VPWR _1038_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_34_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1939_ _1975_/CLK _1939_/D VGND VGND VPWR VPWR _1940_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0270_ _1010_/CLK _0270_/D VGND VGND VPWR VPWR _0271_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1724_ _1833_/CLK _1724_/D VGND VGND VPWR VPWR _1725_/D sky130_fd_sc_hd__dfxtp_1
X_1655_ _1659_/CLK _1655_/D VGND VGND VPWR VPWR _1656_/D sky130_fd_sc_hd__dfxtp_1
X_0606_ _0610_/CLK _0606_/D VGND VGND VPWR VPWR _0607_/D sky130_fd_sc_hd__dfxtp_1
X_1586_ _1587_/CLK _1586_/D VGND VGND VPWR VPWR _1587_/D sky130_fd_sc_hd__dfxtp_1
X_0537_ _0573_/CLK _0537_/D VGND VGND VPWR VPWR _0538_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0468_ _0529_/CLK _0468_/D VGND VGND VPWR VPWR _0469_/D sky130_fd_sc_hd__dfxtp_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0399_ _0642_/CLK _0399_/D VGND VGND VPWR VPWR _0400_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1440_ _1814_/CLK _1440_/D VGND VGND VPWR VPWR _1441_/D sky130_fd_sc_hd__dfxtp_1
X_1371_ _1373_/CLK _1371_/D VGND VGND VPWR VPWR _1372_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0322_ _1055_/CLK _0322_/D VGND VGND VPWR VPWR _0323_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0253_ _1594_/CLK _0253_/D VGND VGND VPWR VPWR _0264_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0184_ _0214_/CLK _0184_/D VGND VGND VPWR VPWR _0185_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_75_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1707_ _1710_/CLK _1707_/D VGND VGND VPWR VPWR _1708_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_105_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1638_ _1659_/CLK _1638_/D VGND VGND VPWR VPWR _1639_/D sky130_fd_sc_hd__dfxtp_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1569_ _1594_/CLK _1569_/D VGND VGND VPWR VPWR _1570_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0940_ _0953_/CLK _0940_/D VGND VGND VPWR VPWR _0941_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0871_ _0874_/CLK _0871_/D VGND VGND VPWR VPWR _0872_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_5_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1423_ _1695_/CLK _1423_/D VGND VGND VPWR VPWR _1424_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1354_ _1364_/CLK _1354_/D VGND VGND VPWR VPWR _1355_/D sky130_fd_sc_hd__dfxtp_1
X_1285_ _1348_/CLK _1285_/D VGND VGND VPWR VPWR _1286_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0305_ _1046_/CLK _0305_/D VGND VGND VPWR VPWR _0306_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0236_ _1980_/CLK _0236_/D VGND VGND VPWR VPWR _0237_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_51_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0167_ _0169_/CLK _0167_/D VGND VGND VPWR VPWR _0168_/D sky130_fd_sc_hd__dfxtp_1
X_0098_ _1226_/CLK _0098_/D VGND VGND VPWR VPWR _0100_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1070_ _1070_/CLK _1070_/D VGND VGND VPWR VPWR _1071_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_33_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0021_ _1858_/CLK _0021_/D VGND VGND VPWR VPWR _0023_/D sky130_fd_sc_hd__dfxtp_1
X_1972_ _1975_/CLK _1972_/D VGND VGND VPWR VPWR _1973_/D sky130_fd_sc_hd__dfxtp_1
X_0923_ _0932_/CLK _0923_/D VGND VGND VPWR VPWR _0925_/D sky130_fd_sc_hd__dfxtp_1
X_0854_ _0874_/CLK _0854_/D VGND VGND VPWR VPWR _0855_/D sky130_fd_sc_hd__dfxtp_1
X_0785_ _0813_/CLK _0785_/D VGND VGND VPWR VPWR _0786_/D sky130_fd_sc_hd__dfxtp_1
X_1406_ _1747_/CLK _1406_/D VGND VGND VPWR VPWR _1407_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1337_ _1772_/CLK _1337_/D VGND VGND VPWR VPWR _1338_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_29_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1268_ _1272_/CLK _1268_/D VGND VGND VPWR VPWR _1269_/D sky130_fd_sc_hd__dfxtp_1
X_1199_ _1808_/CLK _1199_/D VGND VGND VPWR VPWR _1200_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0219_ _0316_/CLK _0219_/D VGND VGND VPWR VPWR _0221_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0570_ _0573_/CLK _0570_/D VGND VGND VPWR VPWR _0571_/D sky130_fd_sc_hd__dfxtp_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1122_ _1841_/CLK _1122_/D VGND VGND VPWR VPWR _1133_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_93_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1053_ _1055_/CLK _1053_/D VGND VGND VPWR VPWR _1054_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0004_ _1997_/CLK _0004_/D VGND VGND VPWR VPWR _0005_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_33_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1955_ _1956_/CLK _1955_/D VGND VGND VPWR VPWR _1956_/D sky130_fd_sc_hd__dfxtp_1
X_0906_ _0906_/CLK _0906_/D VGND VGND VPWR VPWR _0907_/D sky130_fd_sc_hd__dfxtp_1
X_1886_ _1985_/CLK _1886_/D VGND VGND VPWR VPWR _1887_/D sky130_fd_sc_hd__dfxtp_1
X_0837_ _0845_/CLK _0837_/D VGND VGND VPWR VPWR _0838_/D sky130_fd_sc_hd__dfxtp_1
X_0768_ _0791_/CLK _0768_/D VGND VGND VPWR VPWR _0769_/D sky130_fd_sc_hd__dfxtp_1
X_0699_ _0906_/CLK _0699_/D VGND VGND VPWR VPWR _0700_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_69_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_113_clk clkbuf_4_1_0_clk/X VGND VGND VPWR VPWR _1736_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_21_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_104_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _1827_/CLK sky130_fd_sc_hd__clkbuf_16
X_1740_ _1747_/CLK _1740_/D VGND VGND VPWR VPWR _1741_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1671_ _1673_/CLK _1671_/D VGND VGND VPWR VPWR _1672_/D sky130_fd_sc_hd__dfxtp_1
X_0622_ _0622_/CLK _0622_/D VGND VGND VPWR VPWR _0623_/D sky130_fd_sc_hd__dfxtp_1
X_0553_ _0573_/CLK _0553_/D VGND VGND VPWR VPWR _0554_/D sky130_fd_sc_hd__dfxtp_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0484_ _1985_/CLK _0484_/D VGND VGND VPWR VPWR _0495_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_100_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1105_ _1112_/CLK _1105_/D VGND VGND VPWR VPWR _1106_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_26_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1036_ _1046_/CLK _1036_/D VGND VGND VPWR VPWR _1037_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1938_ _1956_/CLK _1938_/D VGND VGND VPWR VPWR _1939_/D sky130_fd_sc_hd__dfxtp_1
X_1869_ _1995_/CLK _1869_/D VGND VGND VPWR VPWR _1870_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_1_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1723_ _1726_/CLK _1723_/D VGND VGND VPWR VPWR _1724_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_104_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1654_ _1659_/CLK _1654_/D VGND VGND VPWR VPWR _1655_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1585_ _1592_/CLK _1585_/D VGND VGND VPWR VPWR _1586_/D sky130_fd_sc_hd__dfxtp_1
X_0605_ _1649_/CLK _0605_/D VGND VGND VPWR VPWR _0616_/D sky130_fd_sc_hd__dfxtp_1
X_0536_ _1182_/CLK _0536_/D VGND VGND VPWR VPWR _0537_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_86_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0467_ _0529_/CLK _0467_/D VGND VGND VPWR VPWR _0468_/D sky130_fd_sc_hd__dfxtp_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0398_ _0642_/CLK _0398_/D VGND VGND VPWR VPWR _0399_/D sky130_fd_sc_hd__dfxtp_1
X_1019_ _1039_/CLK _1019_/D VGND VGND VPWR VPWR _1020_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_34_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1370_ _1373_/CLK _1370_/D VGND VGND VPWR VPWR _1371_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_4_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0321_ _1070_/CLK _0321_/D VGND VGND VPWR VPWR _0322_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0252_ _1980_/CLK _0252_/D VGND VGND VPWR VPWR _0254_/D sky130_fd_sc_hd__dfxtp_1
X_0183_ _1178_/CLK _0183_/D VGND VGND VPWR VPWR _0184_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1706_ _1710_/CLK _1706_/D VGND VGND VPWR VPWR _1707_/D sky130_fd_sc_hd__dfxtp_1
X_1637_ _1659_/CLK _1637_/D VGND VGND VPWR VPWR _1638_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1568_ _1592_/CLK _1568_/D VGND VGND VPWR VPWR _1569_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0519_ _0529_/CLK _0519_/D VGND VGND VPWR VPWR _0520_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_86_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1499_ _1604_/CLK _1499_/D VGND VGND VPWR VPWR _1500_/D sky130_fd_sc_hd__dfxtp_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _1611_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_54_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_84_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _1956_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_45_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0870_ _0874_/CLK _0870_/D VGND VGND VPWR VPWR _0871_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_70_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1422_ _1695_/CLK _1422_/D VGND VGND VPWR VPWR _1423_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_5_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1353_ _1373_/CLK _1353_/D VGND VGND VPWR VPWR _1354_/D sky130_fd_sc_hd__dfxtp_1
X_1284_ _1348_/CLK _1284_/D VGND VGND VPWR VPWR _1285_/D sky130_fd_sc_hd__dfxtp_1
X_0304_ _1046_/CLK _0304_/D VGND VGND VPWR VPWR _0305_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0235_ _1996_/CLK _0235_/D VGND VGND VPWR VPWR _0236_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_75_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _0214_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0166_ _1180_/CLK _0166_/D VGND VGND VPWR VPWR _0167_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_24_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0097_ _1226_/CLK _0097_/D VGND VGND VPWR VPWR _0098_/D sky130_fd_sc_hd__dfxtp_1
X_0999_ _1010_/CLK _0999_/D VGND VGND VPWR VPWR _1000_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_3_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_66_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _1010_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_57_clk clkbuf_4_15_0_clk/X VGND VGND VPWR VPWR _0585_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_92_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0020_ _1858_/CLK _0020_/D VGND VGND VPWR VPWR _0021_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1971_ _1973_/CLK _1971_/D VGND VGND VPWR VPWR _1972_/D sky130_fd_sc_hd__dfxtp_1
X_0922_ _0932_/CLK _0922_/D VGND VGND VPWR VPWR _0923_/D sky130_fd_sc_hd__dfxtp_1
X_0853_ _0874_/CLK _0853_/D VGND VGND VPWR VPWR _0854_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0784_ _0831_/CLK _0784_/D VGND VGND VPWR VPWR _0785_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_96_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1405_ _1747_/CLK _1405_/D VGND VGND VPWR VPWR _1406_/D sky130_fd_sc_hd__dfxtp_1
X_1336_ _1336_/CLK _1336_/D VGND VGND VPWR VPWR _1337_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput1 din VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_48_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _1055_/CLK sky130_fd_sc_hd__clkbuf_16
X_1267_ _1272_/CLK _1267_/D VGND VGND VPWR VPWR _1268_/D sky130_fd_sc_hd__dfxtp_1
X_1198_ _1233_/CLK _1198_/D VGND VGND VPWR VPWR _1199_/D sky130_fd_sc_hd__dfxtp_1
X_0218_ _1996_/CLK _0218_/D VGND VGND VPWR VPWR _0219_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0149_ _1170_/CLK _0149_/D VGND VGND VPWR VPWR _0150_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_51_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_39_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _1104_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1121_ _1127_/CLK _1121_/D VGND VGND VPWR VPWR _1123_/D sky130_fd_sc_hd__dfxtp_1
X_1052_ _1055_/CLK _1052_/D VGND VGND VPWR VPWR _1053_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0003_ _1997_/CLK _0003_/D VGND VGND VPWR VPWR _0004_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_46_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1954_ _1987_/CLK _1954_/D VGND VGND VPWR VPWR _1965_/D sky130_fd_sc_hd__dfxtp_1
X_0905_ _0908_/CLK _0905_/D VGND VGND VPWR VPWR _0906_/D sky130_fd_sc_hd__dfxtp_1
X_1885_ _1985_/CLK _1885_/D VGND VGND VPWR VPWR _1886_/D sky130_fd_sc_hd__dfxtp_1
X_0836_ _1827_/CLK _0836_/D VGND VGND VPWR VPWR _0847_/D sky130_fd_sc_hd__dfxtp_1
X_0767_ _0791_/CLK _0767_/D VGND VGND VPWR VPWR _0768_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_88_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0698_ _1103_/CLK _0698_/D VGND VGND VPWR VPWR _0699_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_96_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1319_ _1788_/CLK _1319_/D VGND VGND VPWR VPWR _1320_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1670_ _1673_/CLK _1670_/D VGND VGND VPWR VPWR _1671_/D sky130_fd_sc_hd__dfxtp_1
X_0621_ _0622_/CLK _0621_/D VGND VGND VPWR VPWR _0622_/D sky130_fd_sc_hd__dfxtp_1
X_0552_ _0573_/CLK _0552_/D VGND VGND VPWR VPWR _0553_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0483_ _0998_/CLK _0483_/D VGND VGND VPWR VPWR _0485_/D sky130_fd_sc_hd__dfxtp_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1104_ _1104_/CLK _1104_/D VGND VGND VPWR VPWR _1105_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1035_ _1046_/CLK _1035_/D VGND VGND VPWR VPWR _1036_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1937_ _1956_/CLK _1937_/D VGND VGND VPWR VPWR _1938_/D sky130_fd_sc_hd__dfxtp_1
X_1868_ _1995_/CLK _1868_/D VGND VGND VPWR VPWR _1869_/D sky130_fd_sc_hd__dfxtp_1
X_0819_ _0898_/CLK _0819_/D VGND VGND VPWR VPWR _0820_/D sky130_fd_sc_hd__dfxtp_1
X_1799_ _1808_/CLK _1799_/D VGND VGND VPWR VPWR _1801_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_1_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1722_ _1736_/CLK _1722_/D VGND VGND VPWR VPWR _1723_/D sky130_fd_sc_hd__dfxtp_1
X_1653_ _1659_/CLK _1653_/D VGND VGND VPWR VPWR _1654_/D sky130_fd_sc_hd__dfxtp_1
X_0604_ _0610_/CLK _0604_/D VGND VGND VPWR VPWR _0606_/D sky130_fd_sc_hd__dfxtp_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1584_ _1587_/CLK _1584_/D VGND VGND VPWR VPWR _1585_/D sky130_fd_sc_hd__dfxtp_1
X_0535_ _0573_/CLK _0535_/D VGND VGND VPWR VPWR _0536_/D sky130_fd_sc_hd__dfxtp_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0466_ _1182_/CLK _0466_/D VGND VGND VPWR VPWR _0467_/D sky130_fd_sc_hd__dfxtp_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0397_ _0642_/CLK _0397_/D VGND VGND VPWR VPWR _0398_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1018_ _1039_/CLK _1018_/D VGND VGND VPWR VPWR _1019_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0320_ _1055_/CLK _0320_/D VGND VGND VPWR VPWR _0321_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_0_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0251_ _1973_/CLK _0251_/D VGND VGND VPWR VPWR _0252_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_82_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0182_ _1178_/CLK _0182_/D VGND VGND VPWR VPWR _0183_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_84_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1705_ _1726_/CLK _1705_/D VGND VGND VPWR VPWR _1706_/D sky130_fd_sc_hd__dfxtp_1
X_1636_ _1673_/CLK _1636_/D VGND VGND VPWR VPWR _1637_/D sky130_fd_sc_hd__dfxtp_1
X_1567_ _1594_/CLK _1567_/D VGND VGND VPWR VPWR _1568_/D sky130_fd_sc_hd__dfxtp_1
X_0518_ _0529_/CLK _0518_/D VGND VGND VPWR VPWR _0519_/D sky130_fd_sc_hd__dfxtp_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1498_ _1600_/CLK _1498_/D VGND VGND VPWR VPWR _1499_/D sky130_fd_sc_hd__dfxtp_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0449_ _0585_/CLK _0449_/D VGND VGND VPWR VPWR _0450_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1421_ _1783_/CLK _1421_/D VGND VGND VPWR VPWR _1422_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1352_ _1364_/CLK _1352_/D VGND VGND VPWR VPWR _1353_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1283_ _1348_/CLK _1283_/D VGND VGND VPWR VPWR _1284_/D sky130_fd_sc_hd__dfxtp_1
X_0303_ _1046_/CLK _0303_/D VGND VGND VPWR VPWR _0304_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0234_ _0316_/CLK _0234_/D VGND VGND VPWR VPWR _0235_/D sky130_fd_sc_hd__dfxtp_1
X_0165_ _1635_/CLK _0165_/D VGND VGND VPWR VPWR _0176_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_24_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0096_ _1226_/CLK _0096_/D VGND VGND VPWR VPWR _0097_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_63_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0998_ _0998_/CLK _0998_/D VGND VGND VPWR VPWR _0999_/D sky130_fd_sc_hd__dfxtp_1
X_1619_ _1673_/CLK _1619_/D VGND VGND VPWR VPWR _1620_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1970_ _1980_/CLK _1970_/D VGND VGND VPWR VPWR _1971_/D sky130_fd_sc_hd__dfxtp_1
X_0921_ _0932_/CLK _0921_/D VGND VGND VPWR VPWR _0922_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_81_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0852_ _0874_/CLK _0852_/D VGND VGND VPWR VPWR _0853_/D sky130_fd_sc_hd__dfxtp_1
X_0783_ _0831_/CLK _0783_/D VGND VGND VPWR VPWR _0784_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1404_ _1747_/CLK _1404_/D VGND VGND VPWR VPWR _1405_/D sky130_fd_sc_hd__dfxtp_1
X_1335_ _1336_/CLK _1335_/D VGND VGND VPWR VPWR _1336_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1266_ _1320_/CLK _1266_/D VGND VGND VPWR VPWR _1267_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_49_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1197_ _1808_/CLK _1197_/D VGND VGND VPWR VPWR _1198_/D sky130_fd_sc_hd__dfxtp_1
X_0217_ _0316_/CLK _0217_/D VGND VGND VPWR VPWR _0218_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0148_ _1162_/CLK _0148_/D VGND VGND VPWR VPWR _0149_/D sky130_fd_sc_hd__dfxtp_1
X_0079_ _1228_/CLK _0079_/D VGND VGND VPWR VPWR _0080_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1120_ _1127_/CLK _1120_/D VGND VGND VPWR VPWR _1121_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_93_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1051_ _1055_/CLK _1051_/D VGND VGND VPWR VPWR _1052_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0002_ _1997_/CLK _0002_/D VGND VGND VPWR VPWR _0003_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_21_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1953_ _1956_/CLK _1953_/D VGND VGND VPWR VPWR _1955_/D sky130_fd_sc_hd__dfxtp_1
X_0904_ _0908_/CLK _0904_/D VGND VGND VPWR VPWR _0905_/D sky130_fd_sc_hd__dfxtp_1
X_1884_ _1985_/CLK _1884_/D VGND VGND VPWR VPWR _1885_/D sky130_fd_sc_hd__dfxtp_1
X_0835_ _0845_/CLK _0835_/D VGND VGND VPWR VPWR _0837_/D sky130_fd_sc_hd__dfxtp_1
X_0766_ _0791_/CLK _0766_/D VGND VGND VPWR VPWR _0767_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0697_ _0906_/CLK _0697_/D VGND VGND VPWR VPWR _0698_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_69_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1318_ _1794_/CLK _1318_/D VGND VGND VPWR VPWR _1319_/D sky130_fd_sc_hd__dfxtp_1
X_1249_ _1272_/CLK _1249_/D VGND VGND VPWR VPWR _1250_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_56_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0620_ _0622_/CLK _0620_/D VGND VGND VPWR VPWR _0621_/D sky130_fd_sc_hd__dfxtp_1
X_0551_ _0573_/CLK _0551_/D VGND VGND VPWR VPWR _0552_/D sky130_fd_sc_hd__dfxtp_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0482_ _0977_/CLK _0482_/D VGND VGND VPWR VPWR _0483_/D sky130_fd_sc_hd__dfxtp_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1103_ _1103_/CLK _1103_/D VGND VGND VPWR VPWR _1104_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_38_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1034_ _1814_/CLK _1034_/D VGND VGND VPWR VPWR _1045_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_61_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1936_ _1936_/CLK _1936_/D VGND VGND VPWR VPWR _1937_/D sky130_fd_sc_hd__dfxtp_1
X_1867_ _1995_/CLK _1867_/D VGND VGND VPWR VPWR _1868_/D sky130_fd_sc_hd__dfxtp_1
X_0818_ _0898_/CLK _0818_/D VGND VGND VPWR VPWR _0819_/D sky130_fd_sc_hd__dfxtp_1
X_1798_ _1808_/CLK _1798_/D VGND VGND VPWR VPWR _1799_/D sky130_fd_sc_hd__dfxtp_1
X_0749_ _0761_/CLK _0749_/D VGND VGND VPWR VPWR _0750_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_88_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1721_ _1726_/CLK _1721_/D VGND VGND VPWR VPWR _1722_/D sky130_fd_sc_hd__dfxtp_1
X_1652_ _1659_/CLK _1652_/D VGND VGND VPWR VPWR _1653_/D sky130_fd_sc_hd__dfxtp_1
X_0603_ _0610_/CLK _0603_/D VGND VGND VPWR VPWR _0604_/D sky130_fd_sc_hd__dfxtp_1
X_1583_ _1587_/CLK _1583_/D VGND VGND VPWR VPWR _1584_/D sky130_fd_sc_hd__dfxtp_1
X_0534_ _1182_/CLK _0534_/D VGND VGND VPWR VPWR _0535_/D sky130_fd_sc_hd__dfxtp_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0465_ _0529_/CLK _0465_/D VGND VGND VPWR VPWR _0466_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_86_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0396_ _1907_/CLK _0396_/D VGND VGND VPWR VPWR _0407_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_39_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1017_ _1017_/CLK _1017_/D VGND VGND VPWR VPWR _1018_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1919_ _1936_/CLK _1919_/D VGND VGND VPWR VPWR _1920_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_103_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0250_ _1980_/CLK _0250_/D VGND VGND VPWR VPWR _0251_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_75_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0181_ _1178_/CLK _0181_/D VGND VGND VPWR VPWR _0182_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_84_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1704_ _1710_/CLK _1704_/D VGND VGND VPWR VPWR _1705_/D sky130_fd_sc_hd__dfxtp_1
X_1635_ _1635_/CLK _1635_/D VGND VGND VPWR VPWR _1636_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1566_ _1592_/CLK _1566_/D VGND VGND VPWR VPWR _1567_/D sky130_fd_sc_hd__dfxtp_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0517_ _0539_/CLK _0517_/D VGND VGND VPWR VPWR _0528_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_59_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1497_ _1604_/CLK _1497_/D VGND VGND VPWR VPWR _1498_/D sky130_fd_sc_hd__dfxtp_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0448_ _0585_/CLK _0448_/D VGND VGND VPWR VPWR _0449_/D sky130_fd_sc_hd__dfxtp_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0379_ _1103_/CLK _0379_/D VGND VGND VPWR VPWR _0380_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_66_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1420_ _1783_/CLK _1420_/D VGND VGND VPWR VPWR _1421_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_79_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1351_ _1364_/CLK _1351_/D VGND VGND VPWR VPWR _1352_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0302_ _1046_/CLK _0302_/D VGND VGND VPWR VPWR _0303_/D sky130_fd_sc_hd__dfxtp_1
X_1282_ _1348_/CLK _1282_/D VGND VGND VPWR VPWR _1283_/D sky130_fd_sc_hd__dfxtp_1
X_0233_ _1996_/CLK _0233_/D VGND VGND VPWR VPWR _0234_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_48_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0164_ _0169_/CLK _0164_/D VGND VGND VPWR VPWR _0166_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_91_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0095_ _1226_/CLK _0095_/D VGND VGND VPWR VPWR _0096_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_51_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0997_ _0998_/CLK _0997_/D VGND VGND VPWR VPWR _0998_/D sky130_fd_sc_hd__dfxtp_1
X_1618_ _1965_/CLK _1618_/D VGND VGND VPWR VPWR _1619_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1549_ _1918_/CLK _1549_/D VGND VGND VPWR VPWR _1550_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0920_ _0932_/CLK _0920_/D VGND VGND VPWR VPWR _0921_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_81_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0851_ _0874_/CLK _0851_/D VGND VGND VPWR VPWR _0852_/D sky130_fd_sc_hd__dfxtp_1
X_0782_ _0831_/CLK _0782_/D VGND VGND VPWR VPWR _0783_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1403_ _1747_/CLK _1403_/D VGND VGND VPWR VPWR _1404_/D sky130_fd_sc_hd__dfxtp_1
X_1334_ _1336_/CLK _1334_/D VGND VGND VPWR VPWR _1335_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1265_ _1320_/CLK _1265_/D VGND VGND VPWR VPWR _1266_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1196_ _1228_/CLK _1196_/D VGND VGND VPWR VPWR _1197_/D sky130_fd_sc_hd__dfxtp_1
X_0216_ _0316_/CLK _0216_/D VGND VGND VPWR VPWR _0217_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0147_ _1162_/CLK _0147_/D VGND VGND VPWR VPWR _0148_/D sky130_fd_sc_hd__dfxtp_1
X_0078_ _1228_/CLK _0078_/D VGND VGND VPWR VPWR _0079_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_116_clk clkbuf_4_1_0_clk/X VGND VGND VPWR VPWR _1783_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1050_ _1055_/CLK _1050_/D VGND VGND VPWR VPWR _1051_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0001_ _1997_/CLK _1997_/Q VGND VGND VPWR VPWR _0002_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_73_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_107_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _1826_/CLK sky130_fd_sc_hd__clkbuf_16
X_1952_ _1956_/CLK _1952_/D VGND VGND VPWR VPWR _1953_/D sky130_fd_sc_hd__dfxtp_1
X_0903_ _0908_/CLK _0903_/D VGND VGND VPWR VPWR _0904_/D sky130_fd_sc_hd__dfxtp_1
X_1883_ _1985_/CLK _1883_/D VGND VGND VPWR VPWR _1884_/D sky130_fd_sc_hd__dfxtp_1
X_0834_ _0845_/CLK _0834_/D VGND VGND VPWR VPWR _0835_/D sky130_fd_sc_hd__dfxtp_1
X_0765_ _0791_/CLK _0765_/D VGND VGND VPWR VPWR _0766_/D sky130_fd_sc_hd__dfxtp_1
X_0696_ _0906_/CLK _0696_/D VGND VGND VPWR VPWR _0697_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_103_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1317_ _1320_/CLK _1317_/D VGND VGND VPWR VPWR _1318_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_56_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1248_ _1272_/CLK _1248_/D VGND VGND VPWR VPWR _1249_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1179_ _1180_/CLK _1179_/D VGND VGND VPWR VPWR _1180_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0550_ _1649_/CLK _0550_/D VGND VGND VPWR VPWR _0561_/D sky130_fd_sc_hd__dfxtp_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0481_ _0977_/CLK _0481_/D VGND VGND VPWR VPWR _0482_/D sky130_fd_sc_hd__dfxtp_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1102_ _1104_/CLK _1102_/D VGND VGND VPWR VPWR _1103_/D sky130_fd_sc_hd__dfxtp_1
X_1033_ _1033_/CLK _1033_/D VGND VGND VPWR VPWR _1035_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_81_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1935_ _1956_/CLK _1935_/D VGND VGND VPWR VPWR _1936_/D sky130_fd_sc_hd__dfxtp_1
X_1866_ _1987_/CLK _1866_/D VGND VGND VPWR VPWR _1877_/D sky130_fd_sc_hd__dfxtp_1
X_0817_ _0831_/CLK _0817_/D VGND VGND VPWR VPWR _0818_/D sky130_fd_sc_hd__dfxtp_1
X_1797_ _1808_/CLK _1797_/D VGND VGND VPWR VPWR _1798_/D sky130_fd_sc_hd__dfxtp_1
X_0748_ _1827_/CLK _0748_/D VGND VGND VPWR VPWR _0759_/D sky130_fd_sc_hd__dfxtp_1
X_0679_ _0898_/CLK _0679_/D VGND VGND VPWR VPWR _0680_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_84_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1720_ _1833_/CLK _1720_/D VGND VGND VPWR VPWR _1721_/D sky130_fd_sc_hd__dfxtp_1
X_1651_ _1659_/CLK _1651_/D VGND VGND VPWR VPWR _1652_/D sky130_fd_sc_hd__dfxtp_1
X_0602_ _0610_/CLK _0602_/D VGND VGND VPWR VPWR _0603_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1582_ _1592_/CLK _1582_/D VGND VGND VPWR VPWR _1583_/D sky130_fd_sc_hd__dfxtp_1
X_0533_ _1182_/CLK _0533_/D VGND VGND VPWR VPWR _0534_/D sky130_fd_sc_hd__dfxtp_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0464_ _1182_/CLK _0464_/D VGND VGND VPWR VPWR _0465_/D sky130_fd_sc_hd__dfxtp_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0395_ _0642_/CLK _0395_/D VGND VGND VPWR VPWR _0397_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_93_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1016_ _1017_/CLK _1016_/D VGND VGND VPWR VPWR _1017_/D sky130_fd_sc_hd__dfxtp_1
X_1918_ _1918_/CLK _1918_/D VGND VGND VPWR VPWR _1919_/D sky130_fd_sc_hd__dfxtp_1
X_1849_ _1862_/CLK _1849_/D VGND VGND VPWR VPWR _1850_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_96_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _1965_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_20_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _1138_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_87_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _1907_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0180_ _1178_/CLK _0180_/D VGND VGND VPWR VPWR _0181_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_29_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _1816_/CLK sky130_fd_sc_hd__clkbuf_16
X_1703_ _1736_/CLK _1703_/D VGND VGND VPWR VPWR _1704_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_8_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1634_ _1673_/CLK _1634_/D VGND VGND VPWR VPWR _1635_/D sky130_fd_sc_hd__dfxtp_1
X_1565_ _1594_/CLK _1565_/D VGND VGND VPWR VPWR _1566_/D sky130_fd_sc_hd__dfxtp_1
X_0516_ _0529_/CLK _0516_/D VGND VGND VPWR VPWR _0518_/D sky130_fd_sc_hd__dfxtp_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1496_ _1600_/CLK _1496_/D VGND VGND VPWR VPWR _1497_/D sky130_fd_sc_hd__dfxtp_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0447_ _0973_/CLK _0447_/D VGND VGND VPWR VPWR _0448_/D sky130_fd_sc_hd__dfxtp_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_78_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _1995_/CLK sky130_fd_sc_hd__clkbuf_16
X_0378_ _1103_/CLK _0378_/D VGND VGND VPWR VPWR _0379_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_69_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _1980_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1350_ _1373_/CLK _1350_/D VGND VGND VPWR VPWR _1351_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0301_ _1046_/CLK _0301_/D VGND VGND VPWR VPWR _0302_/D sky130_fd_sc_hd__dfxtp_1
X_1281_ _1348_/CLK _1281_/D VGND VGND VPWR VPWR _1282_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _1348_/CLK sky130_fd_sc_hd__clkbuf_16
X_0232_ _1996_/CLK _0232_/D VGND VGND VPWR VPWR _0233_/D sky130_fd_sc_hd__dfxtp_1
X_0163_ _0169_/CLK _0163_/D VGND VGND VPWR VPWR _0164_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0094_ _1226_/CLK _0094_/D VGND VGND VPWR VPWR _0095_/D sky130_fd_sc_hd__dfxtp_1
X_0996_ _1017_/CLK _0996_/D VGND VGND VPWR VPWR _0997_/D sky130_fd_sc_hd__dfxtp_1
X_1617_ _1833_/CLK _1617_/D VGND VGND VPWR VPWR _1618_/D sky130_fd_sc_hd__dfxtp_1
X_1548_ _1592_/CLK _1548_/D VGND VGND VPWR VPWR _1549_/D sky130_fd_sc_hd__dfxtp_1
X_1479_ _1833_/CLK _1479_/D VGND VGND VPWR VPWR _1480_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0850_ _0864_/CLK _0850_/D VGND VGND VPWR VPWR _0851_/D sky130_fd_sc_hd__dfxtp_1
X_0781_ _1827_/CLK _0781_/D VGND VGND VPWR VPWR _0792_/D sky130_fd_sc_hd__dfxtp_1
X_1402_ _1747_/CLK _1402_/D VGND VGND VPWR VPWR _1403_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_96_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1333_ _1336_/CLK _1333_/D VGND VGND VPWR VPWR _1334_/D sky130_fd_sc_hd__dfxtp_1
X_1264_ _1320_/CLK _1264_/D VGND VGND VPWR VPWR _1265_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0215_ _0316_/CLK _0215_/D VGND VGND VPWR VPWR _0216_/D sky130_fd_sc_hd__dfxtp_1
X_1195_ _1816_/CLK _1195_/D VGND VGND VPWR VPWR _1196_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0146_ _1162_/CLK _0146_/D VGND VGND VPWR VPWR _0147_/D sky130_fd_sc_hd__dfxtp_1
X_0077_ _1635_/CLK _0077_/D VGND VGND VPWR VPWR _0088_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_24_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0979_ _1826_/CLK _0979_/D VGND VGND VPWR VPWR _0990_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0000_ _1965_/CLK _1987_/Q VGND VGND VPWR VPWR _0011_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_34_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1951_ _1975_/CLK _1951_/D VGND VGND VPWR VPWR _1952_/D sky130_fd_sc_hd__dfxtp_1
X_0902_ _1827_/CLK _0902_/D VGND VGND VPWR VPWR _0913_/D sky130_fd_sc_hd__dfxtp_1
X_1882_ _1985_/CLK _1882_/D VGND VGND VPWR VPWR _1883_/D sky130_fd_sc_hd__dfxtp_1
X_0833_ _0845_/CLK _0833_/D VGND VGND VPWR VPWR _0834_/D sky130_fd_sc_hd__dfxtp_1
X_0764_ _0791_/CLK _0764_/D VGND VGND VPWR VPWR _0765_/D sky130_fd_sc_hd__dfxtp_1
X_0695_ _0906_/CLK _0695_/D VGND VGND VPWR VPWR _0696_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_69_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1316_ _1808_/CLK _1316_/D VGND VGND VPWR VPWR _1317_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_84_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1247_ _1272_/CLK _1247_/D VGND VGND VPWR VPWR _1248_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_56_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1178_ _1178_/CLK _1178_/D VGND VGND VPWR VPWR _1179_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0129_ _1138_/CLK _0129_/D VGND VGND VPWR VPWR _0130_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0480_ _0977_/CLK _0480_/D VGND VGND VPWR VPWR _0481_/D sky130_fd_sc_hd__dfxtp_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1101_ _1103_/CLK _1101_/D VGND VGND VPWR VPWR _1102_/D sky130_fd_sc_hd__dfxtp_1
X_1032_ _1046_/CLK _1032_/D VGND VGND VPWR VPWR _1033_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1934_ _1956_/CLK _1934_/D VGND VGND VPWR VPWR _1935_/D sky130_fd_sc_hd__dfxtp_1
X_1865_ _1995_/CLK _1865_/D VGND VGND VPWR VPWR _1867_/D sky130_fd_sc_hd__dfxtp_1
X_0816_ _0898_/CLK _0816_/D VGND VGND VPWR VPWR _0817_/D sky130_fd_sc_hd__dfxtp_1
X_1796_ _1814_/CLK _1796_/D VGND VGND VPWR VPWR _1797_/D sky130_fd_sc_hd__dfxtp_1
X_0747_ _0750_/CLK _0747_/D VGND VGND VPWR VPWR _0749_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0678_ _0898_/CLK _0678_/D VGND VGND VPWR VPWR _0679_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1650_ _1659_/CLK _1650_/D VGND VGND VPWR VPWR _1651_/D sky130_fd_sc_hd__dfxtp_1
X_0601_ _0610_/CLK _0601_/D VGND VGND VPWR VPWR _0602_/D sky130_fd_sc_hd__dfxtp_1
X_1581_ _1587_/CLK _1581_/D VGND VGND VPWR VPWR _1582_/D sky130_fd_sc_hd__dfxtp_1
X_0532_ _1182_/CLK _0532_/D VGND VGND VPWR VPWR _0533_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0463_ _1182_/CLK _0463_/D VGND VGND VPWR VPWR _0464_/D sky130_fd_sc_hd__dfxtp_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0394_ _0642_/CLK _0394_/D VGND VGND VPWR VPWR _0395_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1015_ _1017_/CLK _1015_/D VGND VGND VPWR VPWR _1016_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_34_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1917_ _1936_/CLK _1917_/D VGND VGND VPWR VPWR _1918_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1848_ _1862_/CLK _1848_/D VGND VGND VPWR VPWR _1849_/D sky130_fd_sc_hd__dfxtp_1
X_1779_ _1783_/CLK _1779_/D VGND VGND VPWR VPWR _1780_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1702_ _1710_/CLK _1702_/D VGND VGND VPWR VPWR _1703_/D sky130_fd_sc_hd__dfxtp_1
X_1633_ _1659_/CLK _1633_/D VGND VGND VPWR VPWR _1634_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1564_ _1594_/CLK _1564_/D VGND VGND VPWR VPWR _1565_/D sky130_fd_sc_hd__dfxtp_1
X_0515_ _0529_/CLK _0515_/D VGND VGND VPWR VPWR _0516_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_86_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1495_ _1600_/CLK _1495_/D VGND VGND VPWR VPWR _1496_/D sky130_fd_sc_hd__dfxtp_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0446_ _0973_/CLK _0446_/D VGND VGND VPWR VPWR _0447_/D sky130_fd_sc_hd__dfxtp_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0377_ _1103_/CLK _0377_/D VGND VGND VPWR VPWR _0378_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_82_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0300_ _1046_/CLK _0300_/D VGND VGND VPWR VPWR _0301_/D sky130_fd_sc_hd__dfxtp_1
X_1280_ _1348_/CLK _1280_/D VGND VGND VPWR VPWR _1281_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0231_ _1594_/CLK _0231_/D VGND VGND VPWR VPWR _0242_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0162_ _0169_/CLK _0162_/D VGND VGND VPWR VPWR _0163_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0093_ _1226_/CLK _0093_/D VGND VGND VPWR VPWR _0094_/D sky130_fd_sc_hd__dfxtp_1
X_0995_ _1017_/CLK _0995_/D VGND VGND VPWR VPWR _0996_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_8_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1616_ _1987_/CLK _1616_/D VGND VGND VPWR VPWR _1617_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1547_ _1578_/CLK _1547_/D VGND VGND VPWR VPWR _1548_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1478_ _1726_/CLK _1478_/D VGND VGND VPWR VPWR _1479_/D sky130_fd_sc_hd__dfxtp_1
X_0429_ _0539_/CLK _0429_/D VGND VGND VPWR VPWR _0440_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_55_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0780_ _0831_/CLK _0780_/D VGND VGND VPWR VPWR _0782_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_5_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1401_ _1747_/CLK _1401_/D VGND VGND VPWR VPWR _1402_/D sky130_fd_sc_hd__dfxtp_1
X_1332_ _1336_/CLK _1332_/D VGND VGND VPWR VPWR _1333_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1263_ _1302_/CLK _1263_/D VGND VGND VPWR VPWR _1264_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_49_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0214_ _0214_/CLK _0214_/D VGND VGND VPWR VPWR _0215_/D sky130_fd_sc_hd__dfxtp_1
X_1194_ _1816_/CLK _1194_/D VGND VGND VPWR VPWR _1195_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_91_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0145_ _1162_/CLK _0145_/D VGND VGND VPWR VPWR _0146_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0076_ _1185_/CLK _0076_/D VGND VGND VPWR VPWR _0078_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0978_ _1039_/CLK _0978_/D VGND VGND VPWR VPWR _0980_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1950_ _1975_/CLK _1950_/D VGND VGND VPWR VPWR _1951_/D sky130_fd_sc_hd__dfxtp_1
X_0901_ _0906_/CLK _0901_/D VGND VGND VPWR VPWR _0903_/D sky130_fd_sc_hd__dfxtp_1
X_1881_ _1985_/CLK _1881_/D VGND VGND VPWR VPWR _1882_/D sky130_fd_sc_hd__dfxtp_1
X_0832_ _0845_/CLK _0832_/D VGND VGND VPWR VPWR _0833_/D sky130_fd_sc_hd__dfxtp_1
X_0763_ _0791_/CLK _0763_/D VGND VGND VPWR VPWR _0764_/D sky130_fd_sc_hd__dfxtp_1
X_0694_ _0906_/CLK _0694_/D VGND VGND VPWR VPWR _0695_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1315_ _1808_/CLK _1315_/D VGND VGND VPWR VPWR _1316_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_56_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1246_ _1272_/CLK _1246_/D VGND VGND VPWR VPWR _1247_/D sky130_fd_sc_hd__dfxtp_1
X_1177_ _1841_/CLK _1177_/D VGND VGND VPWR VPWR _1184_/D sky130_fd_sc_hd__dfxtp_1
X_0128_ _1138_/CLK _0128_/D VGND VGND VPWR VPWR _0129_/D sky130_fd_sc_hd__dfxtp_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0059_ _1170_/CLK _0059_/D VGND VGND VPWR VPWR _0060_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_4_9_0_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1100_ _1846_/CLK _1100_/D VGND VGND VPWR VPWR _1111_/D sky130_fd_sc_hd__dfxtp_1
X_1031_ _1033_/CLK _1031_/D VGND VGND VPWR VPWR _1032_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1933_ _1956_/CLK _1933_/D VGND VGND VPWR VPWR _1934_/D sky130_fd_sc_hd__dfxtp_1
X_1864_ _1997_/CLK _1864_/D VGND VGND VPWR VPWR _1865_/D sky130_fd_sc_hd__dfxtp_1
X_0815_ _0898_/CLK _0815_/D VGND VGND VPWR VPWR _0816_/D sky130_fd_sc_hd__dfxtp_1
X_1795_ _1814_/CLK _1795_/D VGND VGND VPWR VPWR _1796_/D sky130_fd_sc_hd__dfxtp_1
X_0746_ _0761_/CLK _0746_/D VGND VGND VPWR VPWR _0747_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_89_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0677_ _0898_/CLK _0677_/D VGND VGND VPWR VPWR _0678_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_84_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1229_ _1229_/CLK _1229_/D VGND VGND VPWR VPWR _1230_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_25_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0600_ _0610_/CLK _0600_/D VGND VGND VPWR VPWR _0601_/D sky130_fd_sc_hd__dfxtp_1
X_1580_ _1587_/CLK _1580_/D VGND VGND VPWR VPWR _1581_/D sky130_fd_sc_hd__dfxtp_1
X_0531_ _1182_/CLK _0531_/D VGND VGND VPWR VPWR _0532_/D sky130_fd_sc_hd__dfxtp_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0462_ _0539_/CLK _0462_/D VGND VGND VPWR VPWR _0473_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_100_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0393_ _0932_/CLK _0393_/D VGND VGND VPWR VPWR _0394_/D sky130_fd_sc_hd__dfxtp_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1014_ _1017_/CLK _1014_/D VGND VGND VPWR VPWR _1015_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_22_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1916_ _1918_/CLK _1916_/D VGND VGND VPWR VPWR _1917_/D sky130_fd_sc_hd__dfxtp_1
X_1847_ _1862_/CLK _1847_/D VGND VGND VPWR VPWR _1848_/D sky130_fd_sc_hd__dfxtp_1
X_1778_ _1833_/CLK _1778_/D VGND VGND VPWR VPWR _1789_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0729_ _0761_/CLK _0729_/D VGND VGND VPWR VPWR _0730_/D sky130_fd_sc_hd__dfxtp_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1701_ _1710_/CLK _1701_/D VGND VGND VPWR VPWR _1702_/D sky130_fd_sc_hd__dfxtp_1
X_1632_ _1673_/CLK _1632_/D VGND VGND VPWR VPWR _1633_/D sky130_fd_sc_hd__dfxtp_1
X_1563_ _1594_/CLK _1563_/D VGND VGND VPWR VPWR _1564_/D sky130_fd_sc_hd__dfxtp_1
X_0514_ _0529_/CLK _0514_/D VGND VGND VPWR VPWR _0515_/D sky130_fd_sc_hd__dfxtp_1
X_1494_ _1600_/CLK _1494_/D VGND VGND VPWR VPWR _1495_/D sky130_fd_sc_hd__dfxtp_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0445_ _0973_/CLK _0445_/D VGND VGND VPWR VPWR _0446_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_86_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0376_ _1103_/CLK _0376_/D VGND VGND VPWR VPWR _0377_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_82_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0230_ _1996_/CLK _0230_/D VGND VGND VPWR VPWR _0232_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0161_ _0169_/CLK _0161_/D VGND VGND VPWR VPWR _0162_/D sky130_fd_sc_hd__dfxtp_1
X_0092_ _1226_/CLK _0092_/D VGND VGND VPWR VPWR _0093_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_17_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0994_ _0998_/CLK _0994_/D VGND VGND VPWR VPWR _0995_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_105_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1615_ _1833_/CLK _1615_/D VGND VGND VPWR VPWR _1616_/D sky130_fd_sc_hd__dfxtp_1
X_1546_ _1918_/CLK _1546_/D VGND VGND VPWR VPWR _1547_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_59_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1477_ _1833_/CLK _1477_/D VGND VGND VPWR VPWR _1478_/D sky130_fd_sc_hd__dfxtp_1
X_0428_ _0973_/CLK _0428_/D VGND VGND VPWR VPWR _0430_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_86_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0359_ _1112_/CLK _0359_/D VGND VGND VPWR VPWR _0360_/D sky130_fd_sc_hd__dfxtp_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_119_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _1764_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_60_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1400_ _1754_/CLK _1400_/D VGND VGND VPWR VPWR _1401_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_96_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1331_ _1336_/CLK _1331_/D VGND VGND VPWR VPWR _1332_/D sky130_fd_sc_hd__dfxtp_1
X_1262_ _1302_/CLK _1262_/D VGND VGND VPWR VPWR _1263_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0213_ _0316_/CLK _0213_/D VGND VGND VPWR VPWR _0214_/D sky130_fd_sc_hd__dfxtp_1
X_1193_ _1808_/CLK _1193_/D VGND VGND VPWR VPWR _1194_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0144_ _1162_/CLK _0144_/D VGND VGND VPWR VPWR _0145_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0075_ _1185_/CLK _0075_/D VGND VGND VPWR VPWR _0076_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_32_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0977_ _0977_/CLK _0977_/D VGND VGND VPWR VPWR _0978_/D sky130_fd_sc_hd__dfxtp_1
X_1529_ _1578_/CLK _1529_/D VGND VGND VPWR VPWR _1530_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_19_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0900_ _0908_/CLK _0900_/D VGND VGND VPWR VPWR _0901_/D sky130_fd_sc_hd__dfxtp_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1880_ _1995_/CLK _1880_/D VGND VGND VPWR VPWR _1881_/D sky130_fd_sc_hd__dfxtp_1
X_0831_ _0831_/CLK _0831_/D VGND VGND VPWR VPWR _0832_/D sky130_fd_sc_hd__dfxtp_1
X_0762_ _0791_/CLK _0762_/D VGND VGND VPWR VPWR _0763_/D sky130_fd_sc_hd__dfxtp_1
X_0693_ _1665_/CLK _0693_/D VGND VGND VPWR VPWR _0704_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1314_ _1320_/CLK _1314_/D VGND VGND VPWR VPWR _1315_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_69_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1245_ _1272_/CLK _1245_/D VGND VGND VPWR VPWR _1246_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_49_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1176_ _1180_/CLK _1176_/D VGND VGND VPWR VPWR _1178_/D sky130_fd_sc_hd__dfxtp_1
X_0127_ _1138_/CLK _0127_/D VGND VGND VPWR VPWR _0128_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0058_ _1185_/CLK _0058_/D VGND VGND VPWR VPWR _0059_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_50_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _0953_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1030_ _1033_/CLK _1030_/D VGND VGND VPWR VPWR _1031_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_34_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _1112_/CLK sky130_fd_sc_hd__clkbuf_16
X_1932_ _1965_/CLK _1932_/D VGND VGND VPWR VPWR _1943_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1863_ _1995_/CLK _1863_/D VGND VGND VPWR VPWR _1864_/D sky130_fd_sc_hd__dfxtp_1
X_0814_ _1827_/CLK _0814_/D VGND VGND VPWR VPWR _0825_/D sky130_fd_sc_hd__dfxtp_1
X_1794_ _1794_/CLK _1794_/D VGND VGND VPWR VPWR _1795_/D sky130_fd_sc_hd__dfxtp_1
X_0745_ _0750_/CLK _0745_/D VGND VGND VPWR VPWR _0746_/D sky130_fd_sc_hd__dfxtp_1
X_0676_ _0898_/CLK _0676_/D VGND VGND VPWR VPWR _0677_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_69_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1228_ _1228_/CLK _1228_/D VGND VGND VPWR VPWR _1229_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1159_ _1162_/CLK _1159_/D VGND VGND VPWR VPWR _1160_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_32_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _0898_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_99_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _1726_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_23_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _0761_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0530_ _1182_/CLK _0530_/D VGND VGND VPWR VPWR _0531_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0461_ _1182_/CLK _0461_/D VGND VGND VPWR VPWR _0463_/D sky130_fd_sc_hd__dfxtp_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0392_ _1104_/CLK _0392_/D VGND VGND VPWR VPWR _0393_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1013_ _1017_/CLK _1013_/D VGND VGND VPWR VPWR _1014_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_22_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1915_ _1918_/CLK _1915_/D VGND VGND VPWR VPWR _1916_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_14_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _0169_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1846_ _1846_/CLK _1846_/D VGND VGND VPWR VPWR _1847_/D sky130_fd_sc_hd__dfxtp_1
X_1777_ _1783_/CLK _1777_/D VGND VGND VPWR VPWR _1779_/D sky130_fd_sc_hd__dfxtp_1
X_0728_ _0793_/CLK _0728_/D VGND VGND VPWR VPWR _0729_/D sky130_fd_sc_hd__dfxtp_1
X_0659_ _0916_/CLK _0659_/D VGND VGND VPWR VPWR _0661_/D sky130_fd_sc_hd__dfxtp_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_8_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_4_8_0_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1700_ _1710_/CLK _1700_/D VGND VGND VPWR VPWR _1701_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_12_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1631_ _1673_/CLK _1631_/D VGND VGND VPWR VPWR _1632_/D sky130_fd_sc_hd__dfxtp_1
X_1562_ _1594_/CLK _1562_/D VGND VGND VPWR VPWR _1563_/D sky130_fd_sc_hd__dfxtp_1
X_0513_ _0529_/CLK _0513_/D VGND VGND VPWR VPWR _0514_/D sky130_fd_sc_hd__dfxtp_1
X_1493_ _1600_/CLK _1493_/D VGND VGND VPWR VPWR _1494_/D sky130_fd_sc_hd__dfxtp_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0444_ _0973_/CLK _0444_/D VGND VGND VPWR VPWR _0445_/D sky130_fd_sc_hd__dfxtp_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_3_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _1302_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0375_ _1103_/CLK _0375_/D VGND VGND VPWR VPWR _0376_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_94_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1829_ _1846_/CLK _1829_/D VGND VGND VPWR VPWR _1830_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_2_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0160_ _1170_/CLK _0160_/D VGND VGND VPWR VPWR _0161_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_76_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0091_ _1229_/CLK _0091_/D VGND VGND VPWR VPWR _0092_/D sky130_fd_sc_hd__dfxtp_1
X_0993_ _1010_/CLK _0993_/D VGND VGND VPWR VPWR _0994_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1614_ _1833_/CLK _1614_/D VGND VGND VPWR VPWR _1615_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_5_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1545_ _1936_/CLK _1545_/D VGND VGND VPWR VPWR _1546_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1476_ _1726_/CLK _1476_/D VGND VGND VPWR VPWR _1477_/D sky130_fd_sc_hd__dfxtp_1
X_0427_ _0966_/CLK _0427_/D VGND VGND VPWR VPWR _0428_/D sky130_fd_sc_hd__dfxtp_1
X_0358_ _1112_/CLK _0358_/D VGND VGND VPWR VPWR _0359_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_54_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0289_ _0295_/CLK _0289_/D VGND VGND VPWR VPWR _0290_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_70_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1330_ _1336_/CLK _1330_/D VGND VGND VPWR VPWR _1331_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_96_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1261_ _1320_/CLK _1261_/D VGND VGND VPWR VPWR _1262_/D sky130_fd_sc_hd__dfxtp_1
X_1192_ _1816_/CLK _1192_/D VGND VGND VPWR VPWR _1193_/D sky130_fd_sc_hd__dfxtp_1
X_0212_ _0214_/CLK _0212_/D VGND VGND VPWR VPWR _0213_/D sky130_fd_sc_hd__dfxtp_1
X_0143_ _1635_/CLK _0143_/D VGND VGND VPWR VPWR _0154_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0074_ _1816_/CLK _0074_/D VGND VGND VPWR VPWR _0075_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0976_ _0977_/CLK _0976_/D VGND VGND VPWR VPWR _0977_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1528_ _1587_/CLK _1528_/D VGND VGND VPWR VPWR _1529_/D sky130_fd_sc_hd__dfxtp_1
X_1459_ _1695_/CLK _1459_/D VGND VGND VPWR VPWR _1460_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0830_ _0845_/CLK _0830_/D VGND VGND VPWR VPWR _0831_/D sky130_fd_sc_hd__dfxtp_1
X_0761_ _0761_/CLK _0761_/D VGND VGND VPWR VPWR _0762_/D sky130_fd_sc_hd__dfxtp_1
X_0692_ _0906_/CLK _0692_/D VGND VGND VPWR VPWR _0694_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1313_ _1320_/CLK _1313_/D VGND VGND VPWR VPWR _1314_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_84_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1244_ _1244_/CLK _1244_/D VGND VGND VPWR VPWR _1245_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_37_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1175_ _1180_/CLK _1175_/D VGND VGND VPWR VPWR _1176_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0126_ _1138_/CLK _0126_/D VGND VGND VPWR VPWR _0127_/D sky130_fd_sc_hd__dfxtp_1
X_0057_ _1185_/CLK _0057_/D VGND VGND VPWR VPWR _0058_/D sky130_fd_sc_hd__dfxtp_1
X_0959_ _0966_/CLK _0959_/D VGND VGND VPWR VPWR _0960_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_106_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1931_ _1956_/CLK _1931_/D VGND VGND VPWR VPWR _1933_/D sky130_fd_sc_hd__dfxtp_1
X_1862_ _1862_/CLK _1862_/D VGND VGND VPWR VPWR _1863_/D sky130_fd_sc_hd__dfxtp_1
X_0813_ _0813_/CLK _0813_/D VGND VGND VPWR VPWR _0815_/D sky130_fd_sc_hd__dfxtp_1
X_1793_ _1794_/CLK _1793_/D VGND VGND VPWR VPWR _1794_/D sky130_fd_sc_hd__dfxtp_1
X_0744_ _0761_/CLK _0744_/D VGND VGND VPWR VPWR _0745_/D sky130_fd_sc_hd__dfxtp_1
X_0675_ _0874_/CLK _0675_/D VGND VGND VPWR VPWR _0676_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_88_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1227_ _1229_/CLK _1227_/D VGND VGND VPWR VPWR _1228_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_37_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1158_ _1162_/CLK _1158_/D VGND VGND VPWR VPWR _1159_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0109_ _0743_/CLK _0109_/D VGND VGND VPWR VPWR _0111_/D sky130_fd_sc_hd__dfxtp_1
X_1089_ _1841_/CLK _1089_/D VGND VGND VPWR VPWR _1100_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0460_ _0585_/CLK _0460_/D VGND VGND VPWR VPWR _0461_/D sky130_fd_sc_hd__dfxtp_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0391_ _1103_/CLK _0391_/D VGND VGND VPWR VPWR _0392_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1012_ _1686_/CLK _1012_/D VGND VGND VPWR VPWR _1023_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1914_ _1918_/CLK _1914_/D VGND VGND VPWR VPWR _1915_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1845_ _1862_/CLK _1845_/D VGND VGND VPWR VPWR _1846_/D sky130_fd_sc_hd__dfxtp_1
X_1776_ _1783_/CLK _1776_/D VGND VGND VPWR VPWR _1777_/D sky130_fd_sc_hd__dfxtp_1
X_0727_ _0761_/CLK _0727_/D VGND VGND VPWR VPWR _0728_/D sky130_fd_sc_hd__dfxtp_1
X_0658_ _0916_/CLK _0658_/D VGND VGND VPWR VPWR _0659_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_97_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0589_ _0973_/CLK _0589_/D VGND VGND VPWR VPWR _0590_/D sky130_fd_sc_hd__dfxtp_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1630_ _1659_/CLK _1630_/D VGND VGND VPWR VPWR _1631_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1561_ _1594_/CLK _1561_/D VGND VGND VPWR VPWR _1562_/D sky130_fd_sc_hd__dfxtp_1
X_0512_ _0529_/CLK _0512_/D VGND VGND VPWR VPWR _0513_/D sky130_fd_sc_hd__dfxtp_1
X_1492_ _1600_/CLK _1492_/D VGND VGND VPWR VPWR _1493_/D sky130_fd_sc_hd__dfxtp_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0443_ _0973_/CLK _0443_/D VGND VGND VPWR VPWR _0444_/D sky130_fd_sc_hd__dfxtp_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0374_ _1907_/CLK _0374_/D VGND VGND VPWR VPWR _0385_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_81_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1828_ _1846_/CLK _1828_/D VGND VGND VPWR VPWR _1829_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_89_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1759_ _1772_/CLK _1759_/D VGND VGND VPWR VPWR _1760_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0090_ _1229_/CLK _0090_/D VGND VGND VPWR VPWR _0091_/D sky130_fd_sc_hd__dfxtp_1
X_0992_ _1017_/CLK _0992_/D VGND VGND VPWR VPWR _0993_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1613_ _1833_/CLK _1613_/D VGND VGND VPWR VPWR _1614_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_5_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1544_ _1936_/CLK _1544_/D VGND VGND VPWR VPWR _1545_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1475_ _1726_/CLK _1475_/D VGND VGND VPWR VPWR _1476_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_7_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_4_7_0_clk/X sky130_fd_sc_hd__clkbuf_1
X_0426_ _0953_/CLK _0426_/D VGND VGND VPWR VPWR _0427_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_39_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0357_ _1180_/CLK _0357_/D VGND VGND VPWR VPWR _0358_/D sky130_fd_sc_hd__dfxtp_1
X_0288_ _0295_/CLK _0288_/D VGND VGND VPWR VPWR _0289_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1260_ _1302_/CLK _1260_/D VGND VGND VPWR VPWR _1261_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1191_ _1816_/CLK _1191_/D VGND VGND VPWR VPWR _1192_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0211_ _0316_/CLK _0211_/D VGND VGND VPWR VPWR _0212_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_76_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0142_ _1162_/CLK _0142_/D VGND VGND VPWR VPWR _0144_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0073_ _1228_/CLK _0073_/D VGND VGND VPWR VPWR _0074_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0975_ _0977_/CLK _0975_/D VGND VGND VPWR VPWR _0976_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1527_ _1578_/CLK _1527_/D VGND VGND VPWR VPWR _1528_/D sky130_fd_sc_hd__dfxtp_1
X_1458_ _1710_/CLK _1458_/D VGND VGND VPWR VPWR _1459_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0409_ _0622_/CLK _0409_/D VGND VGND VPWR VPWR _0410_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_74_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1389_ _1764_/CLK _1389_/D VGND VGND VPWR VPWR _1390_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0760_ _0791_/CLK _0760_/D VGND VGND VPWR VPWR _0761_/D sky130_fd_sc_hd__dfxtp_1
X_0691_ _0906_/CLK _0691_/D VGND VGND VPWR VPWR _0692_/D sky130_fd_sc_hd__dfxtp_1
X_1312_ _1808_/CLK _1312_/D VGND VGND VPWR VPWR _1313_/D sky130_fd_sc_hd__dfxtp_1
X_1243_ _1244_/CLK _1243_/D VGND VGND VPWR VPWR _1244_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1174_ _1180_/CLK _1174_/D VGND VGND VPWR VPWR _1175_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0125_ _1138_/CLK _0125_/D VGND VGND VPWR VPWR _0126_/D sky130_fd_sc_hd__dfxtp_1
X_0056_ _1185_/CLK _0056_/D VGND VGND VPWR VPWR _0057_/D sky130_fd_sc_hd__dfxtp_1
X_0958_ _0966_/CLK _0958_/D VGND VGND VPWR VPWR _0959_/D sky130_fd_sc_hd__dfxtp_1
X_0889_ _0894_/CLK _0889_/D VGND VGND VPWR VPWR _0890_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1930_ _1956_/CLK _1930_/D VGND VGND VPWR VPWR _1931_/D sky130_fd_sc_hd__dfxtp_1
X_1861_ _1997_/CLK _1861_/D VGND VGND VPWR VPWR _1862_/D sky130_fd_sc_hd__dfxtp_1
X_0812_ _0813_/CLK _0812_/D VGND VGND VPWR VPWR _0813_/D sky130_fd_sc_hd__dfxtp_1
X_1792_ _1794_/CLK _1792_/D VGND VGND VPWR VPWR _1793_/D sky130_fd_sc_hd__dfxtp_1
X_0743_ _0743_/CLK _0743_/D VGND VGND VPWR VPWR _0744_/D sky130_fd_sc_hd__dfxtp_1
X_0674_ _0898_/CLK _0674_/D VGND VGND VPWR VPWR _0675_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_69_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1226_ _1226_/CLK _1226_/D VGND VGND VPWR VPWR _1227_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_25_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1157_ _1162_/CLK _1157_/D VGND VGND VPWR VPWR _1158_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_65_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0108_ _0743_/CLK _0108_/D VGND VGND VPWR VPWR _0109_/D sky130_fd_sc_hd__dfxtp_1
X_1088_ _1088_/CLK _1088_/D VGND VGND VPWR VPWR _1090_/D sky130_fd_sc_hd__dfxtp_1
X_0039_ _0169_/CLK _0039_/D VGND VGND VPWR VPWR _0040_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_100_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _1687_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0390_ _1104_/CLK _0390_/D VGND VGND VPWR VPWR _0391_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1011_ _1017_/CLK _1011_/D VGND VGND VPWR VPWR _1013_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_47_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1913_ _1918_/CLK _1913_/D VGND VGND VPWR VPWR _1914_/D sky130_fd_sc_hd__dfxtp_1
X_1844_ _1987_/CLK _1844_/D VGND VGND VPWR VPWR _1855_/D sky130_fd_sc_hd__dfxtp_1
X_1775_ _1788_/CLK _1775_/D VGND VGND VPWR VPWR _1776_/D sky130_fd_sc_hd__dfxtp_1
X_0726_ _1665_/CLK _0726_/D VGND VGND VPWR VPWR _0737_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_89_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0657_ _0916_/CLK _0657_/D VGND VGND VPWR VPWR _0658_/D sky130_fd_sc_hd__dfxtp_1
X_0588_ _0595_/CLK _0588_/D VGND VGND VPWR VPWR _0589_/D sky130_fd_sc_hd__dfxtp_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1209_ _1320_/CLK _1209_/D VGND VGND VPWR VPWR _1210_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1560_ _1594_/CLK _1560_/D VGND VGND VPWR VPWR _1561_/D sky130_fd_sc_hd__dfxtp_1
X_0511_ _0529_/CLK _0511_/D VGND VGND VPWR VPWR _0512_/D sky130_fd_sc_hd__dfxtp_1
X_1491_ _1965_/CLK _1491_/D VGND VGND VPWR VPWR _1492_/D sky130_fd_sc_hd__dfxtp_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0442_ _0973_/CLK _0442_/D VGND VGND VPWR VPWR _0443_/D sky130_fd_sc_hd__dfxtp_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0373_ _1103_/CLK _0373_/D VGND VGND VPWR VPWR _0375_/D sky130_fd_sc_hd__dfxtp_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1827_ _1827_/CLK _1827_/D VGND VGND VPWR VPWR _1828_/D sky130_fd_sc_hd__dfxtp_1
X_1758_ _1772_/CLK _1758_/D VGND VGND VPWR VPWR _1759_/D sky130_fd_sc_hd__dfxtp_1
X_0709_ _1127_/CLK _0709_/D VGND VGND VPWR VPWR _0710_/D sky130_fd_sc_hd__dfxtp_1
X_1689_ _1695_/CLK _1689_/D VGND VGND VPWR VPWR _1690_/D sky130_fd_sc_hd__dfxtp_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0991_ _1017_/CLK _0991_/D VGND VGND VPWR VPWR _0992_/D sky130_fd_sc_hd__dfxtp_1
X_1612_ _1833_/CLK _1612_/D VGND VGND VPWR VPWR _1613_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1543_ _1918_/CLK _1543_/D VGND VGND VPWR VPWR _1544_/D sky130_fd_sc_hd__dfxtp_1
X_1474_ _1726_/CLK _1474_/D VGND VGND VPWR VPWR _1475_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_5_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0425_ _0953_/CLK _0425_/D VGND VGND VPWR VPWR _0426_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_86_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0356_ _1088_/CLK _0356_/D VGND VGND VPWR VPWR _0357_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0287_ _0295_/CLK _0287_/D VGND VGND VPWR VPWR _0288_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_82_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_80_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _0539_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1190_ _1816_/CLK _1190_/D VGND VGND VPWR VPWR _1191_/D sky130_fd_sc_hd__dfxtp_1
X_0210_ _0214_/CLK _0210_/D VGND VGND VPWR VPWR _0211_/D sky130_fd_sc_hd__dfxtp_1
X_0141_ _1170_/CLK _0141_/D VGND VGND VPWR VPWR _0142_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0072_ _1816_/CLK _0072_/D VGND VGND VPWR VPWR _0073_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_71_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _1033_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0974_ _0977_/CLK _0974_/D VGND VGND VPWR VPWR _0975_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1526_ _1587_/CLK _1526_/D VGND VGND VPWR VPWR _1527_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1457_ _1687_/CLK _1457_/D VGND VGND VPWR VPWR _1458_/D sky130_fd_sc_hd__dfxtp_1
X_0408_ _0622_/CLK _0408_/D VGND VGND VPWR VPWR _0409_/D sky130_fd_sc_hd__dfxtp_1
X_1388_ _1764_/CLK _1388_/D VGND VGND VPWR VPWR _1389_/D sky130_fd_sc_hd__dfxtp_1
X_0339_ _1181_/CLK _0339_/D VGND VGND VPWR VPWR _0340_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_70_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_62_clk clkbuf_4_15_0_clk/X VGND VGND VPWR VPWR _0998_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_53_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _0632_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_6_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_4_6_0_clk/X sky130_fd_sc_hd__clkbuf_1
X_0690_ _0906_/CLK _0690_/D VGND VGND VPWR VPWR _0691_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1311_ _1320_/CLK _1311_/D VGND VGND VPWR VPWR _1312_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_69_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1242_ _1244_/CLK _1242_/D VGND VGND VPWR VPWR _1243_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1173_ _1180_/CLK _1173_/D VGND VGND VPWR VPWR _1174_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0124_ _1138_/CLK _0124_/D VGND VGND VPWR VPWR _0125_/D sky130_fd_sc_hd__dfxtp_1
X_0055_ _1635_/CLK _0055_/D VGND VGND VPWR VPWR _0066_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_44_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _1180_/CLK sky130_fd_sc_hd__clkbuf_16
X_0957_ _1826_/CLK _0957_/D VGND VGND VPWR VPWR _0968_/D sky130_fd_sc_hd__dfxtp_1
X_0888_ _0894_/CLK _0888_/D VGND VGND VPWR VPWR _0889_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1509_ _1604_/CLK _1509_/D VGND VGND VPWR VPWR _1510_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_35_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _0916_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_102_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _0813_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1860_ _1997_/CLK _1860_/D VGND VGND VPWR VPWR _1861_/D sky130_fd_sc_hd__dfxtp_1
X_0811_ _0813_/CLK _0811_/D VGND VGND VPWR VPWR _0812_/D sky130_fd_sc_hd__dfxtp_1
X_1791_ _1794_/CLK _1791_/D VGND VGND VPWR VPWR _1792_/D sky130_fd_sc_hd__dfxtp_1
X_0742_ _0743_/CLK _0742_/D VGND VGND VPWR VPWR _0743_/D sky130_fd_sc_hd__dfxtp_1
X_0673_ _0874_/CLK _0673_/D VGND VGND VPWR VPWR _0674_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1225_ _1226_/CLK _1225_/D VGND VGND VPWR VPWR _1226_/D sky130_fd_sc_hd__dfxtp_1
X_1156_ _1163_/CLK _1156_/D VGND VGND VPWR VPWR _1157_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0107_ _0743_/CLK _0107_/D VGND VGND VPWR VPWR _0108_/D sky130_fd_sc_hd__dfxtp_1
X_1087_ _1088_/CLK _1087_/D VGND VGND VPWR VPWR _1088_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_17_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _1163_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0038_ _0169_/CLK _0038_/D VGND VGND VPWR VPWR _0039_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1989_ _1995_/CLK _1989_/D VGND VGND VPWR VPWR _1990_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1010_ _1010_/CLK _1010_/D VGND VGND VPWR VPWR _1011_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_34_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1912_ _1918_/CLK _1912_/D VGND VGND VPWR VPWR _1913_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1843_ _1846_/CLK _1843_/D VGND VGND VPWR VPWR _1845_/D sky130_fd_sc_hd__dfxtp_1
X_1774_ _1788_/CLK _1774_/D VGND VGND VPWR VPWR _1775_/D sky130_fd_sc_hd__dfxtp_1
X_0725_ _0793_/CLK _0725_/D VGND VGND VPWR VPWR _0727_/D sky130_fd_sc_hd__dfxtp_1
X_0656_ _0916_/CLK _0656_/D VGND VGND VPWR VPWR _0657_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_6_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _1226_/CLK sky130_fd_sc_hd__clkbuf_16
X_0587_ _0595_/CLK _0587_/D VGND VGND VPWR VPWR _0588_/D sky130_fd_sc_hd__dfxtp_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1208_ _1233_/CLK _1208_/D VGND VGND VPWR VPWR _1209_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_53_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1139_ _1147_/CLK _1139_/D VGND VGND VPWR VPWR _1140_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0510_ _0529_/CLK _0510_/D VGND VGND VPWR VPWR _0511_/D sky130_fd_sc_hd__dfxtp_1
X_1490_ _1600_/CLK _1490_/D VGND VGND VPWR VPWR _1491_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0441_ _0973_/CLK _0441_/D VGND VGND VPWR VPWR _0442_/D sky130_fd_sc_hd__dfxtp_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0372_ _1103_/CLK _0372_/D VGND VGND VPWR VPWR _0373_/D sky130_fd_sc_hd__dfxtp_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1826_ _1826_/CLK _1826_/D VGND VGND VPWR VPWR _1827_/D sky130_fd_sc_hd__dfxtp_1
X_1757_ _1772_/CLK _1757_/D VGND VGND VPWR VPWR _1758_/D sky130_fd_sc_hd__dfxtp_1
X_0708_ _1127_/CLK _0708_/D VGND VGND VPWR VPWR _0709_/D sky130_fd_sc_hd__dfxtp_1
X_1688_ _1695_/CLK _1688_/D VGND VGND VPWR VPWR _1689_/D sky130_fd_sc_hd__dfxtp_1
X_0639_ _0919_/CLK _0639_/D VGND VGND VPWR VPWR _0640_/D sky130_fd_sc_hd__dfxtp_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0990_ _1686_/CLK _0990_/D VGND VGND VPWR VPWR _1001_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_8_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1611_ _1611_/CLK _1611_/D VGND VGND VPWR VPWR _1612_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1542_ _1918_/CLK _1542_/D VGND VGND VPWR VPWR _1543_/D sky130_fd_sc_hd__dfxtp_1
X_1473_ _1726_/CLK _1473_/D VGND VGND VPWR VPWR _1474_/D sky130_fd_sc_hd__dfxtp_1
X_0424_ _0953_/CLK _0424_/D VGND VGND VPWR VPWR _0425_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0355_ _1088_/CLK _0355_/D VGND VGND VPWR VPWR _0356_/D sky130_fd_sc_hd__dfxtp_1
X_0286_ _0539_/CLK _0286_/D VGND VGND VPWR VPWR _0297_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1809_ _1814_/CLK _1809_/D VGND VGND VPWR VPWR _1810_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0140_ _1170_/CLK _0140_/D VGND VGND VPWR VPWR _0141_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0071_ _1816_/CLK _0071_/D VGND VGND VPWR VPWR _0072_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_51_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0973_ _0973_/CLK _0973_/D VGND VGND VPWR VPWR _0974_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1525_ _1587_/CLK _1525_/D VGND VGND VPWR VPWR _1526_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1456_ _1710_/CLK _1456_/D VGND VGND VPWR VPWR _1457_/D sky130_fd_sc_hd__dfxtp_1
X_1387_ _1764_/CLK _1387_/D VGND VGND VPWR VPWR _1388_/D sky130_fd_sc_hd__dfxtp_1
X_0407_ _1907_/CLK _0407_/D VGND VGND VPWR VPWR _0418_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0338_ _1070_/CLK _0338_/D VGND VGND VPWR VPWR _0339_/D sky130_fd_sc_hd__dfxtp_1
X_0269_ _0280_/CLK _0269_/D VGND VGND VPWR VPWR _0270_/D sky130_fd_sc_hd__dfxtp_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1310_ _1320_/CLK _1310_/D VGND VGND VPWR VPWR _1311_/D sky130_fd_sc_hd__dfxtp_1
X_1241_ _1244_/CLK _1241_/D VGND VGND VPWR VPWR _1242_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_2_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1172_ _1180_/CLK _1172_/D VGND VGND VPWR VPWR _1173_/D sky130_fd_sc_hd__dfxtp_1
X_0123_ _1138_/CLK _0123_/D VGND VGND VPWR VPWR _0124_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0054_ _0169_/CLK _0054_/D VGND VGND VPWR VPWR _0056_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0956_ _0966_/CLK _0956_/D VGND VGND VPWR VPWR _0958_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0887_ _0916_/CLK _0887_/D VGND VGND VPWR VPWR _0888_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_102_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1508_ _1611_/CLK _1508_/D VGND VGND VPWR VPWR _1509_/D sky130_fd_sc_hd__dfxtp_1
X_1439_ _1686_/CLK _1439_/D VGND VGND VPWR VPWR _1440_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0810_ _0831_/CLK _0810_/D VGND VGND VPWR VPWR _0811_/D sky130_fd_sc_hd__dfxtp_1
X_1790_ _1794_/CLK _1790_/D VGND VGND VPWR VPWR _1791_/D sky130_fd_sc_hd__dfxtp_1
X_0741_ _0743_/CLK _0741_/D VGND VGND VPWR VPWR _0742_/D sky130_fd_sc_hd__dfxtp_1
X_0672_ _0874_/CLK _0672_/D VGND VGND VPWR VPWR _0673_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1224_ _1226_/CLK _1224_/D VGND VGND VPWR VPWR _1225_/D sky130_fd_sc_hd__dfxtp_1
X_1155_ _1185_/CLK _1155_/D VGND VGND VPWR VPWR _1166_/D sky130_fd_sc_hd__dfxtp_1
X_0106_ _0743_/CLK _0106_/D VGND VGND VPWR VPWR _0107_/D sky130_fd_sc_hd__dfxtp_1
X_1086_ _1088_/CLK _1086_/D VGND VGND VPWR VPWR _1087_/D sky130_fd_sc_hd__dfxtp_1
X_0037_ _0169_/CLK _0037_/D VGND VGND VPWR VPWR _0038_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_21_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1988_ _1991_/CLK _1988_/D VGND VGND VPWR VPWR _1989_/D sky130_fd_sc_hd__dfxtp_1
X_0939_ _1077_/CLK _0939_/D VGND VGND VPWR VPWR _0940_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_106_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_5_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_4_5_0_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1911_ _1918_/CLK _1911_/D VGND VGND VPWR VPWR _1912_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1842_ _1862_/CLK _1842_/D VGND VGND VPWR VPWR _1843_/D sky130_fd_sc_hd__dfxtp_1
X_1773_ _1788_/CLK _1773_/D VGND VGND VPWR VPWR _1774_/D sky130_fd_sc_hd__dfxtp_1
X_0724_ _0791_/CLK _0724_/D VGND VGND VPWR VPWR _0725_/D sky130_fd_sc_hd__dfxtp_1
X_0655_ _0916_/CLK _0655_/D VGND VGND VPWR VPWR _0656_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_89_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0586_ _0595_/CLK _0586_/D VGND VGND VPWR VPWR _0587_/D sky130_fd_sc_hd__dfxtp_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1207_ _1233_/CLK _1207_/D VGND VGND VPWR VPWR _1208_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_53_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1138_ _1138_/CLK _1138_/D VGND VGND VPWR VPWR _1139_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1069_ _1071_/CLK _1069_/D VGND VGND VPWR VPWR _1070_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_13_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0440_ _0539_/CLK _0440_/D VGND VGND VPWR VPWR _0451_/D sky130_fd_sc_hd__dfxtp_1
X_0371_ _1112_/CLK _0371_/D VGND VGND VPWR VPWR _0372_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_39_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1825_ _1826_/CLK _1825_/D VGND VGND VPWR VPWR _1826_/D sky130_fd_sc_hd__dfxtp_1
X_1756_ _1833_/CLK input1/X VGND VGND VPWR VPWR _1767_/D sky130_fd_sc_hd__dfxtp_1
X_0707_ _0813_/CLK _0707_/D VGND VGND VPWR VPWR _0708_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_104_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1687_ _1687_/CLK _1687_/D VGND VGND VPWR VPWR _1688_/D sky130_fd_sc_hd__dfxtp_1
X_0638_ _1649_/CLK _0638_/D VGND VGND VPWR VPWR _0649_/D sky130_fd_sc_hd__dfxtp_1
X_0569_ _0595_/CLK _0569_/D VGND VGND VPWR VPWR _0570_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_97_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1610_ _1987_/CLK _1610_/D VGND VGND VPWR VPWR _1611_/D sky130_fd_sc_hd__dfxtp_1
X_1541_ _1578_/CLK _1541_/D VGND VGND VPWR VPWR _1542_/D sky130_fd_sc_hd__dfxtp_1
X_1472_ _1726_/CLK _1472_/D VGND VGND VPWR VPWR _1473_/D sky130_fd_sc_hd__dfxtp_1
X_0423_ _0622_/CLK _0423_/D VGND VGND VPWR VPWR _0424_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0354_ _1112_/CLK _0354_/D VGND VGND VPWR VPWR _0355_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_94_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0285_ _1033_/CLK _0285_/D VGND VGND VPWR VPWR _0287_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_82_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1808_ _1808_/CLK _1808_/D VGND VGND VPWR VPWR _1809_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1739_ _1747_/CLK _1739_/D VGND VGND VPWR VPWR _1740_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0070_ _1816_/CLK _0070_/D VGND VGND VPWR VPWR _0071_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_17_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0972_ _0977_/CLK _0972_/D VGND VGND VPWR VPWR _0973_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1524_ _1587_/CLK _1524_/D VGND VGND VPWR VPWR _1525_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1455_ _1710_/CLK _1455_/D VGND VGND VPWR VPWR _1456_/D sky130_fd_sc_hd__dfxtp_1
X_0406_ _0622_/CLK _0406_/D VGND VGND VPWR VPWR _0408_/D sky130_fd_sc_hd__dfxtp_1
X_1386_ _1764_/CLK _1386_/D VGND VGND VPWR VPWR _1387_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_28_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0337_ _1070_/CLK _0337_/D VGND VGND VPWR VPWR _0338_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_55_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0268_ _0280_/CLK _0268_/D VGND VGND VPWR VPWR _0269_/D sky130_fd_sc_hd__dfxtp_1
X_0199_ _1178_/CLK _0199_/D VGND VGND VPWR VPWR _0200_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_23_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1240_ _1244_/CLK _1240_/D VGND VGND VPWR VPWR _1241_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1171_ _1180_/CLK _1171_/D VGND VGND VPWR VPWR _1172_/D sky130_fd_sc_hd__dfxtp_1
X_0122_ _1138_/CLK _0122_/D VGND VGND VPWR VPWR _0123_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0053_ _1841_/CLK _0053_/D VGND VGND VPWR VPWR _0054_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0955_ _0966_/CLK _0955_/D VGND VGND VPWR VPWR _0956_/D sky130_fd_sc_hd__dfxtp_1
X_0886_ _0916_/CLK _0886_/D VGND VGND VPWR VPWR _0887_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_121_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _1364_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_101_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1507_ _1604_/CLK _1507_/D VGND VGND VPWR VPWR _1508_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1438_ _1814_/CLK _1438_/D VGND VGND VPWR VPWR _1439_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1369_ _1373_/CLK _1369_/D VGND VGND VPWR VPWR _1370_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_112_clk clkbuf_4_1_0_clk/X VGND VGND VPWR VPWR _1710_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_3_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_103_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _1665_/CLK sky130_fd_sc_hd__clkbuf_16
X_0740_ _1138_/CLK _0740_/D VGND VGND VPWR VPWR _0741_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_10_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0671_ _1665_/CLK _0671_/D VGND VGND VPWR VPWR _0682_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1223_ _1228_/CLK _1223_/D VGND VGND VPWR VPWR _1224_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1154_ _1163_/CLK _1154_/D VGND VGND VPWR VPWR _1156_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1085_ _1088_/CLK _1085_/D VGND VGND VPWR VPWR _1086_/D sky130_fd_sc_hd__dfxtp_1
X_0105_ _0750_/CLK _0105_/D VGND VGND VPWR VPWR _0106_/D sky130_fd_sc_hd__dfxtp_1
X_0036_ _1846_/CLK _0036_/D VGND VGND VPWR VPWR _0037_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1987_ _1987_/CLK _1987_/D VGND VGND VPWR VPWR _1987_/Q sky130_fd_sc_hd__dfxtp_1
X_0938_ _1077_/CLK _0938_/D VGND VGND VPWR VPWR _0939_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0869_ _1665_/CLK _0869_/D VGND VGND VPWR VPWR _0880_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_88_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1910_ _1987_/CLK _1910_/D VGND VGND VPWR VPWR _1921_/D sky130_fd_sc_hd__dfxtp_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1841_ _1841_/CLK _1841_/D VGND VGND VPWR VPWR _1842_/D sky130_fd_sc_hd__dfxtp_1
X_1772_ _1772_/CLK _1772_/D VGND VGND VPWR VPWR _1773_/D sky130_fd_sc_hd__dfxtp_1
X_0723_ _0791_/CLK _0723_/D VGND VGND VPWR VPWR _0724_/D sky130_fd_sc_hd__dfxtp_1
X_0654_ _0916_/CLK _0654_/D VGND VGND VPWR VPWR _0655_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_6_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0585_ _0585_/CLK _0585_/D VGND VGND VPWR VPWR _0586_/D sky130_fd_sc_hd__dfxtp_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1206_ _1233_/CLK _1206_/D VGND VGND VPWR VPWR _1207_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1137_ _1147_/CLK _1137_/D VGND VGND VPWR VPWR _1138_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_65_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1068_ _1071_/CLK _1068_/D VGND VGND VPWR VPWR _1069_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_33_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0019_ _1858_/CLK _0019_/D VGND VGND VPWR VPWR _0020_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0370_ _1112_/CLK _0370_/D VGND VGND VPWR VPWR _0371_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_4_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_4_4_0_clk/X sky130_fd_sc_hd__clkbuf_1
X_1824_ _1846_/CLK _1824_/D VGND VGND VPWR VPWR _1825_/D sky130_fd_sc_hd__dfxtp_1
X_1755_ _1783_/CLK _1755_/D VGND VGND VPWR VPWR _1757_/D sky130_fd_sc_hd__dfxtp_1
X_0706_ _1127_/CLK _0706_/D VGND VGND VPWR VPWR _0707_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_7_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1686_ _1686_/CLK _1686_/D VGND VGND VPWR VPWR _1687_/D sky130_fd_sc_hd__dfxtp_1
X_0637_ _0642_/CLK _0637_/D VGND VGND VPWR VPWR _0639_/D sky130_fd_sc_hd__dfxtp_1
X_0568_ _0595_/CLK _0568_/D VGND VGND VPWR VPWR _0569_/D sky130_fd_sc_hd__dfxtp_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0499_ _0508_/CLK _0499_/D VGND VGND VPWR VPWR _0500_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_38_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_92_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _1604_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_38_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_83_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _1975_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1540_ _1578_/CLK _1540_/D VGND VGND VPWR VPWR _1541_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1471_ _1673_/CLK _1471_/D VGND VGND VPWR VPWR _1472_/D sky130_fd_sc_hd__dfxtp_1
X_0422_ _0953_/CLK _0422_/D VGND VGND VPWR VPWR _0423_/D sky130_fd_sc_hd__dfxtp_1
X_0353_ _1088_/CLK _0353_/D VGND VGND VPWR VPWR _0354_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0284_ _1980_/CLK _0284_/D VGND VGND VPWR VPWR _0285_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_94_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_74_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _1996_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1807_ _1814_/CLK _1807_/D VGND VGND VPWR VPWR _1808_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_104_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1738_ _1747_/CLK _1738_/D VGND VGND VPWR VPWR _1739_/D sky130_fd_sc_hd__dfxtp_1
X_1669_ _1673_/CLK _1669_/D VGND VGND VPWR VPWR _1670_/D sky130_fd_sc_hd__dfxtp_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_65_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _1017_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_56_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _0973_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0971_ _1039_/CLK _0971_/D VGND VGND VPWR VPWR _0972_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_9_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1523_ _1587_/CLK _1523_/D VGND VGND VPWR VPWR _1524_/D sky130_fd_sc_hd__dfxtp_1
X_1454_ _1695_/CLK _1454_/D VGND VGND VPWR VPWR _1455_/D sky130_fd_sc_hd__dfxtp_1
X_0405_ _0622_/CLK _0405_/D VGND VGND VPWR VPWR _0406_/D sky130_fd_sc_hd__dfxtp_1
X_1385_ _1764_/CLK _1385_/D VGND VGND VPWR VPWR _1386_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0336_ _1070_/CLK _0336_/D VGND VGND VPWR VPWR _0337_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_27_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0267_ _0280_/CLK _0267_/D VGND VGND VPWR VPWR _0268_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_47_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _1071_/CLK sky130_fd_sc_hd__clkbuf_16
X_0198_ _1594_/CLK _0198_/D VGND VGND VPWR VPWR _0209_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_38_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _0932_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1170_ _1170_/CLK _1170_/D VGND VGND VPWR VPWR _1171_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0121_ _1635_/CLK _0121_/D VGND VGND VPWR VPWR _0132_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_29_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _0864_/CLK sky130_fd_sc_hd__clkbuf_16
X_0052_ _1185_/CLK _0052_/D VGND VGND VPWR VPWR _0053_/D sky130_fd_sc_hd__dfxtp_1
X_0954_ _0966_/CLK _0954_/D VGND VGND VPWR VPWR _0955_/D sky130_fd_sc_hd__dfxtp_1
X_0885_ _0894_/CLK _0885_/D VGND VGND VPWR VPWR _0886_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1506_ _1604_/CLK _1506_/D VGND VGND VPWR VPWR _1507_/D sky130_fd_sc_hd__dfxtp_1
X_1437_ _1814_/CLK _1437_/D VGND VGND VPWR VPWR _1438_/D sky130_fd_sc_hd__dfxtp_1
X_1368_ _1373_/CLK _1368_/D VGND VGND VPWR VPWR _1369_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0319_ _0539_/CLK _0319_/D VGND VGND VPWR VPWR _0330_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1299_ _1302_/CLK _1299_/D VGND VGND VPWR VPWR _1300_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0670_ _0874_/CLK _0670_/D VGND VGND VPWR VPWR _0672_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_10_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1222_ _1229_/CLK _1222_/D VGND VGND VPWR VPWR _1223_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1153_ _1163_/CLK _1153_/D VGND VGND VPWR VPWR _1154_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1084_ _1088_/CLK _1084_/D VGND VGND VPWR VPWR _1085_/D sky130_fd_sc_hd__dfxtp_1
X_0104_ _0750_/CLK _0104_/D VGND VGND VPWR VPWR _0105_/D sky130_fd_sc_hd__dfxtp_1
X_0035_ _1858_/CLK _0035_/D VGND VGND VPWR VPWR _0036_/D sky130_fd_sc_hd__dfxtp_1
X_1986_ _1991_/CLK _1986_/D VGND VGND VPWR VPWR _1988_/D sky130_fd_sc_hd__dfxtp_1
X_0937_ _0953_/CLK _0937_/D VGND VGND VPWR VPWR _0938_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_9_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _1233_/CLK sky130_fd_sc_hd__clkbuf_16
X_0868_ _0874_/CLK _0868_/D VGND VGND VPWR VPWR _0870_/D sky130_fd_sc_hd__dfxtp_1
X_0799_ _0813_/CLK _0799_/D VGND VGND VPWR VPWR _0800_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_88_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1840_ _1846_/CLK _1840_/D VGND VGND VPWR VPWR _1841_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1771_ _1772_/CLK _1771_/D VGND VGND VPWR VPWR _1772_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_6_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0722_ _0791_/CLK _0722_/D VGND VGND VPWR VPWR _0723_/D sky130_fd_sc_hd__dfxtp_1
X_0653_ _0916_/CLK _0653_/D VGND VGND VPWR VPWR _0654_/D sky130_fd_sc_hd__dfxtp_1
X_0584_ _0973_/CLK _0584_/D VGND VGND VPWR VPWR _0585_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1205_ _1808_/CLK _1205_/D VGND VGND VPWR VPWR _1206_/D sky130_fd_sc_hd__dfxtp_1
X_1136_ _1138_/CLK _1136_/D VGND VGND VPWR VPWR _1137_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1067_ _1826_/CLK _1067_/D VGND VGND VPWR VPWR _1078_/D sky130_fd_sc_hd__dfxtp_1
X_0018_ _1858_/CLK _0018_/D VGND VGND VPWR VPWR _0019_/D sky130_fd_sc_hd__dfxtp_1
X_1969_ _1973_/CLK _1969_/D VGND VGND VPWR VPWR _1970_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1823_ _1826_/CLK _1823_/D VGND VGND VPWR VPWR _1824_/D sky130_fd_sc_hd__dfxtp_1
X_1754_ _1754_/CLK _1754_/D VGND VGND VPWR VPWR _1755_/D sky130_fd_sc_hd__dfxtp_1
X_0705_ _0813_/CLK _0705_/D VGND VGND VPWR VPWR _0706_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_104_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1685_ _1686_/CLK _1685_/D VGND VGND VPWR VPWR _1686_/D sky130_fd_sc_hd__dfxtp_1
X_0636_ _0642_/CLK _0636_/D VGND VGND VPWR VPWR _0637_/D sky130_fd_sc_hd__dfxtp_1
X_0567_ _0595_/CLK _0567_/D VGND VGND VPWR VPWR _0568_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_97_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0498_ _0508_/CLK _0498_/D VGND VGND VPWR VPWR _0499_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1119_ _1163_/CLK _1119_/D VGND VGND VPWR VPWR _1120_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1470_ _1726_/CLK _1470_/D VGND VGND VPWR VPWR _1471_/D sky130_fd_sc_hd__dfxtp_1
X_0421_ _0953_/CLK _0421_/D VGND VGND VPWR VPWR _0422_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_79_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0352_ _1907_/CLK _0352_/D VGND VGND VPWR VPWR _0363_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_94_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0283_ _1033_/CLK _0283_/D VGND VGND VPWR VPWR _0284_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_90_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1806_ _1808_/CLK _1806_/D VGND VGND VPWR VPWR _1807_/D sky130_fd_sc_hd__dfxtp_1
X_1737_ _1747_/CLK _1737_/D VGND VGND VPWR VPWR _1738_/D sky130_fd_sc_hd__dfxtp_1
X_1668_ _1687_/CLK _1668_/D VGND VGND VPWR VPWR _1669_/D sky130_fd_sc_hd__dfxtp_1
X_0619_ _0632_/CLK _0619_/D VGND VGND VPWR VPWR _0620_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_100_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1599_ _1600_/CLK _1599_/D VGND VGND VPWR VPWR _1600_/D sky130_fd_sc_hd__dfxtp_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_3_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_4_3_0_clk/X sky130_fd_sc_hd__clkbuf_1
X_0970_ _1046_/CLK _0970_/D VGND VGND VPWR VPWR _0971_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1522_ _1587_/CLK _1522_/D VGND VGND VPWR VPWR _1523_/D sky130_fd_sc_hd__dfxtp_1
X_1453_ _1695_/CLK _1453_/D VGND VGND VPWR VPWR _1454_/D sky130_fd_sc_hd__dfxtp_1
X_0404_ _0642_/CLK _0404_/D VGND VGND VPWR VPWR _0405_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1384_ _1764_/CLK _1384_/D VGND VGND VPWR VPWR _1385_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0335_ _1070_/CLK _0335_/D VGND VGND VPWR VPWR _0336_/D sky130_fd_sc_hd__dfxtp_1
X_0266_ _0280_/CLK _0266_/D VGND VGND VPWR VPWR _0267_/D sky130_fd_sc_hd__dfxtp_1
X_0197_ _1178_/CLK _0197_/D VGND VGND VPWR VPWR _0199_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_63_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0120_ _1138_/CLK _0120_/D VGND VGND VPWR VPWR _0122_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0051_ _0169_/CLK _0051_/D VGND VGND VPWR VPWR _0052_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0953_ _0953_/CLK _0953_/D VGND VGND VPWR VPWR _0954_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0884_ _0894_/CLK _0884_/D VGND VGND VPWR VPWR _0885_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1505_ _1604_/CLK _1505_/D VGND VGND VPWR VPWR _1506_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_87_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1436_ _1814_/CLK _1436_/D VGND VGND VPWR VPWR _1437_/D sky130_fd_sc_hd__dfxtp_1
X_1367_ _1373_/CLK _1367_/D VGND VGND VPWR VPWR _1368_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0318_ _1055_/CLK _0318_/D VGND VGND VPWR VPWR _0320_/D sky130_fd_sc_hd__dfxtp_1
X_1298_ _1302_/CLK _1298_/D VGND VGND VPWR VPWR _1299_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0249_ _1980_/CLK _0249_/D VGND VGND VPWR VPWR _0250_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1221_ _1816_/CLK _1221_/D VGND VGND VPWR VPWR _1222_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_65_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1152_ _1163_/CLK _1152_/D VGND VGND VPWR VPWR _1153_/D sky130_fd_sc_hd__dfxtp_1
X_1083_ _1181_/CLK _1083_/D VGND VGND VPWR VPWR _1084_/D sky130_fd_sc_hd__dfxtp_1
X_0103_ _1226_/CLK _0103_/D VGND VGND VPWR VPWR _0104_/D sky130_fd_sc_hd__dfxtp_1
X_0034_ _1846_/CLK _0034_/D VGND VGND VPWR VPWR _0035_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1985_ _1985_/CLK _1985_/D VGND VGND VPWR VPWR _1986_/D sky130_fd_sc_hd__dfxtp_1
X_0936_ _1077_/CLK _0936_/D VGND VGND VPWR VPWR _0937_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0867_ _0874_/CLK _0867_/D VGND VGND VPWR VPWR _0868_/D sky130_fd_sc_hd__dfxtp_1
X_0798_ _0813_/CLK _0798_/D VGND VGND VPWR VPWR _0799_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_87_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1419_ _1783_/CLK _1419_/D VGND VGND VPWR VPWR _1420_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1770_ _1788_/CLK _1770_/D VGND VGND VPWR VPWR _1771_/D sky130_fd_sc_hd__dfxtp_1
X_0721_ _1127_/CLK _0721_/D VGND VGND VPWR VPWR _0722_/D sky130_fd_sc_hd__dfxtp_1
X_0652_ _0919_/CLK _0652_/D VGND VGND VPWR VPWR _0653_/D sky130_fd_sc_hd__dfxtp_1
X_0583_ _1649_/CLK _0583_/D VGND VGND VPWR VPWR _0594_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1204_ _1808_/CLK _1204_/D VGND VGND VPWR VPWR _1205_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_65_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1135_ _1147_/CLK _1135_/D VGND VGND VPWR VPWR _1136_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_65_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1066_ _1071_/CLK _1066_/D VGND VGND VPWR VPWR _1068_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_21_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0017_ _0214_/CLK _0017_/D VGND VGND VPWR VPWR _0018_/D sky130_fd_sc_hd__dfxtp_1
X_1968_ _1975_/CLK _1968_/D VGND VGND VPWR VPWR _1969_/D sky130_fd_sc_hd__dfxtp_1
X_0919_ _0919_/CLK _0919_/D VGND VGND VPWR VPWR _0920_/D sky130_fd_sc_hd__dfxtp_1
X_1899_ _1987_/CLK _1899_/D VGND VGND VPWR VPWR _1910_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_88_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1822_ _1987_/CLK _1822_/D VGND VGND VPWR VPWR _1833_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1753_ _1772_/CLK _1753_/D VGND VGND VPWR VPWR _1754_/D sky130_fd_sc_hd__dfxtp_1
X_1684_ _1686_/CLK _1684_/D VGND VGND VPWR VPWR _1685_/D sky130_fd_sc_hd__dfxtp_1
X_0704_ _1665_/CLK _0704_/D VGND VGND VPWR VPWR _0715_/D sky130_fd_sc_hd__dfxtp_1
X_0635_ _0642_/CLK _0635_/D VGND VGND VPWR VPWR _0636_/D sky130_fd_sc_hd__dfxtp_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0566_ _0595_/CLK _0566_/D VGND VGND VPWR VPWR _0567_/D sky130_fd_sc_hd__dfxtp_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0497_ _0508_/CLK _0497_/D VGND VGND VPWR VPWR _0498_/D sky130_fd_sc_hd__dfxtp_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1118_ _1163_/CLK _1118_/D VGND VGND VPWR VPWR _1119_/D sky130_fd_sc_hd__dfxtp_1
X_1049_ _1055_/CLK _1049_/D VGND VGND VPWR VPWR _1050_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0420_ _0953_/CLK _0420_/D VGND VGND VPWR VPWR _0421_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0351_ _1088_/CLK _0351_/D VGND VGND VPWR VPWR _0353_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0282_ _0295_/CLK _0282_/D VGND VGND VPWR VPWR _0283_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_90_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1805_ _1808_/CLK _1805_/D VGND VGND VPWR VPWR _1806_/D sky130_fd_sc_hd__dfxtp_1
X_1736_ _1736_/CLK _1736_/D VGND VGND VPWR VPWR _1737_/D sky130_fd_sc_hd__dfxtp_1
X_1667_ _1687_/CLK _1667_/D VGND VGND VPWR VPWR _1668_/D sky130_fd_sc_hd__dfxtp_1
X_0618_ _0632_/CLK _0618_/D VGND VGND VPWR VPWR _0619_/D sky130_fd_sc_hd__dfxtp_1
X_1598_ _1600_/CLK _1598_/D VGND VGND VPWR VPWR _1599_/D sky130_fd_sc_hd__dfxtp_1
X_0549_ _0573_/CLK _0549_/D VGND VGND VPWR VPWR _0551_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1521_ _1587_/CLK _1521_/D VGND VGND VPWR VPWR _1522_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1452_ _1695_/CLK _1452_/D VGND VGND VPWR VPWR _1453_/D sky130_fd_sc_hd__dfxtp_1
X_0403_ _0622_/CLK _0403_/D VGND VGND VPWR VPWR _0404_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1383_ _1764_/CLK _1383_/D VGND VGND VPWR VPWR _1384_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0334_ _1070_/CLK _0334_/D VGND VGND VPWR VPWR _0335_/D sky130_fd_sc_hd__dfxtp_1
X_0265_ _0280_/CLK _0265_/D VGND VGND VPWR VPWR _0266_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_82_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0196_ _0214_/CLK _0196_/D VGND VGND VPWR VPWR _0197_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_90_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1719_ _1833_/CLK _1719_/D VGND VGND VPWR VPWR _1720_/D sky130_fd_sc_hd__dfxtp_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_115_clk clkbuf_4_1_0_clk/X VGND VGND VPWR VPWR _1754_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0050_ _1841_/CLK _0050_/D VGND VGND VPWR VPWR _0051_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_17_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0952_ _0953_/CLK _0952_/D VGND VGND VPWR VPWR _0953_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_106_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _1846_/CLK sky130_fd_sc_hd__clkbuf_16
X_0883_ _0894_/CLK _0883_/D VGND VGND VPWR VPWR _0884_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1504_ _1604_/CLK _1504_/D VGND VGND VPWR VPWR _1505_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_102_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1435_ _1814_/CLK _1435_/D VGND VGND VPWR VPWR _1436_/D sky130_fd_sc_hd__dfxtp_1
X_1366_ _1373_/CLK _1366_/D VGND VGND VPWR VPWR _1367_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0317_ _1055_/CLK _0317_/D VGND VGND VPWR VPWR _0318_/D sky130_fd_sc_hd__dfxtp_1
X_1297_ _1348_/CLK _1297_/D VGND VGND VPWR VPWR _1298_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0248_ _1980_/CLK _0248_/D VGND VGND VPWR VPWR _0249_/D sky130_fd_sc_hd__dfxtp_1
X_0179_ _1178_/CLK _0179_/D VGND VGND VPWR VPWR _0180_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_2_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_4_2_0_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1220_ _1228_/CLK _1220_/D VGND VGND VPWR VPWR _1221_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_77_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1151_ _1163_/CLK _1151_/D VGND VGND VPWR VPWR _1152_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0102_ _1226_/CLK _0102_/D VGND VGND VPWR VPWR _0103_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1082_ _1181_/CLK _1082_/D VGND VGND VPWR VPWR _1083_/D sky130_fd_sc_hd__dfxtp_1
X_0033_ _1635_/CLK _0033_/D VGND VGND VPWR VPWR _0044_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_33_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1984_ _1991_/CLK _1984_/D VGND VGND VPWR VPWR _1985_/D sky130_fd_sc_hd__dfxtp_1
X_0935_ _1826_/CLK _0935_/D VGND VGND VPWR VPWR _0946_/D sky130_fd_sc_hd__dfxtp_1
X_0866_ _0874_/CLK _0866_/D VGND VGND VPWR VPWR _0867_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_106_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0797_ _0813_/CLK _0797_/D VGND VGND VPWR VPWR _0798_/D sky130_fd_sc_hd__dfxtp_1
X_1418_ _1783_/CLK _1418_/D VGND VGND VPWR VPWR _1419_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1349_ _1373_/CLK _1349_/D VGND VGND VPWR VPWR _1350_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_56_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0720_ _0793_/CLK _0720_/D VGND VGND VPWR VPWR _0721_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0651_ _0919_/CLK _0651_/D VGND VGND VPWR VPWR _0652_/D sky130_fd_sc_hd__dfxtp_1
X_0582_ _0595_/CLK _0582_/D VGND VGND VPWR VPWR _0584_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_97_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1203_ _1808_/CLK _1203_/D VGND VGND VPWR VPWR _1204_/D sky130_fd_sc_hd__dfxtp_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1134_ _1147_/CLK _1134_/D VGND VGND VPWR VPWR _1135_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1065_ _1071_/CLK _1065_/D VGND VGND VPWR VPWR _1066_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_18_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0016_ _0214_/CLK _0016_/D VGND VGND VPWR VPWR _0017_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_21_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1967_ _1973_/CLK _1967_/D VGND VGND VPWR VPWR _1968_/D sky130_fd_sc_hd__dfxtp_1
X_0918_ _0919_/CLK _0918_/D VGND VGND VPWR VPWR _0919_/D sky130_fd_sc_hd__dfxtp_1
X_1898_ _1985_/CLK _1898_/D VGND VGND VPWR VPWR _1900_/D sky130_fd_sc_hd__dfxtp_1
X_0849_ _0874_/CLK _0849_/D VGND VGND VPWR VPWR _0850_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_95_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _1635_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_86_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _1918_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1821_ _1826_/CLK _1821_/D VGND VGND VPWR VPWR _1823_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1752_ _1783_/CLK _1752_/D VGND VGND VPWR VPWR _1753_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_10_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _1808_/CLK sky130_fd_sc_hd__clkbuf_16
X_0703_ _0906_/CLK _0703_/D VGND VGND VPWR VPWR _0705_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_7_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1683_ _1687_/CLK _1683_/D VGND VGND VPWR VPWR _1684_/D sky130_fd_sc_hd__dfxtp_1
X_0634_ _0642_/CLK _0634_/D VGND VGND VPWR VPWR _0635_/D sky130_fd_sc_hd__dfxtp_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0565_ _0595_/CLK _0565_/D VGND VGND VPWR VPWR _0566_/D sky130_fd_sc_hd__dfxtp_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0496_ _0998_/CLK _0496_/D VGND VGND VPWR VPWR _0497_/D sky130_fd_sc_hd__dfxtp_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_77_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _1997_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1117_ _1127_/CLK _1117_/D VGND VGND VPWR VPWR _1118_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1048_ _1055_/CLK _1048_/D VGND VGND VPWR VPWR _1049_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_21_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_68_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _1973_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0350_ _1088_/CLK _0350_/D VGND VGND VPWR VPWR _0351_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_94_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0281_ _1033_/CLK _0281_/D VGND VGND VPWR VPWR _0282_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_59_clk clkbuf_4_15_0_clk/X VGND VGND VPWR VPWR _1182_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_85_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1804_ _1814_/CLK _1804_/D VGND VGND VPWR VPWR _1805_/D sky130_fd_sc_hd__dfxtp_1
X_1735_ _1736_/CLK _1735_/D VGND VGND VPWR VPWR _1736_/D sky130_fd_sc_hd__dfxtp_1
X_1666_ _1673_/CLK _1666_/D VGND VGND VPWR VPWR _1667_/D sky130_fd_sc_hd__dfxtp_1
X_0617_ _0632_/CLK _0617_/D VGND VGND VPWR VPWR _0618_/D sky130_fd_sc_hd__dfxtp_1
X_1597_ _1600_/CLK _1597_/D VGND VGND VPWR VPWR _1598_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0548_ _0573_/CLK _0548_/D VGND VGND VPWR VPWR _0549_/D sky130_fd_sc_hd__dfxtp_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0479_ _0998_/CLK _0479_/D VGND VGND VPWR VPWR _0480_/D sky130_fd_sc_hd__dfxtp_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1520_ _1587_/CLK _1520_/D VGND VGND VPWR VPWR _1521_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1451_ _1695_/CLK _1451_/D VGND VGND VPWR VPWR _1452_/D sky130_fd_sc_hd__dfxtp_1
X_0402_ _0642_/CLK _0402_/D VGND VGND VPWR VPWR _0403_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1382_ _1764_/CLK _1382_/D VGND VGND VPWR VPWR _1383_/D sky130_fd_sc_hd__dfxtp_1
X_0333_ _1070_/CLK _0333_/D VGND VGND VPWR VPWR _0334_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0264_ _0539_/CLK _0264_/D VGND VGND VPWR VPWR _0275_/D sky130_fd_sc_hd__dfxtp_1
X_0195_ _0214_/CLK _0195_/D VGND VGND VPWR VPWR _0196_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1718_ _1833_/CLK _1718_/D VGND VGND VPWR VPWR _1719_/D sky130_fd_sc_hd__dfxtp_1
X_1649_ _1649_/CLK _1649_/D VGND VGND VPWR VPWR _1650_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0951_ _0966_/CLK _0951_/D VGND VGND VPWR VPWR _0952_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0882_ _0894_/CLK _0882_/D VGND VGND VPWR VPWR _0883_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_9_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1503_ _1604_/CLK _1503_/D VGND VGND VPWR VPWR _1504_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1434_ _1814_/CLK _1434_/D VGND VGND VPWR VPWR _1435_/D sky130_fd_sc_hd__dfxtp_1
X_1365_ _1373_/CLK _1365_/D VGND VGND VPWR VPWR _1366_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0316_ _0316_/CLK _0316_/D VGND VGND VPWR VPWR _0317_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1296_ _1348_/CLK _1296_/D VGND VGND VPWR VPWR _1297_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0247_ _0295_/CLK _0247_/D VGND VGND VPWR VPWR _0248_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0178_ _1180_/CLK _0178_/D VGND VGND VPWR VPWR _0179_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_11_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1150_ _1163_/CLK _1150_/D VGND VGND VPWR VPWR _1151_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0101_ _1226_/CLK _0101_/D VGND VGND VPWR VPWR _0102_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_65_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1081_ _1104_/CLK _1081_/D VGND VGND VPWR VPWR _1082_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0032_ _1846_/CLK _0032_/D VGND VGND VPWR VPWR _0034_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_33_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1983_ _1991_/CLK _1983_/D VGND VGND VPWR VPWR _1984_/D sky130_fd_sc_hd__dfxtp_1
X_0934_ _1077_/CLK _0934_/D VGND VGND VPWR VPWR _0936_/D sky130_fd_sc_hd__dfxtp_1
X_0865_ _0874_/CLK _0865_/D VGND VGND VPWR VPWR _0866_/D sky130_fd_sc_hd__dfxtp_1
X_0796_ _0813_/CLK _0796_/D VGND VGND VPWR VPWR _0797_/D sky130_fd_sc_hd__dfxtp_1
X_1417_ _1783_/CLK _1417_/D VGND VGND VPWR VPWR _1418_/D sky130_fd_sc_hd__dfxtp_1
X_1348_ _1348_/CLK _1348_/D VGND VGND VPWR VPWR _1349_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1279_ _1348_/CLK _1279_/D VGND VGND VPWR VPWR _1280_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0650_ _0916_/CLK _0650_/D VGND VGND VPWR VPWR _0651_/D sky130_fd_sc_hd__dfxtp_1
X_0581_ _0585_/CLK _0581_/D VGND VGND VPWR VPWR _0582_/D sky130_fd_sc_hd__dfxtp_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1202_ _1233_/CLK _1202_/D VGND VGND VPWR VPWR _1203_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_1_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_4_1_0_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1133_ _1841_/CLK _1133_/D VGND VGND VPWR VPWR _1144_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_53_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1064_ _1071_/CLK _1064_/D VGND VGND VPWR VPWR _1065_/D sky130_fd_sc_hd__dfxtp_1
X_0015_ _1996_/CLK _0015_/D VGND VGND VPWR VPWR _0016_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_33_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1966_ _1975_/CLK _1966_/D VGND VGND VPWR VPWR _1967_/D sky130_fd_sc_hd__dfxtp_1
X_0917_ _0919_/CLK _0917_/D VGND VGND VPWR VPWR _0918_/D sky130_fd_sc_hd__dfxtp_1
X_1897_ _1975_/CLK _1897_/D VGND VGND VPWR VPWR _1898_/D sky130_fd_sc_hd__dfxtp_1
X_0848_ _0864_/CLK _0848_/D VGND VGND VPWR VPWR _0849_/D sky130_fd_sc_hd__dfxtp_1
X_0779_ _0831_/CLK _0779_/D VGND VGND VPWR VPWR _0780_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1820_ _1826_/CLK _1820_/D VGND VGND VPWR VPWR _1821_/D sky130_fd_sc_hd__dfxtp_1
X_1751_ _1783_/CLK _1751_/D VGND VGND VPWR VPWR _1752_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0702_ _0813_/CLK _0702_/D VGND VGND VPWR VPWR _0703_/D sky130_fd_sc_hd__dfxtp_1
X_1682_ _1827_/CLK _1682_/D VGND VGND VPWR VPWR _1683_/D sky130_fd_sc_hd__dfxtp_1
X_0633_ _0642_/CLK _0633_/D VGND VGND VPWR VPWR _0634_/D sky130_fd_sc_hd__dfxtp_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0564_ _0595_/CLK _0564_/D VGND VGND VPWR VPWR _0565_/D sky130_fd_sc_hd__dfxtp_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0495_ _0539_/CLK _0495_/D VGND VGND VPWR VPWR _0506_/D sky130_fd_sc_hd__dfxtp_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1116_ _1127_/CLK _1116_/D VGND VGND VPWR VPWR _1117_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1047_ _1055_/CLK _1047_/D VGND VGND VPWR VPWR _1048_/D sky130_fd_sc_hd__dfxtp_1
X_1949_ _1956_/CLK _1949_/D VGND VGND VPWR VPWR _1950_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_103_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0280_ _0280_/CLK _0280_/D VGND VGND VPWR VPWR _0281_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_94_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1803_ _1808_/CLK _1803_/D VGND VGND VPWR VPWR _1804_/D sky130_fd_sc_hd__dfxtp_1
X_1734_ _1736_/CLK _1734_/D VGND VGND VPWR VPWR _1735_/D sky130_fd_sc_hd__dfxtp_1
X_1665_ _1665_/CLK _1665_/D VGND VGND VPWR VPWR _1666_/D sky130_fd_sc_hd__dfxtp_1
X_1596_ _1600_/CLK _1596_/D VGND VGND VPWR VPWR _1597_/D sky130_fd_sc_hd__dfxtp_1
X_0616_ _1649_/CLK _0616_/D VGND VGND VPWR VPWR _0627_/D sky130_fd_sc_hd__dfxtp_1
X_0547_ _0573_/CLK _0547_/D VGND VGND VPWR VPWR _0548_/D sky130_fd_sc_hd__dfxtp_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0478_ _0977_/CLK _0478_/D VGND VGND VPWR VPWR _0479_/D sky130_fd_sc_hd__dfxtp_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1450_ _1695_/CLK _1450_/D VGND VGND VPWR VPWR _1451_/D sky130_fd_sc_hd__dfxtp_1
X_0401_ _0622_/CLK _0401_/D VGND VGND VPWR VPWR _0402_/D sky130_fd_sc_hd__dfxtp_1
X_1381_ _1764_/CLK _1381_/D VGND VGND VPWR VPWR _1382_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0332_ _1070_/CLK _0332_/D VGND VGND VPWR VPWR _0333_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0263_ _1973_/CLK _0263_/D VGND VGND VPWR VPWR _0265_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_82_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0194_ _0214_/CLK _0194_/D VGND VGND VPWR VPWR _0195_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_23_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1717_ _1833_/CLK _1717_/D VGND VGND VPWR VPWR _1718_/D sky130_fd_sc_hd__dfxtp_1
X_1648_ _1659_/CLK _1648_/D VGND VGND VPWR VPWR _1649_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1579_ _1592_/CLK _1579_/D VGND VGND VPWR VPWR _1580_/D sky130_fd_sc_hd__dfxtp_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0950_ _0953_/CLK _0950_/D VGND VGND VPWR VPWR _0951_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0881_ _0894_/CLK _0881_/D VGND VGND VPWR VPWR _0882_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_9_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1502_ _1604_/CLK _1502_/D VGND VGND VPWR VPWR _1503_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1433_ _1686_/CLK _1433_/D VGND VGND VPWR VPWR _1434_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1364_ _1364_/CLK _1364_/D VGND VGND VPWR VPWR _1365_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1295_ _1348_/CLK _1295_/D VGND VGND VPWR VPWR _1296_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0315_ _1055_/CLK _0315_/D VGND VGND VPWR VPWR _0316_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0246_ _1980_/CLK _0246_/D VGND VGND VPWR VPWR _0247_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_91_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0177_ _1178_/CLK _0177_/D VGND VGND VPWR VPWR _0178_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_51_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0100_ _1226_/CLK _0100_/D VGND VGND VPWR VPWR _0101_/D sky130_fd_sc_hd__dfxtp_1
X_1080_ _1104_/CLK _1080_/D VGND VGND VPWR VPWR _1081_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0031_ _1858_/CLK _0031_/D VGND VGND VPWR VPWR _0032_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_21_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1982_ _1991_/CLK _1982_/D VGND VGND VPWR VPWR _1983_/D sky130_fd_sc_hd__dfxtp_1
X_0933_ _1077_/CLK _0933_/D VGND VGND VPWR VPWR _0934_/D sky130_fd_sc_hd__dfxtp_1
X_0864_ _0864_/CLK _0864_/D VGND VGND VPWR VPWR _0865_/D sky130_fd_sc_hd__dfxtp_1
X_0795_ _0813_/CLK _0795_/D VGND VGND VPWR VPWR _0796_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_88_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1416_ _1783_/CLK _1416_/D VGND VGND VPWR VPWR _1417_/D sky130_fd_sc_hd__dfxtp_1
X_1347_ _1364_/CLK _1347_/D VGND VGND VPWR VPWR _1348_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1278_ _1348_/CLK _1278_/D VGND VGND VPWR VPWR _1279_/D sky130_fd_sc_hd__dfxtp_1
X_0229_ _1996_/CLK _0229_/D VGND VGND VPWR VPWR _0230_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0580_ _0585_/CLK _0580_/D VGND VGND VPWR VPWR _0581_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_40_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1201_ _1808_/CLK _1201_/D VGND VGND VPWR VPWR _1202_/D sky130_fd_sc_hd__dfxtp_1
X_1132_ _1147_/CLK _1132_/D VGND VGND VPWR VPWR _1134_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1063_ _1071_/CLK _1063_/D VGND VGND VPWR VPWR _1064_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0014_ _1996_/CLK _0014_/D VGND VGND VPWR VPWR _0015_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_33_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1965_ _1965_/CLK _1965_/D VGND VGND VPWR VPWR _1976_/D sky130_fd_sc_hd__dfxtp_1
X_0916_ _0916_/CLK _0916_/D VGND VGND VPWR VPWR _0917_/D sky130_fd_sc_hd__dfxtp_1
X_1896_ _1975_/CLK _1896_/D VGND VGND VPWR VPWR _1897_/D sky130_fd_sc_hd__dfxtp_1
X_0847_ _1827_/CLK _0847_/D VGND VGND VPWR VPWR _0858_/D sky130_fd_sc_hd__dfxtp_1
X_0778_ _0831_/CLK _0778_/D VGND VGND VPWR VPWR _0779_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_88_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1750_ _1754_/CLK _1750_/D VGND VGND VPWR VPWR _1751_/D sky130_fd_sc_hd__dfxtp_1
X_0701_ _0906_/CLK _0701_/D VGND VGND VPWR VPWR _0702_/D sky130_fd_sc_hd__dfxtp_1
X_1681_ _1827_/CLK _1681_/D VGND VGND VPWR VPWR _1682_/D sky130_fd_sc_hd__dfxtp_1
X_0632_ _0632_/CLK _0632_/D VGND VGND VPWR VPWR _0633_/D sky130_fd_sc_hd__dfxtp_1
X_0563_ _0610_/CLK _0563_/D VGND VGND VPWR VPWR _0564_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0494_ _0508_/CLK _0494_/D VGND VGND VPWR VPWR _0496_/D sky130_fd_sc_hd__dfxtp_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1115_ _1163_/CLK _1115_/D VGND VGND VPWR VPWR _1116_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1046_ _1046_/CLK _1046_/D VGND VGND VPWR VPWR _1047_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_61_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1948_ _1975_/CLK _1948_/D VGND VGND VPWR VPWR _1949_/D sky130_fd_sc_hd__dfxtp_1
X_1879_ _1995_/CLK _1879_/D VGND VGND VPWR VPWR _1880_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_0_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_4_0_0_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1802_ _1808_/CLK _1802_/D VGND VGND VPWR VPWR _1803_/D sky130_fd_sc_hd__dfxtp_1
X_1733_ _1736_/CLK _1733_/D VGND VGND VPWR VPWR _1734_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1664_ _1665_/CLK _1664_/D VGND VGND VPWR VPWR _1665_/D sky130_fd_sc_hd__dfxtp_1
X_0615_ _0632_/CLK _0615_/D VGND VGND VPWR VPWR _0617_/D sky130_fd_sc_hd__dfxtp_1
X_1595_ _1600_/CLK _1595_/D VGND VGND VPWR VPWR _1596_/D sky130_fd_sc_hd__dfxtp_1
X_0546_ _0573_/CLK _0546_/D VGND VGND VPWR VPWR _0547_/D sky130_fd_sc_hd__dfxtp_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0477_ _0977_/CLK _0477_/D VGND VGND VPWR VPWR _0478_/D sky130_fd_sc_hd__dfxtp_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1029_ _1033_/CLK _1029_/D VGND VGND VPWR VPWR _1030_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_22_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_118_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _1772_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0400_ _0642_/CLK _0400_/D VGND VGND VPWR VPWR _0401_/D sky130_fd_sc_hd__dfxtp_1
X_1380_ _1764_/CLK _1380_/D VGND VGND VPWR VPWR _1381_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0331_ _1070_/CLK _0331_/D VGND VGND VPWR VPWR _0332_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0262_ _0280_/CLK _0262_/D VGND VGND VPWR VPWR _0263_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0193_ _0214_/CLK _0193_/D VGND VGND VPWR VPWR _0194_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_35_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_109_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _1814_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1716_ _1726_/CLK _1716_/D VGND VGND VPWR VPWR _1717_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_105_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1647_ _1649_/CLK _1647_/D VGND VGND VPWR VPWR _1648_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1578_ _1578_/CLK _1578_/D VGND VGND VPWR VPWR _1579_/D sky130_fd_sc_hd__dfxtp_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0529_ _0529_/CLK _0529_/D VGND VGND VPWR VPWR _0530_/D sky130_fd_sc_hd__dfxtp_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0880_ _1827_/CLK _0880_/D VGND VGND VPWR VPWR _0891_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_40_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1501_ _1604_/CLK _1501_/D VGND VGND VPWR VPWR _1502_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1432_ _1794_/CLK _1432_/D VGND VGND VPWR VPWR _1433_/D sky130_fd_sc_hd__dfxtp_1
X_1363_ _1373_/CLK _1363_/D VGND VGND VPWR VPWR _1364_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1294_ _1336_/CLK _1294_/D VGND VGND VPWR VPWR _1295_/D sky130_fd_sc_hd__dfxtp_1
X_0314_ _0316_/CLK _0314_/D VGND VGND VPWR VPWR _0315_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0245_ _1980_/CLK _0245_/D VGND VGND VPWR VPWR _0246_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0176_ _1600_/CLK _0176_/D VGND VGND VPWR VPWR _0187_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0030_ _1858_/CLK _0030_/D VGND VGND VPWR VPWR _0031_/D sky130_fd_sc_hd__dfxtp_1
X_1981_ _1991_/CLK _1981_/D VGND VGND VPWR VPWR _1982_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_60_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0932_ _0932_/CLK _0932_/D VGND VGND VPWR VPWR _0933_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_40_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _1103_/CLK sky130_fd_sc_hd__clkbuf_16
X_0863_ _0864_/CLK _0863_/D VGND VGND VPWR VPWR _0864_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0794_ _0813_/CLK _0794_/D VGND VGND VPWR VPWR _0795_/D sky130_fd_sc_hd__dfxtp_1
X_1415_ _1783_/CLK _1415_/D VGND VGND VPWR VPWR _1416_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1346_ _1364_/CLK _1346_/D VGND VGND VPWR VPWR _1347_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1277_ _1348_/CLK _1277_/D VGND VGND VPWR VPWR _1278_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0228_ _1996_/CLK _0228_/D VGND VGND VPWR VPWR _0229_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0159_ _0169_/CLK _0159_/D VGND VGND VPWR VPWR _0160_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_24_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_31_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _0894_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_105_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_98_clk clkbuf_4_4_0_clk/X VGND VGND VPWR VPWR _1833_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _0750_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_89_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _1592_/CLK sky130_fd_sc_hd__clkbuf_16
X_1200_ _1808_/CLK _1200_/D VGND VGND VPWR VPWR _1201_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_38_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1131_ _1147_/CLK _1131_/D VGND VGND VPWR VPWR _1132_/D sky130_fd_sc_hd__dfxtp_1
X_1062_ _1071_/CLK _1062_/D VGND VGND VPWR VPWR _1063_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0013_ _1996_/CLK _0013_/D VGND VGND VPWR VPWR _0014_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_clk clkbuf_4_3_0_clk/X VGND VGND VPWR VPWR _1841_/CLK sky130_fd_sc_hd__clkbuf_16
X_1964_ _1973_/CLK _1964_/D VGND VGND VPWR VPWR _1966_/D sky130_fd_sc_hd__dfxtp_1
X_0915_ _0919_/CLK _0915_/D VGND VGND VPWR VPWR _0916_/D sky130_fd_sc_hd__dfxtp_1
X_1895_ _1975_/CLK _1895_/D VGND VGND VPWR VPWR _1896_/D sky130_fd_sc_hd__dfxtp_1
X_0846_ _0864_/CLK _0846_/D VGND VGND VPWR VPWR _0848_/D sky130_fd_sc_hd__dfxtp_1
X_0777_ _0831_/CLK _0777_/D VGND VGND VPWR VPWR _0778_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1329_ _1336_/CLK _1329_/D VGND VGND VPWR VPWR _1330_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0700_ _1112_/CLK _0700_/D VGND VGND VPWR VPWR _0701_/D sky130_fd_sc_hd__dfxtp_1
X_1680_ _1687_/CLK _1680_/D VGND VGND VPWR VPWR _1681_/D sky130_fd_sc_hd__dfxtp_1
X_0631_ _0632_/CLK _0631_/D VGND VGND VPWR VPWR _0632_/D sky130_fd_sc_hd__dfxtp_1
X_0562_ _0610_/CLK _0562_/D VGND VGND VPWR VPWR _0563_/D sky130_fd_sc_hd__dfxtp_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0493_ _0998_/CLK _0493_/D VGND VGND VPWR VPWR _0494_/D sky130_fd_sc_hd__dfxtp_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_2_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _1320_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1114_ _1163_/CLK _1114_/D VGND VGND VPWR VPWR _1115_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_93_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1045_ _1826_/CLK _1045_/D VGND VGND VPWR VPWR _1056_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_80_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1947_ _1975_/CLK _1947_/D VGND VGND VPWR VPWR _1948_/D sky130_fd_sc_hd__dfxtp_1
X_1878_ _1985_/CLK _1878_/D VGND VGND VPWR VPWR _1879_/D sky130_fd_sc_hd__dfxtp_1
X_0829_ _0831_/CLK _0829_/D VGND VGND VPWR VPWR _0830_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_1_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1801_ _1814_/CLK _1801_/D VGND VGND VPWR VPWR _1802_/D sky130_fd_sc_hd__dfxtp_1
X_1732_ _1736_/CLK _1732_/D VGND VGND VPWR VPWR _1733_/D sky130_fd_sc_hd__dfxtp_1
X_1663_ _1665_/CLK _1663_/D VGND VGND VPWR VPWR _1664_/D sky130_fd_sc_hd__dfxtp_1
X_0614_ _0632_/CLK _0614_/D VGND VGND VPWR VPWR _0615_/D sky130_fd_sc_hd__dfxtp_1
X_1594_ _1594_/CLK _1594_/D VGND VGND VPWR VPWR _1595_/D sky130_fd_sc_hd__dfxtp_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0545_ _0573_/CLK _0545_/D VGND VGND VPWR VPWR _0546_/D sky130_fd_sc_hd__dfxtp_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0476_ _0977_/CLK _0476_/D VGND VGND VPWR VPWR _0477_/D sky130_fd_sc_hd__dfxtp_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1028_ _1033_/CLK _1028_/D VGND VGND VPWR VPWR _1029_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0330_ _1907_/CLK _0330_/D VGND VGND VPWR VPWR _0341_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0261_ _0280_/CLK _0261_/D VGND VGND VPWR VPWR _0262_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0192_ _0214_/CLK _0192_/D VGND VGND VPWR VPWR _0193_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_90_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1715_ _1726_/CLK _1715_/D VGND VGND VPWR VPWR _1716_/D sky130_fd_sc_hd__dfxtp_1
X_1646_ _1649_/CLK _1646_/D VGND VGND VPWR VPWR _1647_/D sky130_fd_sc_hd__dfxtp_1
X_1577_ _1578_/CLK _1577_/D VGND VGND VPWR VPWR _1578_/D sky130_fd_sc_hd__dfxtp_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0528_ _1649_/CLK _0528_/D VGND VGND VPWR VPWR _0539_/D sky130_fd_sc_hd__dfxtp_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0459_ _1182_/CLK _0459_/D VGND VGND VPWR VPWR _0460_/D sky130_fd_sc_hd__dfxtp_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1500_ _1604_/CLK _1500_/D VGND VGND VPWR VPWR _1501_/D sky130_fd_sc_hd__dfxtp_1
X_1431_ _1794_/CLK _1431_/D VGND VGND VPWR VPWR _1432_/D sky130_fd_sc_hd__dfxtp_1
X_1362_ _1364_/CLK _1362_/D VGND VGND VPWR VPWR _1363_/D sky130_fd_sc_hd__dfxtp_1
X_1293_ _1336_/CLK _1293_/D VGND VGND VPWR VPWR _1294_/D sky130_fd_sc_hd__dfxtp_1
X_0313_ _1055_/CLK _0313_/D VGND VGND VPWR VPWR _0314_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0244_ _1980_/CLK _0244_/D VGND VGND VPWR VPWR _0245_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0175_ _1178_/CLK _0175_/D VGND VGND VPWR VPWR _0177_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_63_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1629_ _1673_/CLK _1629_/D VGND VGND VPWR VPWR _1630_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_86_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1980_ _1980_/CLK _1980_/D VGND VGND VPWR VPWR _1981_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_60_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0931_ _1077_/CLK _0931_/D VGND VGND VPWR VPWR _0932_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0862_ _0874_/CLK _0862_/D VGND VGND VPWR VPWR _0863_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0793_ _0793_/CLK _0793_/D VGND VGND VPWR VPWR _0794_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1414_ _1747_/CLK _1414_/D VGND VGND VPWR VPWR _1415_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1345_ _1772_/CLK _1345_/D VGND VGND VPWR VPWR _1346_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1276_ _1348_/CLK _1276_/D VGND VGND VPWR VPWR _1277_/D sky130_fd_sc_hd__dfxtp_1
X_0227_ _1996_/CLK _0227_/D VGND VGND VPWR VPWR _0228_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_51_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0158_ _1170_/CLK _0158_/D VGND VGND VPWR VPWR _0159_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0089_ _1229_/CLK _0089_/D VGND VGND VPWR VPWR _0090_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_105_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1130_ _1147_/CLK _1130_/D VGND VGND VPWR VPWR _1131_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_92_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1061_ _1071_/CLK _1061_/D VGND VGND VPWR VPWR _1062_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_46_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0012_ _1996_/CLK _0012_/D VGND VGND VPWR VPWR _0013_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_61_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1963_ _1973_/CLK _1963_/D VGND VGND VPWR VPWR _1964_/D sky130_fd_sc_hd__dfxtp_1
X_0914_ _0919_/CLK _0914_/D VGND VGND VPWR VPWR _0915_/D sky130_fd_sc_hd__dfxtp_1
X_1894_ _1975_/CLK _1894_/D VGND VGND VPWR VPWR _1895_/D sky130_fd_sc_hd__dfxtp_1
X_0845_ _0845_/CLK _0845_/D VGND VGND VPWR VPWR _0846_/D sky130_fd_sc_hd__dfxtp_1
X_0776_ _0831_/CLK _0776_/D VGND VGND VPWR VPWR _0777_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_29_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1328_ _1336_/CLK _1328_/D VGND VGND VPWR VPWR _1329_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1259_ _1302_/CLK _1259_/D VGND VGND VPWR VPWR _1260_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0630_ _0632_/CLK _0630_/D VGND VGND VPWR VPWR _0631_/D sky130_fd_sc_hd__dfxtp_1
X_0561_ _1649_/CLK _0561_/D VGND VGND VPWR VPWR _0572_/D sky130_fd_sc_hd__dfxtp_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0492_ _0508_/CLK _0492_/D VGND VGND VPWR VPWR _0493_/D sky130_fd_sc_hd__dfxtp_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1113_ _1163_/CLK _1113_/D VGND VGND VPWR VPWR _1114_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1044_ _1046_/CLK _1044_/D VGND VGND VPWR VPWR _1046_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_34_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1946_ _1956_/CLK _1946_/D VGND VGND VPWR VPWR _1947_/D sky130_fd_sc_hd__dfxtp_1
X_1877_ _1987_/CLK _1877_/D VGND VGND VPWR VPWR _1888_/D sky130_fd_sc_hd__dfxtp_1
X_0828_ _0831_/CLK _0828_/D VGND VGND VPWR VPWR _0829_/D sky130_fd_sc_hd__dfxtp_1
X_0759_ _1665_/CLK _0759_/D VGND VGND VPWR VPWR _0770_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_88_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1800_ _1833_/CLK _1800_/D VGND VGND VPWR VPWR _1811_/D sky130_fd_sc_hd__dfxtp_1
X_1731_ _1736_/CLK _1731_/D VGND VGND VPWR VPWR _1732_/D sky130_fd_sc_hd__dfxtp_1
X_1662_ _1665_/CLK _1662_/D VGND VGND VPWR VPWR _1663_/D sky130_fd_sc_hd__dfxtp_1
X_0613_ _0632_/CLK _0613_/D VGND VGND VPWR VPWR _0614_/D sky130_fd_sc_hd__dfxtp_1
X_1593_ _1600_/CLK _1593_/D VGND VGND VPWR VPWR _1594_/D sky130_fd_sc_hd__dfxtp_1
X_0544_ _0573_/CLK _0544_/D VGND VGND VPWR VPWR _0545_/D sky130_fd_sc_hd__dfxtp_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0475_ _0998_/CLK _0475_/D VGND VGND VPWR VPWR _0476_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1027_ _1033_/CLK _1027_/D VGND VGND VPWR VPWR _1028_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1929_ _1956_/CLK _1929_/D VGND VGND VPWR VPWR _1930_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_89_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0260_ _1973_/CLK _0260_/D VGND VGND VPWR VPWR _0261_/D sky130_fd_sc_hd__dfxtp_1
X_0191_ _0214_/CLK _0191_/D VGND VGND VPWR VPWR _0192_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_51_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1714_ _1726_/CLK _1714_/D VGND VGND VPWR VPWR _1715_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1645_ _1649_/CLK _1645_/D VGND VGND VPWR VPWR _1646_/D sky130_fd_sc_hd__dfxtp_1
X_1576_ _1592_/CLK _1576_/D VGND VGND VPWR VPWR _1577_/D sky130_fd_sc_hd__dfxtp_1
X_0527_ _1182_/CLK _0527_/D VGND VGND VPWR VPWR _0529_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0458_ _0585_/CLK _0458_/D VGND VGND VPWR VPWR _0459_/D sky130_fd_sc_hd__dfxtp_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0389_ _0932_/CLK _0389_/D VGND VGND VPWR VPWR _0390_/D sky130_fd_sc_hd__dfxtp_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1430_ _1794_/CLK _1430_/D VGND VGND VPWR VPWR _1431_/D sky130_fd_sc_hd__dfxtp_1
X_1361_ _1364_/CLK _1361_/D VGND VGND VPWR VPWR _1362_/D sky130_fd_sc_hd__dfxtp_1
X_0312_ _1046_/CLK _0312_/D VGND VGND VPWR VPWR _0313_/D sky130_fd_sc_hd__dfxtp_1
X_1292_ _1336_/CLK _1292_/D VGND VGND VPWR VPWR _1293_/D sky130_fd_sc_hd__dfxtp_1
X_0243_ _1980_/CLK _0243_/D VGND VGND VPWR VPWR _0244_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0174_ _1180_/CLK _0174_/D VGND VGND VPWR VPWR _0175_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_24_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1628_ _1673_/CLK _1628_/D VGND VGND VPWR VPWR _1629_/D sky130_fd_sc_hd__dfxtp_1
X_1559_ _1907_/CLK _1559_/D VGND VGND VPWR VPWR _1560_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_74_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0930_ _0932_/CLK _0930_/D VGND VGND VPWR VPWR _0931_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_60_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0861_ _0864_/CLK _0861_/D VGND VGND VPWR VPWR _0862_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_9_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0792_ _1827_/CLK _0792_/D VGND VGND VPWR VPWR _0803_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1413_ _1783_/CLK _1413_/D VGND VGND VPWR VPWR _1414_/D sky130_fd_sc_hd__dfxtp_1
X_1344_ _1772_/CLK _1344_/D VGND VGND VPWR VPWR _1345_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1275_ _1348_/CLK _1275_/D VGND VGND VPWR VPWR _1276_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0226_ _1996_/CLK _0226_/D VGND VGND VPWR VPWR _0227_/D sky130_fd_sc_hd__dfxtp_1
X_0157_ _1170_/CLK _0157_/D VGND VGND VPWR VPWR _0158_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0088_ _1635_/CLK _0088_/D VGND VGND VPWR VPWR _0099_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_24_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1060_ _1071_/CLK _1060_/D VGND VGND VPWR VPWR _1061_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_18_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0011_ _1965_/CLK _0011_/D VGND VGND VPWR VPWR _0022_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_46_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1962_ _1973_/CLK _1962_/D VGND VGND VPWR VPWR _1963_/D sky130_fd_sc_hd__dfxtp_1
X_0913_ _1826_/CLK _0913_/D VGND VGND VPWR VPWR _0924_/D sky130_fd_sc_hd__dfxtp_1
X_1893_ _1991_/CLK _1893_/D VGND VGND VPWR VPWR _1894_/D sky130_fd_sc_hd__dfxtp_1
X_0844_ _0864_/CLK _0844_/D VGND VGND VPWR VPWR _0845_/D sky130_fd_sc_hd__dfxtp_1
X_0775_ _0831_/CLK _0775_/D VGND VGND VPWR VPWR _0776_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_96_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1327_ _1336_/CLK _1327_/D VGND VGND VPWR VPWR _1328_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_29_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1258_ _1302_/CLK _1258_/D VGND VGND VPWR VPWR _1259_/D sky130_fd_sc_hd__dfxtp_1
X_0209_ _1594_/CLK _0209_/D VGND VGND VPWR VPWR _0220_/D sky130_fd_sc_hd__dfxtp_1
X_1189_ _1816_/CLK _1189_/D VGND VGND VPWR VPWR _1190_/D sky130_fd_sc_hd__dfxtp_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0560_ _0610_/CLK _0560_/D VGND VGND VPWR VPWR _0562_/D sky130_fd_sc_hd__dfxtp_1
X_0491_ _0998_/CLK _0491_/D VGND VGND VPWR VPWR _0492_/D sky130_fd_sc_hd__dfxtp_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1112_ _1112_/CLK _1112_/D VGND VGND VPWR VPWR _1113_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_93_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1043_ _1046_/CLK _1043_/D VGND VGND VPWR VPWR _1044_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1945_ _1975_/CLK _1945_/D VGND VGND VPWR VPWR _1946_/D sky130_fd_sc_hd__dfxtp_1
X_1876_ _1995_/CLK _1876_/D VGND VGND VPWR VPWR _1878_/D sky130_fd_sc_hd__dfxtp_1
X_0827_ _0831_/CLK _0827_/D VGND VGND VPWR VPWR _0828_/D sky130_fd_sc_hd__dfxtp_1
X_0758_ _0761_/CLK _0758_/D VGND VGND VPWR VPWR _0760_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_103_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0689_ _0898_/CLK _0689_/D VGND VGND VPWR VPWR _0690_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1730_ _1736_/CLK _1730_/D VGND VGND VPWR VPWR _1731_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_7_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1661_ _1665_/CLK _1661_/D VGND VGND VPWR VPWR _1662_/D sky130_fd_sc_hd__dfxtp_1
X_0612_ _0632_/CLK _0612_/D VGND VGND VPWR VPWR _0613_/D sky130_fd_sc_hd__dfxtp_1
X_1592_ _1592_/CLK _1592_/D VGND VGND VPWR VPWR _1593_/D sky130_fd_sc_hd__dfxtp_1
X_0543_ _0573_/CLK _0543_/D VGND VGND VPWR VPWR _0544_/D sky130_fd_sc_hd__dfxtp_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0474_ _0998_/CLK _0474_/D VGND VGND VPWR VPWR _0475_/D sky130_fd_sc_hd__dfxtp_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1026_ _1033_/CLK _1026_/D VGND VGND VPWR VPWR _1027_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1928_ _1956_/CLK _1928_/D VGND VGND VPWR VPWR _1929_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1859_ _1997_/CLK _1859_/D VGND VGND VPWR VPWR _1860_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0190_ _1178_/CLK _0190_/D VGND VGND VPWR VPWR _0191_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_35_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_70_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _0295_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_31_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1713_ _1726_/CLK _1713_/D VGND VGND VPWR VPWR _1714_/D sky130_fd_sc_hd__dfxtp_1
XANTENNA_0 _1181_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1644_ _1649_/CLK _1644_/D VGND VGND VPWR VPWR _1645_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1575_ _1592_/CLK _1575_/D VGND VGND VPWR VPWR _1576_/D sky130_fd_sc_hd__dfxtp_1
X_0526_ _1182_/CLK _0526_/D VGND VGND VPWR VPWR _0527_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0457_ _0585_/CLK _0457_/D VGND VGND VPWR VPWR _0458_/D sky130_fd_sc_hd__dfxtp_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0388_ _1103_/CLK _0388_/D VGND VGND VPWR VPWR _0389_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1009_ _1010_/CLK _1009_/D VGND VGND VPWR VPWR _1010_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_61_clk clkbuf_4_15_0_clk/X VGND VGND VPWR VPWR _0508_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_52_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _0622_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput2 _1181_/D VGND VGND VPWR VPWR out_window[0] sky130_fd_sc_hd__clkbuf_2
X_1360_ _1364_/CLK _1360_/D VGND VGND VPWR VPWR _1361_/D sky130_fd_sc_hd__dfxtp_1
X_0311_ _1046_/CLK _0311_/D VGND VGND VPWR VPWR _0312_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1291_ _1336_/CLK _1291_/D VGND VGND VPWR VPWR _1292_/D sky130_fd_sc_hd__dfxtp_1
X_0242_ _0539_/CLK _0242_/D VGND VGND VPWR VPWR _0253_/D sky130_fd_sc_hd__dfxtp_1
X_0173_ _1180_/CLK _0173_/D VGND VGND VPWR VPWR _0174_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_63_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_43_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _1181_/CLK sky130_fd_sc_hd__clkbuf_16
X_1627_ _1673_/CLK _1627_/D VGND VGND VPWR VPWR _1628_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1558_ _1594_/CLK _1558_/D VGND VGND VPWR VPWR _1559_/D sky130_fd_sc_hd__dfxtp_1
X_0509_ _0529_/CLK _0509_/D VGND VGND VPWR VPWR _0510_/D sky130_fd_sc_hd__dfxtp_1
X_1489_ _1600_/CLK _1489_/D VGND VGND VPWR VPWR _1490_/D sky130_fd_sc_hd__dfxtp_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_34_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _0908_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_22_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_25_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _0793_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0860_ _0864_/CLK _0860_/D VGND VGND VPWR VPWR _0861_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_9_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0791_ _0791_/CLK _0791_/D VGND VGND VPWR VPWR _0793_/D sky130_fd_sc_hd__dfxtp_1
X_1412_ _1747_/CLK _1412_/D VGND VGND VPWR VPWR _1413_/D sky130_fd_sc_hd__dfxtp_1
X_1343_ _1373_/CLK _1343_/D VGND VGND VPWR VPWR _1344_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_3_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1274_ _1302_/CLK _1274_/D VGND VGND VPWR VPWR _1275_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0225_ _1996_/CLK _0225_/D VGND VGND VPWR VPWR _0226_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0156_ _1170_/CLK _0156_/D VGND VGND VPWR VPWR _0157_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0087_ _1229_/CLK _0087_/D VGND VGND VPWR VPWR _0089_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_16_clk clkbuf_4_9_0_clk/X VGND VGND VPWR VPWR _1162_/CLK sky130_fd_sc_hd__clkbuf_16
X_0989_ _0998_/CLK _0989_/D VGND VGND VPWR VPWR _0991_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_3_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0010_ _1997_/CLK _0010_/D VGND VGND VPWR VPWR _0012_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_61_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1961_ _1973_/CLK _1961_/D VGND VGND VPWR VPWR _1962_/D sky130_fd_sc_hd__dfxtp_1
X_0912_ _0916_/CLK _0912_/D VGND VGND VPWR VPWR _0914_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_14_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1892_ _1991_/CLK _1892_/D VGND VGND VPWR VPWR _1893_/D sky130_fd_sc_hd__dfxtp_1
X_0843_ _0864_/CLK _0843_/D VGND VGND VPWR VPWR _0844_/D sky130_fd_sc_hd__dfxtp_1
X_0774_ _0845_/CLK _0774_/D VGND VGND VPWR VPWR _0775_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _1244_/CLK sky130_fd_sc_hd__clkbuf_16
X_1326_ _1788_/CLK _1326_/D VGND VGND VPWR VPWR _1327_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_56_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1257_ _1302_/CLK _1257_/D VGND VGND VPWR VPWR _1258_/D sky130_fd_sc_hd__dfxtp_1
X_1188_ _1816_/CLK _1188_/D VGND VGND VPWR VPWR _1189_/D sky130_fd_sc_hd__dfxtp_1
X_0208_ _0316_/CLK _0208_/D VGND VGND VPWR VPWR _0210_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_24_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0139_ _1162_/CLK _0139_/D VGND VGND VPWR VPWR _0140_/D sky130_fd_sc_hd__dfxtp_1
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0490_ _0998_/CLK _0490_/D VGND VGND VPWR VPWR _0491_/D sky130_fd_sc_hd__dfxtp_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1111_ _1841_/CLK _1111_/D VGND VGND VPWR VPWR _1122_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1042_ _1046_/CLK _1042_/D VGND VGND VPWR VPWR _1043_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1944_ _1975_/CLK _1944_/D VGND VGND VPWR VPWR _1945_/D sky130_fd_sc_hd__dfxtp_1
X_1875_ _1995_/CLK _1875_/D VGND VGND VPWR VPWR _1876_/D sky130_fd_sc_hd__dfxtp_1
X_0826_ _0845_/CLK _0826_/D VGND VGND VPWR VPWR _0827_/D sky130_fd_sc_hd__dfxtp_1
X_0757_ _0761_/CLK _0757_/D VGND VGND VPWR VPWR _0758_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0688_ _0906_/CLK _0688_/D VGND VGND VPWR VPWR _0689_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_15_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_4_15_0_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1309_ _1320_/CLK _1309_/D VGND VGND VPWR VPWR _1310_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1660_ _1665_/CLK _1660_/D VGND VGND VPWR VPWR _1661_/D sky130_fd_sc_hd__dfxtp_1
X_0611_ _0632_/CLK _0611_/D VGND VGND VPWR VPWR _0612_/D sky130_fd_sc_hd__dfxtp_1
X_1591_ _1600_/CLK _1591_/D VGND VGND VPWR VPWR _1592_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_7_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0542_ _0573_/CLK _0542_/D VGND VGND VPWR VPWR _0543_/D sky130_fd_sc_hd__dfxtp_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0473_ _0539_/CLK _0473_/D VGND VGND VPWR VPWR _0484_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1025_ _1033_/CLK _1025_/D VGND VGND VPWR VPWR _1026_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1927_ _1936_/CLK _1927_/D VGND VGND VPWR VPWR _1928_/D sky130_fd_sc_hd__dfxtp_1
X_1858_ _1858_/CLK _1858_/D VGND VGND VPWR VPWR _1859_/D sky130_fd_sc_hd__dfxtp_1
X_0809_ _0813_/CLK _0809_/D VGND VGND VPWR VPWR _0810_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1789_ _1833_/CLK _1789_/D VGND VGND VPWR VPWR _1800_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_1_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1712_ _1726_/CLK _1712_/D VGND VGND VPWR VPWR _1713_/D sky130_fd_sc_hd__dfxtp_1
XANTENNA_1 _1182_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1643_ _1649_/CLK _1643_/D VGND VGND VPWR VPWR _1644_/D sky130_fd_sc_hd__dfxtp_1
X_1574_ _1592_/CLK _1574_/D VGND VGND VPWR VPWR _1575_/D sky130_fd_sc_hd__dfxtp_1
X_0525_ _1182_/CLK _0525_/D VGND VGND VPWR VPWR _0526_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0456_ _0585_/CLK _0456_/D VGND VGND VPWR VPWR _0457_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_86_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0387_ _0908_/CLK _0387_/D VGND VGND VPWR VPWR _0388_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1008_ _1017_/CLK _1008_/D VGND VGND VPWR VPWR _1009_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_1_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput3 _1182_/D VGND VGND VPWR VPWR out_window[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_68_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0310_ _1046_/CLK _0310_/D VGND VGND VPWR VPWR _0311_/D sky130_fd_sc_hd__dfxtp_1
X_1290_ _1336_/CLK _1290_/D VGND VGND VPWR VPWR _1291_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_48_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0241_ _1980_/CLK _0241_/D VGND VGND VPWR VPWR _0243_/D sky130_fd_sc_hd__dfxtp_1
X_0172_ _1178_/CLK _0172_/D VGND VGND VPWR VPWR _0173_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1626_ _1673_/CLK _1626_/D VGND VGND VPWR VPWR _1627_/D sky130_fd_sc_hd__dfxtp_1
X_1557_ _1907_/CLK _1557_/D VGND VGND VPWR VPWR _1558_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0508_ _0508_/CLK _0508_/D VGND VGND VPWR VPWR _0509_/D sky130_fd_sc_hd__dfxtp_1
X_1488_ _1965_/CLK _1488_/D VGND VGND VPWR VPWR _1489_/D sky130_fd_sc_hd__dfxtp_1
X_0439_ _0973_/CLK _0439_/D VGND VGND VPWR VPWR _0441_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_39_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0790_ _0793_/CLK _0790_/D VGND VGND VPWR VPWR _0791_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_42_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1411_ _1710_/CLK _1411_/D VGND VGND VPWR VPWR _1412_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_96_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1342_ _1772_/CLK _1342_/D VGND VGND VPWR VPWR _1343_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_3_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1273_ _1348_/CLK _1273_/D VGND VGND VPWR VPWR _1274_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0224_ _1996_/CLK _0224_/D VGND VGND VPWR VPWR _0225_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0155_ _1170_/CLK _0155_/D VGND VGND VPWR VPWR _0156_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0086_ _1229_/CLK _0086_/D VGND VGND VPWR VPWR _0087_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0988_ _1017_/CLK _0988_/D VGND VGND VPWR VPWR _0989_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_87_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1609_ _1965_/CLK _1609_/D VGND VGND VPWR VPWR _1610_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1960_ _1973_/CLK _1960_/D VGND VGND VPWR VPWR _1961_/D sky130_fd_sc_hd__dfxtp_1
X_0911_ _0919_/CLK _0911_/D VGND VGND VPWR VPWR _0912_/D sky130_fd_sc_hd__dfxtp_1
X_1891_ _1991_/CLK _1891_/D VGND VGND VPWR VPWR _1892_/D sky130_fd_sc_hd__dfxtp_1
X_0842_ _0864_/CLK _0842_/D VGND VGND VPWR VPWR _0843_/D sky130_fd_sc_hd__dfxtp_1
X_0773_ _0845_/CLK _0773_/D VGND VGND VPWR VPWR _0774_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1325_ _1336_/CLK _1325_/D VGND VGND VPWR VPWR _1326_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1256_ _1302_/CLK _1256_/D VGND VGND VPWR VPWR _1257_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1187_ _1841_/CLK _1187_/D VGND VGND VPWR VPWR _1188_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0207_ _0214_/CLK _0207_/D VGND VGND VPWR VPWR _0208_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_24_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0138_ _1162_/CLK _0138_/D VGND VGND VPWR VPWR _0139_/D sky130_fd_sc_hd__dfxtp_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0069_ _1816_/CLK _0069_/D VGND VGND VPWR VPWR _0070_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_3_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1110_ _1163_/CLK _1110_/D VGND VGND VPWR VPWR _1112_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1041_ _1055_/CLK _1041_/D VGND VGND VPWR VPWR _1042_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1943_ _1987_/CLK _1943_/D VGND VGND VPWR VPWR _1954_/D sky130_fd_sc_hd__dfxtp_1
X_1874_ _1995_/CLK _1874_/D VGND VGND VPWR VPWR _1875_/D sky130_fd_sc_hd__dfxtp_1
X_0825_ _1827_/CLK _0825_/D VGND VGND VPWR VPWR _0836_/D sky130_fd_sc_hd__dfxtp_1
X_0756_ _0761_/CLK _0756_/D VGND VGND VPWR VPWR _0757_/D sky130_fd_sc_hd__dfxtp_1
X_0687_ _0898_/CLK _0687_/D VGND VGND VPWR VPWR _0688_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_84_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1308_ _1320_/CLK _1308_/D VGND VGND VPWR VPWR _1309_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_25_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1239_ _1244_/CLK _1239_/D VGND VGND VPWR VPWR _1240_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_25_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0610_ _0610_/CLK _0610_/D VGND VGND VPWR VPWR _0611_/D sky130_fd_sc_hd__dfxtp_1
X_1590_ _1600_/CLK _1590_/D VGND VGND VPWR VPWR _1591_/D sky130_fd_sc_hd__dfxtp_1
X_0541_ _0573_/CLK _0541_/D VGND VGND VPWR VPWR _0542_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0472_ _0998_/CLK _0472_/D VGND VGND VPWR VPWR _0474_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_3_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1024_ _1039_/CLK _1024_/D VGND VGND VPWR VPWR _1025_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_22_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1926_ _1956_/CLK _1926_/D VGND VGND VPWR VPWR _1927_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1857_ _1997_/CLK _1857_/D VGND VGND VPWR VPWR _1858_/D sky130_fd_sc_hd__dfxtp_1
X_0808_ _0906_/CLK _0808_/D VGND VGND VPWR VPWR _0809_/D sky130_fd_sc_hd__dfxtp_1
X_1788_ _1788_/CLK _1788_/D VGND VGND VPWR VPWR _1790_/D sky130_fd_sc_hd__dfxtp_1
X_0739_ _0761_/CLK _0739_/D VGND VGND VPWR VPWR _0740_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_57_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_14_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_4_14_0_clk/X sky130_fd_sc_hd__clkbuf_1
X_1711_ _1726_/CLK _1711_/D VGND VGND VPWR VPWR _1712_/D sky130_fd_sc_hd__dfxtp_1
X_1642_ _1649_/CLK _1642_/D VGND VGND VPWR VPWR _1643_/D sky130_fd_sc_hd__dfxtp_1
X_1573_ _1592_/CLK _1573_/D VGND VGND VPWR VPWR _1574_/D sky130_fd_sc_hd__dfxtp_1
X_0524_ _0529_/CLK _0524_/D VGND VGND VPWR VPWR _0525_/D sky130_fd_sc_hd__dfxtp_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0455_ _0585_/CLK _0455_/D VGND VGND VPWR VPWR _0456_/D sky130_fd_sc_hd__dfxtp_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0386_ _1103_/CLK _0386_/D VGND VGND VPWR VPWR _0387_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_27_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1007_ _1010_/CLK _1007_/D VGND VGND VPWR VPWR _1008_/D sky130_fd_sc_hd__dfxtp_1
X_1909_ _1918_/CLK _1909_/D VGND VGND VPWR VPWR _1911_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_1_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput4 _1183_/D VGND VGND VPWR VPWR out_window[2] sky130_fd_sc_hd__clkbuf_2
X_0240_ _0295_/CLK _0240_/D VGND VGND VPWR VPWR _0241_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0171_ _1180_/CLK _0171_/D VGND VGND VPWR VPWR _0172_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_48_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_120_clk clkbuf_4_0_0_clk/X VGND VGND VPWR VPWR _1373_/CLK sky130_fd_sc_hd__clkbuf_16
X_1625_ _1673_/CLK _1625_/D VGND VGND VPWR VPWR _1626_/D sky130_fd_sc_hd__dfxtp_1
X_1556_ _1592_/CLK _1556_/D VGND VGND VPWR VPWR _1557_/D sky130_fd_sc_hd__dfxtp_1
X_0507_ _0508_/CLK _0507_/D VGND VGND VPWR VPWR _0508_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1487_ _1965_/CLK _1487_/D VGND VGND VPWR VPWR _1488_/D sky130_fd_sc_hd__dfxtp_1
X_0438_ _0973_/CLK _0438_/D VGND VGND VPWR VPWR _0439_/D sky130_fd_sc_hd__dfxtp_1
X_0369_ _1088_/CLK _0369_/D VGND VGND VPWR VPWR _0370_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_94_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_111_clk clkbuf_4_1_0_clk/X VGND VGND VPWR VPWR _1695_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_89_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_102_clk clkbuf_4_6_0_clk/X VGND VGND VPWR VPWR _1659_/CLK sky130_fd_sc_hd__clkbuf_16
X_1410_ _1710_/CLK _1410_/D VGND VGND VPWR VPWR _1411_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_68_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1341_ _1373_/CLK _1341_/D VGND VGND VPWR VPWR _1342_/D sky130_fd_sc_hd__dfxtp_1
X_1272_ _1272_/CLK _1272_/D VGND VGND VPWR VPWR _1273_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0223_ _1996_/CLK _0223_/D VGND VGND VPWR VPWR _0224_/D sky130_fd_sc_hd__dfxtp_1
X_0154_ _1600_/CLK _0154_/D VGND VGND VPWR VPWR _0165_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0085_ _1229_/CLK _0085_/D VGND VGND VPWR VPWR _0086_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0987_ _1017_/CLK _0987_/D VGND VGND VPWR VPWR _0988_/D sky130_fd_sc_hd__dfxtp_1
X_1608_ _1611_/CLK _1608_/D VGND VGND VPWR VPWR _1609_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_87_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1539_ _1578_/CLK _1539_/D VGND VGND VPWR VPWR _1540_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0910_ _0916_/CLK _0910_/D VGND VGND VPWR VPWR _0911_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1890_ _1991_/CLK _1890_/D VGND VGND VPWR VPWR _1891_/D sky130_fd_sc_hd__dfxtp_1
X_0841_ _0864_/CLK _0841_/D VGND VGND VPWR VPWR _0842_/D sky130_fd_sc_hd__dfxtp_1
X_0772_ _0791_/CLK _0772_/D VGND VGND VPWR VPWR _0773_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_102_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1324_ _1788_/CLK _1324_/D VGND VGND VPWR VPWR _1325_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_56_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1255_ _1272_/CLK _1255_/D VGND VGND VPWR VPWR _1256_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_37_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1186_ _1816_/CLK _1186_/D VGND VGND VPWR VPWR _1187_/D sky130_fd_sc_hd__dfxtp_1
X_0206_ _1178_/CLK _0206_/D VGND VGND VPWR VPWR _0207_/D sky130_fd_sc_hd__dfxtp_1
X_0137_ _1185_/CLK _0137_/D VGND VGND VPWR VPWR _0138_/D sky130_fd_sc_hd__dfxtp_1
X_0068_ _1816_/CLK _0068_/D VGND VGND VPWR VPWR _0069_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1040_ _1046_/CLK _1040_/D VGND VGND VPWR VPWR _1041_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1942_ _1975_/CLK _1942_/D VGND VGND VPWR VPWR _1944_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1873_ _1995_/CLK _1873_/D VGND VGND VPWR VPWR _1874_/D sky130_fd_sc_hd__dfxtp_1
X_0824_ _0845_/CLK _0824_/D VGND VGND VPWR VPWR _0826_/D sky130_fd_sc_hd__dfxtp_1
X_0755_ _0761_/CLK _0755_/D VGND VGND VPWR VPWR _0756_/D sky130_fd_sc_hd__dfxtp_1
X_0686_ _0898_/CLK _0686_/D VGND VGND VPWR VPWR _0687_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_103_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1307_ _1320_/CLK _1307_/D VGND VGND VPWR VPWR _1308_/D sky130_fd_sc_hd__dfxtp_1
X_1238_ _1272_/CLK _1238_/D VGND VGND VPWR VPWR _1239_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_91_clk clkbuf_4_5_0_clk/X VGND VGND VPWR VPWR _1587_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1169_ _1180_/CLK _1169_/D VGND VGND VPWR VPWR _1170_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_52_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_82_clk clkbuf_4_7_0_clk/X VGND VGND VPWR VPWR _1991_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0540_ _1182_/CLK _0540_/D VGND VGND VPWR VPWR _0541_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_98_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0471_ _0998_/CLK _0471_/D VGND VGND VPWR VPWR _0472_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_3_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1023_ _1686_/CLK _1023_/D VGND VGND VPWR VPWR _1034_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_53_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_73_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _0316_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1925_ _1936_/CLK _1925_/D VGND VGND VPWR VPWR _1926_/D sky130_fd_sc_hd__dfxtp_1
X_1856_ _1862_/CLK _1856_/D VGND VGND VPWR VPWR _1857_/D sky130_fd_sc_hd__dfxtp_1
X_0807_ _0906_/CLK _0807_/D VGND VGND VPWR VPWR _0808_/D sky130_fd_sc_hd__dfxtp_1
X_1787_ _1794_/CLK _1787_/D VGND VGND VPWR VPWR _1788_/D sky130_fd_sc_hd__dfxtp_1
X_0738_ _1138_/CLK _0738_/D VGND VGND VPWR VPWR _0739_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_103_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0669_ _0874_/CLK _0669_/D VGND VGND VPWR VPWR _0670_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_64_clk clkbuf_4_13_0_clk/X VGND VGND VPWR VPWR _1039_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_55_clk clkbuf_4_14_0_clk/X VGND VGND VPWR VPWR _0595_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1710_ _1710_/CLK _1710_/D VGND VGND VPWR VPWR _1711_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_8_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1641_ _1659_/CLK _1641_/D VGND VGND VPWR VPWR _1642_/D sky130_fd_sc_hd__dfxtp_1
X_1572_ _1592_/CLK _1572_/D VGND VGND VPWR VPWR _1573_/D sky130_fd_sc_hd__dfxtp_1
X_0523_ _0529_/CLK _0523_/D VGND VGND VPWR VPWR _0524_/D sky130_fd_sc_hd__dfxtp_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0454_ _0585_/CLK _0454_/D VGND VGND VPWR VPWR _0455_/D sky130_fd_sc_hd__dfxtp_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0385_ _1918_/CLK _0385_/D VGND VGND VPWR VPWR _0396_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_54_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_46_clk clkbuf_4_12_0_clk/X VGND VGND VPWR VPWR _1070_/CLK sky130_fd_sc_hd__clkbuf_16
X_1006_ _1010_/CLK _1006_/D VGND VGND VPWR VPWR _1007_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_22_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1908_ _1936_/CLK _1908_/D VGND VGND VPWR VPWR _1909_/D sky130_fd_sc_hd__dfxtp_1
X_1839_ _1846_/CLK _1839_/D VGND VGND VPWR VPWR _1840_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk clkbuf_4_11_0_clk/X VGND VGND VPWR VPWR _0642_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput5 _1183_/Q VGND VGND VPWR VPWR out_window[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0170_ _1180_/CLK _0170_/D VGND VGND VPWR VPWR _0171_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_91_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_28_clk clkbuf_4_10_0_clk/X VGND VGND VPWR VPWR _0845_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1624_ _1673_/CLK _1624_/D VGND VGND VPWR VPWR _1625_/D sky130_fd_sc_hd__dfxtp_1
X_1555_ _1918_/CLK _1555_/D VGND VGND VPWR VPWR _1556_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0506_ _0539_/CLK _0506_/D VGND VGND VPWR VPWR _0517_/D sky130_fd_sc_hd__dfxtp_1
X_1486_ _1965_/CLK _1486_/D VGND VGND VPWR VPWR _1487_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_100_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0437_ _0973_/CLK _0437_/D VGND VGND VPWR VPWR _0438_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_86_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0368_ _1112_/CLK _0368_/D VGND VGND VPWR VPWR _0369_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_clk clkbuf_4_8_0_clk/X VGND VGND VPWR VPWR _1147_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0299_ _0316_/CLK _0299_/D VGND VGND VPWR VPWR _0300_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_35_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_13_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_4_13_0_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1340_ _1772_/CLK _1340_/D VGND VGND VPWR VPWR _1341_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_3_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1271_ _1272_/CLK _1271_/D VGND VGND VPWR VPWR _1272_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_49_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0222_ _1996_/CLK _0222_/D VGND VGND VPWR VPWR _0223_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0153_ _1170_/CLK _0153_/D VGND VGND VPWR VPWR _0155_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0084_ _1229_/CLK _0084_/D VGND VGND VPWR VPWR _0085_/D sky130_fd_sc_hd__dfxtp_1
X_0986_ _1039_/CLK _0986_/D VGND VGND VPWR VPWR _0987_/D sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_8_clk clkbuf_4_2_0_clk/X VGND VGND VPWR VPWR _1228_/CLK sky130_fd_sc_hd__clkbuf_16
X_1607_ _1611_/CLK _1607_/D VGND VGND VPWR VPWR _1608_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_99_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1538_ _1592_/CLK _1538_/D VGND VGND VPWR VPWR _1539_/D sky130_fd_sc_hd__dfxtp_1
X_1469_ _1726_/CLK _1469_/D VGND VGND VPWR VPWR _1470_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_86_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0840_ _0864_/CLK _0840_/D VGND VGND VPWR VPWR _0841_/D sky130_fd_sc_hd__dfxtp_1
X_0771_ _0791_/CLK _0771_/D VGND VGND VPWR VPWR _0772_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1323_ _1788_/CLK _1323_/D VGND VGND VPWR VPWR _1324_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1254_ _1302_/CLK _1254_/D VGND VGND VPWR VPWR _1255_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_37_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0205_ _1178_/CLK _0205_/D VGND VGND VPWR VPWR _0206_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_76_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1185_ _1185_/CLK _1185_/D VGND VGND VPWR VPWR _1186_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_37_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0136_ _1147_/CLK _0136_/D VGND VGND VPWR VPWR _0137_/D sky130_fd_sc_hd__dfxtp_1
X_0067_ _1185_/CLK _0067_/D VGND VGND VPWR VPWR _0068_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_20_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0969_ _0973_/CLK _0969_/D VGND VGND VPWR VPWR _0970_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_106_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1941_ _1975_/CLK _1941_/D VGND VGND VPWR VPWR _1942_/D sky130_fd_sc_hd__dfxtp_1
X_1872_ _1995_/CLK _1872_/D VGND VGND VPWR VPWR _1873_/D sky130_fd_sc_hd__dfxtp_1
X_0823_ _0831_/CLK _0823_/D VGND VGND VPWR VPWR _0824_/D sky130_fd_sc_hd__dfxtp_1
X_0754_ _0761_/CLK _0754_/D VGND VGND VPWR VPWR _0755_/D sky130_fd_sc_hd__dfxtp_1
X_0685_ _0898_/CLK _0685_/D VGND VGND VPWR VPWR _0686_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_69_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1306_ _1336_/CLK _1306_/D VGND VGND VPWR VPWR _1307_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1237_ _1272_/CLK _1237_/D VGND VGND VPWR VPWR _1238_/D sky130_fd_sc_hd__dfxtp_1
X_1168_ _1180_/CLK _1168_/D VGND VGND VPWR VPWR _1169_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0119_ _1138_/CLK _0119_/D VGND VGND VPWR VPWR _0120_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1099_ _1104_/CLK _1099_/D VGND VGND VPWR VPWR _1101_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_40_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0470_ _0977_/CLK _0470_/D VGND VGND VPWR VPWR _0471_/D sky130_fd_sc_hd__dfxtp_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1022_ _1033_/CLK _1022_/D VGND VGND VPWR VPWR _1024_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1924_ _1936_/CLK _1924_/D VGND VGND VPWR VPWR _1925_/D sky130_fd_sc_hd__dfxtp_1
X_1855_ _1987_/CLK _1855_/D VGND VGND VPWR VPWR _1866_/D sky130_fd_sc_hd__dfxtp_1
X_0806_ _0813_/CLK _0806_/D VGND VGND VPWR VPWR _0807_/D sky130_fd_sc_hd__dfxtp_1
X_1786_ _1794_/CLK _1786_/D VGND VGND VPWR VPWR _1787_/D sky130_fd_sc_hd__dfxtp_1
X_0737_ _1827_/CLK _0737_/D VGND VGND VPWR VPWR _0748_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_89_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0668_ _0916_/CLK _0668_/D VGND VGND VPWR VPWR _0669_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_39_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0599_ _0632_/CLK _0599_/D VGND VGND VPWR VPWR _0600_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1640_ _1649_/CLK _1640_/D VGND VGND VPWR VPWR _1641_/D sky130_fd_sc_hd__dfxtp_1
X_1571_ _1592_/CLK _1571_/D VGND VGND VPWR VPWR _1572_/D sky130_fd_sc_hd__dfxtp_1
X_0522_ _1182_/CLK _0522_/D VGND VGND VPWR VPWR _0523_/D sky130_fd_sc_hd__dfxtp_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0453_ _0585_/CLK _0453_/D VGND VGND VPWR VPWR _0454_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_79_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0384_ _0908_/CLK _0384_/D VGND VGND VPWR VPWR _0386_/D sky130_fd_sc_hd__dfxtp_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1005_ _1010_/CLK _1005_/D VGND VGND VPWR VPWR _1006_/D sky130_fd_sc_hd__dfxtp_1
X_1907_ _1907_/CLK _1907_/D VGND VGND VPWR VPWR _1908_/D sky130_fd_sc_hd__dfxtp_1
X_1838_ _1846_/CLK _1838_/D VGND VGND VPWR VPWR _1839_/D sky130_fd_sc_hd__dfxtp_1
X_1769_ _1788_/CLK _1769_/D VGND VGND VPWR VPWR _1770_/D sky130_fd_sc_hd__dfxtp_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1623_ _1673_/CLK _1623_/D VGND VGND VPWR VPWR _1624_/D sky130_fd_sc_hd__dfxtp_1
X_1554_ _1907_/CLK _1554_/D VGND VGND VPWR VPWR _1555_/D sky130_fd_sc_hd__dfxtp_1
X_0505_ _0508_/CLK _0505_/D VGND VGND VPWR VPWR _0507_/D sky130_fd_sc_hd__dfxtp_1
X_1485_ _1965_/CLK _1485_/D VGND VGND VPWR VPWR _1486_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0436_ _0966_/CLK _0436_/D VGND VGND VPWR VPWR _0437_/D sky130_fd_sc_hd__dfxtp_1
.ends

