magic
tech sky130A
magscale 1 2
timestamp 1636908413
<< locali >>
rect 39681 60027 39715 60197
rect 14657 56287 14691 56457
rect 59461 49215 59495 54485
rect 59461 32895 59495 34901
rect 59461 24123 59495 28373
rect 59553 24395 59587 29461
rect 59461 6987 59495 9945
<< viali >>
rect 27353 60197 27387 60231
rect 38853 60197 38887 60231
rect 39681 60197 39715 60231
rect 58633 60197 58667 60231
rect 6469 60061 6503 60095
rect 11713 60061 11747 60095
rect 29929 60061 29963 60095
rect 32137 60061 32171 60095
rect 35357 60061 35391 60095
rect 37473 60061 37507 60095
rect 39865 60061 39899 60095
rect 45017 60061 45051 60095
rect 47777 60061 47811 60095
rect 50169 60061 50203 60095
rect 53389 60061 53423 60095
rect 6736 59993 6770 60027
rect 11980 59993 12014 60027
rect 27261 59993 27295 60027
rect 27537 59993 27571 60027
rect 30196 59993 30230 60027
rect 32382 59993 32416 60027
rect 35624 59993 35658 60027
rect 37740 59993 37774 60027
rect 39681 59993 39715 60027
rect 40110 59993 40144 60027
rect 45284 59993 45318 60027
rect 48044 59993 48078 60027
rect 50436 59993 50470 60027
rect 53656 59993 53690 60027
rect 58449 59993 58483 60027
rect 7849 59925 7883 59959
rect 13093 59925 13127 59959
rect 31309 59925 31343 59959
rect 33517 59925 33551 59959
rect 36737 59925 36771 59959
rect 41245 59925 41279 59959
rect 46397 59925 46431 59959
rect 49157 59925 49191 59959
rect 51549 59925 51583 59959
rect 54769 59925 54803 59959
rect 7757 59721 7791 59755
rect 12909 59721 12943 59755
rect 31585 59721 31619 59755
rect 33977 59721 34011 59755
rect 38945 59721 38979 59755
rect 46949 59721 46983 59755
rect 54953 59721 54987 59755
rect 30472 59653 30506 59687
rect 6377 59585 6411 59619
rect 6644 59585 6678 59619
rect 8217 59585 8251 59619
rect 8484 59585 8518 59619
rect 11796 59585 11830 59619
rect 13369 59585 13403 59619
rect 13636 59585 13670 59619
rect 19901 59585 19935 59619
rect 20168 59585 20202 59619
rect 22744 59585 22778 59619
rect 24317 59585 24351 59619
rect 24584 59585 24618 59619
rect 26985 59585 27019 59619
rect 27252 59585 27286 59619
rect 30205 59585 30239 59619
rect 32853 59585 32887 59619
rect 34704 59585 34738 59619
rect 37565 59585 37599 59619
rect 37832 59585 37866 59619
rect 40684 59585 40718 59619
rect 43904 59585 43938 59619
rect 45569 59585 45603 59619
rect 45836 59585 45870 59619
rect 48881 59585 48915 59619
rect 49148 59585 49182 59619
rect 51080 59585 51114 59619
rect 53840 59585 53874 59619
rect 56221 59585 56255 59619
rect 11529 59517 11563 59551
rect 22477 59517 22511 59551
rect 32597 59517 32631 59551
rect 34437 59517 34471 59551
rect 40417 59517 40451 59551
rect 43637 59517 43671 59551
rect 50813 59517 50847 59551
rect 53573 59517 53607 59551
rect 55965 59517 55999 59551
rect 9597 59381 9631 59415
rect 14749 59381 14783 59415
rect 21281 59381 21315 59415
rect 23857 59381 23891 59415
rect 25697 59381 25731 59415
rect 28365 59381 28399 59415
rect 35817 59381 35851 59415
rect 41797 59381 41831 59415
rect 45017 59381 45051 59415
rect 50261 59381 50295 59415
rect 52193 59381 52227 59415
rect 57345 59381 57379 59415
rect 8125 59177 8159 59211
rect 23857 59177 23891 59211
rect 39037 59177 39071 59211
rect 44465 59177 44499 59211
rect 54769 59177 54803 59211
rect 56701 59177 56735 59211
rect 25789 59041 25823 59075
rect 37657 59041 37691 59075
rect 4905 58973 4939 59007
rect 6745 58973 6779 59007
rect 8953 58973 8987 59007
rect 9220 58973 9254 59007
rect 10793 58973 10827 59007
rect 14105 58973 14139 59007
rect 14372 58973 14406 59007
rect 15945 58973 15979 59007
rect 20545 58973 20579 59007
rect 22477 58973 22511 59007
rect 26056 58973 26090 59007
rect 27629 58973 27663 59007
rect 27896 58973 27930 59007
rect 30297 58973 30331 59007
rect 32137 58973 32171 59007
rect 35633 58973 35667 59007
rect 35900 58973 35934 59007
rect 41245 58973 41279 59007
rect 43085 58973 43119 59007
rect 46397 58973 46431 59007
rect 48237 58973 48271 59007
rect 51549 58973 51583 59007
rect 51816 58973 51850 59007
rect 53389 58973 53423 59007
rect 55321 58973 55355 59007
rect 55577 58973 55611 59007
rect 57253 58973 57287 59007
rect 5172 58905 5206 58939
rect 7012 58905 7046 58939
rect 11060 58905 11094 58939
rect 16190 58905 16224 58939
rect 20812 58905 20846 58939
rect 22744 58905 22778 58939
rect 30564 58905 30598 58939
rect 32382 58905 32416 58939
rect 37924 58905 37958 58939
rect 41512 58905 41546 58939
rect 43352 58905 43386 58939
rect 46664 58905 46698 58939
rect 48504 58905 48538 58939
rect 53656 58905 53690 58939
rect 57498 58905 57532 58939
rect 6285 58837 6319 58871
rect 10333 58837 10367 58871
rect 12173 58837 12207 58871
rect 15485 58837 15519 58871
rect 17325 58837 17359 58871
rect 21925 58837 21959 58871
rect 27169 58837 27203 58871
rect 29009 58837 29043 58871
rect 31677 58837 31711 58871
rect 33517 58837 33551 58871
rect 37013 58837 37047 58871
rect 42625 58837 42659 58871
rect 47777 58837 47811 58871
rect 49617 58837 49651 58871
rect 52929 58837 52963 58871
rect 58633 58837 58667 58871
rect 7757 58633 7791 58667
rect 9597 58633 9631 58667
rect 14749 58633 14783 58667
rect 21281 58633 21315 58667
rect 25973 58633 26007 58667
rect 31585 58633 31619 58667
rect 38853 58633 38887 58667
rect 41889 58633 41923 58667
rect 45201 58633 45235 58667
rect 47041 58633 47075 58667
rect 6622 58565 6656 58599
rect 8484 58565 8518 58599
rect 11796 58565 11830 58599
rect 13614 58565 13648 58599
rect 20168 58565 20202 58599
rect 23020 58565 23054 58599
rect 28172 58565 28206 58599
rect 30472 58565 30506 58599
rect 33885 58565 33919 58599
rect 40776 58565 40810 58599
rect 44088 58565 44122 58599
rect 45928 58565 45962 58599
rect 54392 58565 54426 58599
rect 56232 58565 56266 58599
rect 4169 58497 4203 58531
rect 4436 58497 4470 58531
rect 8217 58497 8251 58531
rect 13369 58497 13403 58531
rect 18328 58497 18362 58531
rect 19901 58497 19935 58531
rect 22753 58497 22787 58531
rect 24593 58497 24627 58531
rect 24860 58497 24894 58531
rect 30205 58497 30239 58531
rect 37473 58497 37507 58531
rect 37740 58497 37774 58531
rect 43821 58497 43855 58531
rect 45661 58497 45695 58531
rect 47961 58497 47995 58531
rect 51080 58497 51114 58531
rect 54125 58497 54159 58531
rect 6377 58429 6411 58463
rect 11529 58429 11563 58463
rect 18061 58429 18095 58463
rect 27905 58429 27939 58463
rect 40509 58429 40543 58463
rect 50813 58429 50847 58463
rect 55965 58429 55999 58463
rect 5549 58293 5583 58327
rect 12909 58293 12943 58327
rect 19441 58293 19475 58327
rect 24133 58293 24167 58327
rect 29285 58293 29319 58327
rect 35357 58293 35391 58327
rect 49249 58293 49283 58327
rect 52193 58293 52227 58327
rect 55505 58293 55539 58327
rect 57345 58293 57379 58327
rect 5181 58089 5215 58123
rect 38577 58089 38611 58123
rect 47777 58089 47811 58123
rect 52929 58089 52963 58123
rect 54769 58089 54803 58123
rect 10333 58021 10367 58055
rect 21741 58021 21775 58055
rect 40417 57953 40451 57987
rect 48237 57953 48271 57987
rect 3801 57885 3835 57919
rect 5641 57885 5675 57919
rect 8953 57885 8987 57919
rect 9220 57885 9254 57919
rect 10793 57885 10827 57919
rect 17325 57885 17359 57919
rect 25789 57885 25823 57919
rect 27629 57885 27663 57919
rect 27896 57885 27930 57919
rect 30941 57885 30975 57919
rect 32781 57885 32815 57919
rect 33048 57885 33082 57919
rect 35357 57885 35391 57919
rect 35624 57885 35658 57919
rect 37197 57885 37231 57919
rect 40684 57885 40718 57919
rect 43085 57885 43119 57919
rect 43352 57885 43386 57919
rect 46397 57885 46431 57919
rect 51549 57885 51583 57919
rect 53389 57885 53423 57919
rect 53656 57885 53690 57919
rect 55321 57885 55355 57919
rect 57161 57885 57195 57919
rect 4068 57817 4102 57851
rect 5886 57817 5920 57851
rect 11038 57817 11072 57851
rect 14473 57817 14507 57851
rect 17592 57817 17626 57851
rect 20453 57817 20487 57851
rect 26056 57817 26090 57851
rect 31208 57817 31242 57851
rect 37464 57817 37498 57851
rect 46664 57817 46698 57851
rect 48504 57817 48538 57851
rect 51816 57817 51850 57851
rect 55588 57817 55622 57851
rect 57428 57817 57462 57851
rect 7021 57749 7055 57783
rect 12173 57749 12207 57783
rect 15761 57749 15795 57783
rect 18705 57749 18739 57783
rect 27169 57749 27203 57783
rect 29009 57749 29043 57783
rect 32321 57749 32355 57783
rect 34161 57749 34195 57783
rect 36737 57749 36771 57783
rect 41797 57749 41831 57783
rect 44465 57749 44499 57783
rect 49617 57749 49651 57783
rect 56701 57749 56735 57783
rect 58541 57749 58575 57783
rect 4997 57545 5031 57579
rect 12909 57545 12943 57579
rect 21281 57545 21315 57579
rect 26433 57545 26467 57579
rect 31585 57545 31619 57579
rect 40325 57545 40359 57579
rect 50353 57545 50387 57579
rect 54401 57545 54435 57579
rect 11796 57477 11830 57511
rect 14372 57477 14406 57511
rect 18328 57477 18362 57511
rect 23480 57477 23514 57511
rect 25320 57477 25354 57511
rect 27896 57477 27930 57511
rect 30472 57477 30506 57511
rect 34958 57477 34992 57511
rect 39037 57477 39071 57511
rect 51080 57477 51114 57511
rect 53113 57477 53147 57511
rect 3884 57409 3918 57443
rect 7196 57409 7230 57443
rect 8769 57409 8803 57443
rect 14105 57409 14139 57443
rect 18061 57409 18095 57443
rect 19901 57409 19935 57443
rect 20168 57409 20202 57443
rect 30205 57409 30239 57443
rect 33140 57409 33174 57443
rect 42441 57409 42475 57443
rect 42708 57409 42742 57443
rect 44281 57409 44315 57443
rect 44548 57409 44582 57443
rect 49240 57409 49274 57443
rect 55321 57409 55355 57443
rect 55588 57409 55622 57443
rect 3617 57341 3651 57375
rect 6929 57341 6963 57375
rect 10517 57341 10551 57375
rect 11529 57341 11563 57375
rect 23213 57341 23247 57375
rect 25053 57341 25087 57375
rect 27629 57341 27663 57375
rect 32873 57341 32907 57375
rect 34713 57341 34747 57375
rect 48973 57341 49007 57375
rect 50813 57341 50847 57375
rect 8309 57205 8343 57239
rect 15485 57205 15519 57239
rect 19441 57205 19475 57239
rect 24593 57205 24627 57239
rect 29009 57205 29043 57239
rect 34253 57205 34287 57239
rect 36093 57205 36127 57239
rect 43821 57205 43855 57239
rect 45661 57205 45695 57239
rect 52193 57205 52227 57239
rect 56701 57205 56735 57239
rect 5181 57001 5215 57035
rect 8309 57001 8343 57035
rect 12909 57001 12943 57035
rect 15853 57001 15887 57035
rect 18705 57001 18739 57035
rect 23857 57001 23891 57035
rect 26065 57001 26099 57035
rect 28917 57001 28951 57035
rect 32321 57001 32355 57035
rect 34161 57001 34195 57035
rect 38669 57001 38703 57035
rect 49617 57001 49651 57035
rect 52929 57001 52963 57035
rect 54769 57001 54803 57035
rect 56701 57001 56735 57035
rect 58541 57001 58575 57035
rect 8953 56865 8987 56899
rect 14473 56865 14507 56899
rect 19901 56865 19935 56899
rect 22477 56865 22511 56899
rect 32781 56865 32815 56899
rect 37289 56865 37323 56899
rect 40877 56865 40911 56899
rect 42717 56865 42751 56899
rect 45017 56865 45051 56899
rect 51549 56865 51583 56899
rect 55321 56865 55355 56899
rect 3801 56797 3835 56831
rect 6929 56797 6963 56831
rect 7196 56797 7230 56831
rect 11529 56797 11563 56831
rect 11796 56797 11830 56831
rect 14740 56797 14774 56831
rect 17325 56797 17359 56831
rect 20168 56797 20202 56831
rect 22744 56797 22778 56831
rect 27537 56797 27571 56831
rect 27804 56797 27838 56831
rect 30941 56797 30975 56831
rect 31208 56797 31242 56831
rect 34713 56797 34747 56831
rect 34980 56797 35014 56831
rect 41144 56797 41178 56831
rect 48237 56797 48271 56831
rect 48504 56797 48538 56831
rect 51816 56797 51850 56831
rect 53389 56797 53423 56831
rect 57161 56797 57195 56831
rect 57417 56797 57451 56831
rect 4068 56729 4102 56763
rect 9220 56729 9254 56763
rect 17592 56729 17626 56763
rect 24777 56729 24811 56763
rect 33048 56729 33082 56763
rect 37556 56729 37590 56763
rect 42962 56729 42996 56763
rect 45284 56729 45318 56763
rect 53656 56729 53690 56763
rect 55588 56729 55622 56763
rect 10333 56661 10367 56695
rect 21281 56661 21315 56695
rect 36093 56661 36127 56695
rect 42257 56661 42291 56695
rect 44097 56661 44131 56695
rect 46397 56661 46431 56695
rect 4997 56457 5031 56491
rect 8309 56457 8343 56491
rect 14657 56457 14691 56491
rect 23765 56457 23799 56491
rect 34253 56457 34287 56491
rect 39037 56457 39071 56491
rect 41797 56457 41831 56491
rect 43821 56457 43855 56491
rect 45661 56457 45695 56491
rect 50353 56457 50387 56491
rect 55689 56457 55723 56491
rect 9036 56389 9070 56423
rect 3884 56321 3918 56355
rect 7196 56321 7230 56355
rect 8769 56321 8803 56355
rect 12817 56321 12851 56355
rect 13084 56321 13118 56355
rect 15016 56389 15050 56423
rect 18328 56389 18362 56423
rect 20168 56389 20202 56423
rect 22652 56389 22686 56423
rect 27997 56389 28031 56423
rect 34980 56389 35014 56423
rect 40684 56389 40718 56423
rect 44548 56389 44582 56423
rect 49240 56389 49274 56423
rect 51080 56389 51114 56423
rect 19901 56321 19935 56355
rect 22385 56321 22419 56355
rect 24492 56321 24526 56355
rect 30461 56321 30495 56355
rect 32873 56321 32907 56355
rect 33140 56321 33174 56355
rect 37657 56321 37691 56355
rect 37924 56321 37958 56355
rect 40417 56321 40451 56355
rect 42697 56321 42731 56355
rect 48973 56321 49007 56355
rect 50813 56321 50847 56355
rect 54576 56321 54610 56355
rect 3617 56253 3651 56287
rect 6929 56253 6963 56287
rect 14657 56253 14691 56287
rect 14749 56253 14783 56287
rect 18061 56253 18095 56287
rect 24225 56253 24259 56287
rect 30205 56253 30239 56287
rect 34713 56253 34747 56287
rect 42441 56253 42475 56287
rect 44281 56253 44315 56287
rect 54309 56253 54343 56287
rect 19441 56185 19475 56219
rect 36093 56185 36127 56219
rect 52193 56185 52227 56219
rect 10149 56117 10183 56151
rect 14197 56117 14231 56151
rect 16129 56117 16163 56151
rect 21281 56117 21315 56151
rect 25605 56117 25639 56151
rect 29285 56117 29319 56151
rect 31585 56117 31619 56151
rect 21281 55913 21315 55947
rect 28549 55913 28583 55947
rect 39037 55913 39071 55947
rect 43177 55913 43211 55947
rect 46397 55913 46431 55947
rect 49433 55913 49467 55947
rect 54769 55913 54803 55947
rect 8953 55777 8987 55811
rect 14657 55777 14691 55811
rect 37657 55777 37691 55811
rect 45017 55777 45051 55811
rect 9220 55709 9254 55743
rect 12173 55709 12207 55743
rect 14924 55709 14958 55743
rect 17325 55709 17359 55743
rect 17592 55709 17626 55743
rect 19901 55709 19935 55743
rect 20168 55709 20202 55743
rect 21741 55709 21775 55743
rect 24409 55709 24443 55743
rect 27169 55709 27203 55743
rect 27425 55709 27459 55743
rect 32137 55709 32171 55743
rect 35817 55709 35851 55743
rect 40049 55709 40083 55743
rect 40316 55709 40350 55743
rect 45284 55709 45318 55743
rect 48053 55709 48087 55743
rect 48320 55709 48354 55743
rect 50169 55709 50203 55743
rect 53389 55709 53423 55743
rect 53656 55709 53690 55743
rect 4997 55641 5031 55675
rect 12440 55641 12474 55675
rect 22008 55641 22042 55675
rect 24676 55641 24710 55675
rect 32404 55641 32438 55675
rect 36084 55641 36118 55675
rect 37902 55641 37936 55675
rect 41889 55641 41923 55675
rect 50436 55641 50470 55675
rect 56149 55641 56183 55675
rect 6285 55573 6319 55607
rect 10333 55573 10367 55607
rect 13553 55573 13587 55607
rect 16037 55573 16071 55607
rect 18705 55573 18739 55607
rect 23121 55573 23155 55607
rect 25789 55573 25823 55607
rect 33517 55573 33551 55607
rect 37197 55573 37231 55607
rect 41429 55573 41463 55607
rect 51549 55573 51583 55607
rect 57437 55573 57471 55607
rect 5181 55369 5215 55403
rect 8217 55369 8251 55403
rect 13737 55369 13771 55403
rect 15577 55369 15611 55403
rect 19165 55369 19199 55403
rect 21005 55369 21039 55403
rect 23213 55369 23247 55403
rect 25053 55369 25087 55403
rect 30573 55369 30607 55403
rect 33517 55369 33551 55403
rect 36737 55369 36771 55403
rect 40049 55369 40083 55403
rect 41889 55369 41923 55403
rect 49433 55369 49467 55403
rect 54125 55369 54159 55403
rect 55965 55369 55999 55403
rect 4068 55301 4102 55335
rect 9588 55301 9622 55335
rect 12624 55301 12658 55335
rect 14464 55301 14498 55335
rect 18052 55301 18086 55335
rect 19870 55301 19904 55335
rect 40776 55301 40810 55335
rect 45376 55301 45410 55335
rect 52990 55301 53024 55335
rect 3801 55233 3835 55267
rect 6837 55233 6871 55267
rect 7104 55233 7138 55267
rect 12357 55233 12391 55267
rect 17785 55233 17819 55267
rect 19625 55233 19659 55267
rect 22100 55233 22134 55267
rect 23673 55233 23707 55267
rect 23940 55233 23974 55267
rect 27620 55233 27654 55267
rect 29460 55233 29494 55267
rect 32404 55233 32438 55267
rect 35357 55233 35391 55267
rect 35624 55233 35658 55267
rect 38669 55233 38703 55267
rect 38936 55233 38970 55267
rect 45109 55233 45143 55267
rect 48320 55233 48354 55267
rect 49893 55233 49927 55267
rect 50160 55233 50194 55267
rect 52745 55233 52779 55267
rect 54585 55233 54619 55267
rect 54852 55233 54886 55267
rect 9321 55165 9355 55199
rect 14197 55165 14231 55199
rect 21833 55165 21867 55199
rect 27353 55165 27387 55199
rect 29193 55165 29227 55199
rect 32137 55165 32171 55199
rect 40509 55165 40543 55199
rect 48053 55165 48087 55199
rect 28733 55097 28767 55131
rect 10701 55029 10735 55063
rect 46489 55029 46523 55063
rect 51273 55029 51307 55063
rect 23121 54825 23155 54859
rect 25789 54825 25823 54859
rect 28273 54825 28307 54859
rect 36645 54825 36679 54859
rect 41429 54825 41463 54859
rect 49065 54825 49099 54859
rect 51549 54825 51583 54859
rect 6929 54689 6963 54723
rect 14105 54689 14139 54723
rect 21741 54689 21775 54723
rect 57069 54689 57103 54723
rect 5089 54621 5123 54655
rect 9505 54621 9539 54655
rect 9772 54621 9806 54655
rect 14372 54621 14406 54655
rect 15945 54621 15979 54655
rect 19901 54621 19935 54655
rect 24409 54621 24443 54655
rect 24676 54621 24710 54655
rect 26893 54621 26927 54655
rect 29561 54621 29595 54655
rect 35265 54621 35299 54655
rect 37105 54621 37139 54655
rect 40049 54621 40083 54655
rect 42993 54621 43027 54655
rect 45845 54621 45879 54655
rect 46112 54621 46146 54655
rect 47685 54621 47719 54655
rect 50169 54621 50203 54655
rect 50436 54621 50470 54655
rect 52009 54621 52043 54655
rect 52276 54621 52310 54655
rect 5356 54553 5390 54587
rect 7196 54553 7230 54587
rect 16212 54553 16246 54587
rect 20168 54553 20202 54587
rect 22008 54553 22042 54587
rect 27160 54553 27194 54587
rect 29806 54553 29840 54587
rect 32413 54553 32447 54587
rect 33977 54553 34011 54587
rect 35532 54553 35566 54587
rect 37372 54553 37406 54587
rect 40316 54553 40350 54587
rect 43260 54553 43294 54587
rect 47952 54553 47986 54587
rect 57336 54553 57370 54587
rect 6469 54485 6503 54519
rect 8309 54485 8343 54519
rect 10885 54485 10919 54519
rect 15485 54485 15519 54519
rect 17325 54485 17359 54519
rect 21281 54485 21315 54519
rect 30941 54485 30975 54519
rect 38485 54485 38519 54519
rect 44373 54485 44407 54519
rect 47225 54485 47259 54519
rect 53389 54485 53423 54519
rect 58449 54485 58483 54519
rect 59461 54485 59495 54519
rect 7757 54281 7791 54315
rect 23213 54281 23247 54315
rect 25053 54281 25087 54315
rect 28365 54281 28399 54315
rect 30205 54281 30239 54315
rect 33517 54281 33551 54315
rect 48973 54281 49007 54315
rect 50905 54281 50939 54315
rect 56885 54281 56919 54315
rect 6622 54213 6656 54247
rect 9864 54213 9898 54247
rect 14924 54213 14958 54247
rect 18705 54213 18739 54247
rect 22078 54213 22112 54247
rect 23940 54213 23974 54247
rect 29092 54213 29126 54247
rect 45928 54213 45962 54247
rect 49792 54213 49826 54247
rect 3148 54145 3182 54179
rect 6377 54145 6411 54179
rect 9597 54145 9631 54179
rect 11785 54145 11819 54179
rect 14657 54145 14691 54179
rect 16681 54145 16715 54179
rect 16948 54145 16982 54179
rect 23673 54145 23707 54179
rect 26985 54145 27019 54179
rect 27252 54145 27286 54179
rect 28825 54145 28859 54179
rect 32137 54145 32171 54179
rect 32404 54145 32438 54179
rect 34233 54145 34267 54179
rect 38669 54145 38703 54179
rect 38936 54145 38970 54179
rect 40776 54145 40810 54179
rect 43821 54145 43855 54179
rect 44088 54145 44122 54179
rect 47860 54145 47894 54179
rect 49525 54145 49559 54179
rect 53001 54145 53035 54179
rect 55761 54145 55795 54179
rect 2881 54077 2915 54111
rect 11529 54077 11563 54111
rect 20453 54077 20487 54111
rect 21833 54077 21867 54111
rect 33977 54077 34011 54111
rect 40509 54077 40543 54111
rect 45661 54077 45695 54111
rect 47593 54077 47627 54111
rect 52745 54077 52779 54111
rect 55505 54077 55539 54111
rect 4261 53941 4295 53975
rect 10977 53941 11011 53975
rect 12909 53941 12943 53975
rect 16037 53941 16071 53975
rect 18061 53941 18095 53975
rect 35357 53941 35391 53975
rect 40049 53941 40083 53975
rect 41889 53941 41923 53975
rect 45201 53941 45235 53975
rect 47041 53941 47075 53975
rect 54125 53941 54159 53975
rect 11253 53737 11287 53771
rect 15945 53737 15979 53771
rect 17785 53737 17819 53771
rect 22477 53737 22511 53771
rect 27353 53737 27387 53771
rect 32781 53737 32815 53771
rect 39313 53737 39347 53771
rect 42625 53737 42659 53771
rect 52469 53737 52503 53771
rect 3801 53601 3835 53635
rect 5641 53601 5675 53635
rect 14565 53601 14599 53635
rect 43085 53601 43119 53635
rect 51089 53601 51123 53635
rect 4068 53533 4102 53567
rect 9873 53533 9907 53567
rect 10140 53533 10174 53567
rect 11713 53533 11747 53567
rect 11980 53533 12014 53567
rect 14832 53533 14866 53567
rect 16405 53533 16439 53567
rect 16672 53533 16706 53567
rect 19257 53533 19291 53567
rect 21097 53533 21131 53567
rect 25973 53533 26007 53567
rect 29561 53533 29595 53567
rect 29828 53533 29862 53567
rect 31401 53533 31435 53567
rect 34713 53533 34747 53567
rect 37933 53533 37967 53567
rect 38200 53533 38234 53567
rect 41245 53533 41279 53567
rect 45293 53533 45327 53567
rect 45560 53533 45594 53567
rect 47133 53533 47167 53567
rect 51356 53533 51390 53567
rect 52929 53533 52963 53567
rect 53196 53533 53230 53567
rect 56793 53533 56827 53567
rect 5886 53465 5920 53499
rect 19524 53465 19558 53499
rect 21342 53465 21376 53499
rect 26240 53465 26274 53499
rect 31646 53465 31680 53499
rect 34958 53465 34992 53499
rect 41512 53465 41546 53499
rect 43352 53465 43386 53499
rect 57060 53465 57094 53499
rect 5181 53397 5215 53431
rect 7021 53397 7055 53431
rect 13093 53397 13127 53431
rect 20637 53397 20671 53431
rect 30941 53397 30975 53431
rect 36093 53397 36127 53431
rect 44465 53397 44499 53431
rect 46673 53397 46707 53431
rect 48421 53397 48455 53431
rect 54309 53397 54343 53431
rect 58173 53397 58207 53431
rect 3525 53193 3559 53227
rect 5365 53193 5399 53227
rect 7941 53193 7975 53227
rect 19901 53193 19935 53227
rect 26433 53193 26467 53227
rect 30849 53193 30883 53227
rect 33517 53193 33551 53227
rect 40049 53193 40083 53227
rect 41889 53193 41923 53227
rect 44833 53193 44867 53227
rect 48973 53193 49007 53227
rect 55045 53193 55079 53227
rect 57345 53193 57379 53227
rect 4230 53125 4264 53159
rect 6828 53125 6862 53159
rect 13093 53125 13127 53159
rect 14657 53125 14691 53159
rect 16948 53125 16982 53159
rect 23480 53125 23514 53159
rect 29736 53125 29770 53159
rect 32404 53125 32438 53159
rect 34244 53125 34278 53159
rect 38936 53125 38970 53159
rect 40776 53125 40810 53159
rect 45560 53125 45594 53159
rect 56232 53125 56266 53159
rect 2145 53057 2179 53091
rect 2412 53057 2446 53091
rect 3985 53057 4019 53091
rect 6561 53057 6595 53091
rect 16681 53057 16715 53091
rect 18521 53057 18555 53091
rect 18777 53057 18811 53091
rect 23213 53057 23247 53091
rect 25053 53057 25087 53091
rect 25320 53057 25354 53091
rect 29469 53057 29503 53091
rect 32137 53057 32171 53091
rect 33977 53057 34011 53091
rect 38669 53057 38703 53091
rect 40509 53057 40543 53091
rect 43720 53057 43754 53091
rect 47860 53057 47894 53091
rect 53665 53057 53699 53091
rect 53932 53057 53966 53091
rect 55965 53057 55999 53091
rect 43453 52989 43487 53023
rect 45293 52989 45327 53023
rect 47593 52989 47627 53023
rect 46673 52921 46707 52955
rect 18061 52853 18095 52887
rect 24593 52853 24627 52887
rect 35357 52853 35391 52887
rect 3249 52649 3283 52683
rect 5825 52649 5859 52683
rect 18521 52649 18555 52683
rect 26249 52649 26283 52683
rect 34069 52649 34103 52683
rect 41797 52649 41831 52683
rect 44465 52649 44499 52683
rect 48329 52649 48363 52683
rect 54769 52649 54803 52683
rect 57713 52649 57747 52683
rect 10517 52581 10551 52615
rect 23213 52581 23247 52615
rect 9137 52513 9171 52547
rect 24869 52513 24903 52547
rect 43085 52513 43119 52547
rect 56333 52513 56367 52547
rect 1869 52445 1903 52479
rect 2136 52445 2170 52479
rect 4445 52445 4479 52479
rect 4712 52445 4746 52479
rect 9404 52445 9438 52479
rect 11529 52445 11563 52479
rect 11796 52445 11830 52479
rect 14105 52445 14139 52479
rect 17141 52445 17175 52479
rect 17408 52445 17442 52479
rect 19993 52445 20027 52479
rect 20260 52445 20294 52479
rect 21833 52445 21867 52479
rect 22100 52445 22134 52479
rect 25136 52445 25170 52479
rect 26709 52445 26743 52479
rect 26965 52445 26999 52479
rect 32689 52445 32723 52479
rect 32956 52445 32990 52479
rect 40417 52445 40451 52479
rect 40684 52445 40718 52479
rect 43352 52445 43386 52479
rect 46949 52445 46983 52479
rect 47216 52445 47250 52479
rect 51089 52445 51123 52479
rect 51356 52445 51390 52479
rect 53389 52445 53423 52479
rect 53656 52445 53690 52479
rect 14350 52377 14384 52411
rect 56600 52377 56634 52411
rect 12909 52309 12943 52343
rect 15485 52309 15519 52343
rect 21373 52309 21407 52343
rect 28089 52309 28123 52343
rect 52469 52309 52503 52343
rect 3433 52105 3467 52139
rect 10977 52105 11011 52139
rect 13369 52105 13403 52139
rect 20637 52105 20671 52139
rect 40325 52105 40359 52139
rect 44557 52105 44591 52139
rect 46857 52105 46891 52139
rect 48973 52105 49007 52139
rect 54493 52105 54527 52139
rect 57345 52105 57379 52139
rect 11796 52037 11830 52071
rect 19524 52037 19558 52071
rect 27252 52037 27286 52071
rect 33416 52037 33450 52071
rect 43444 52037 43478 52071
rect 51080 52037 51114 52071
rect 2320 51969 2354 52003
rect 6561 51969 6595 52003
rect 6828 51969 6862 52003
rect 9597 51969 9631 52003
rect 9864 51969 9898 52003
rect 11529 51969 11563 52003
rect 13553 51969 13587 52003
rect 14361 51969 14395 52003
rect 16681 51969 16715 52003
rect 16948 51969 16982 52003
rect 22100 51969 22134 52003
rect 23940 51969 23974 52003
rect 28825 51969 28859 52003
rect 29092 51969 29126 52003
rect 33149 51969 33183 52003
rect 35173 51969 35207 52003
rect 35440 51969 35474 52003
rect 38016 51969 38050 52003
rect 40509 51969 40543 52003
rect 47041 51969 47075 52003
rect 47860 51969 47894 52003
rect 53113 51969 53147 52003
rect 53380 51969 53414 52003
rect 55965 51969 55999 52003
rect 56232 51969 56266 52003
rect 2053 51901 2087 51935
rect 14105 51901 14139 51935
rect 19257 51901 19291 51935
rect 21833 51901 21867 51935
rect 23673 51901 23707 51935
rect 26985 51901 27019 51935
rect 37749 51901 37783 51935
rect 43177 51901 43211 51935
rect 47593 51901 47627 51935
rect 50813 51901 50847 51935
rect 12909 51833 12943 51867
rect 7941 51765 7975 51799
rect 15485 51765 15519 51799
rect 18061 51765 18095 51799
rect 23213 51765 23247 51799
rect 25053 51765 25087 51799
rect 28365 51765 28399 51799
rect 30205 51765 30239 51799
rect 34529 51765 34563 51799
rect 36553 51765 36587 51799
rect 39129 51765 39163 51799
rect 52193 51765 52227 51799
rect 3249 51561 3283 51595
rect 8401 51561 8435 51595
rect 13461 51561 13495 51595
rect 49065 51561 49099 51595
rect 54309 51561 54343 51595
rect 57161 51561 57195 51595
rect 19993 51493 20027 51527
rect 14105 51425 14139 51459
rect 24409 51425 24443 51459
rect 39865 51425 39899 51459
rect 45845 51425 45879 51459
rect 1869 51357 1903 51391
rect 5181 51357 5215 51391
rect 7021 51357 7055 51391
rect 10241 51357 10275 51391
rect 12081 51357 12115 51391
rect 14372 51357 14406 51391
rect 15945 51357 15979 51391
rect 20177 51357 20211 51391
rect 20729 51357 20763 51391
rect 27261 51357 27295 51391
rect 29561 51357 29595 51391
rect 32781 51357 32815 51391
rect 33048 51357 33082 51391
rect 34713 51357 34747 51391
rect 36553 51357 36587 51391
rect 47685 51357 47719 51391
rect 50905 51357 50939 51391
rect 51172 51357 51206 51391
rect 52929 51357 52963 51391
rect 53196 51357 53230 51391
rect 2136 51289 2170 51323
rect 5448 51289 5482 51323
rect 7288 51289 7322 51323
rect 10508 51289 10542 51323
rect 12348 51289 12382 51323
rect 16190 51289 16224 51323
rect 20996 51289 21030 51323
rect 24676 51289 24710 51323
rect 29828 51289 29862 51323
rect 34958 51289 34992 51323
rect 36820 51289 36854 51323
rect 40132 51289 40166 51323
rect 46112 51289 46146 51323
rect 47952 51289 47986 51323
rect 55873 51289 55907 51323
rect 6561 51221 6595 51255
rect 11621 51221 11655 51255
rect 15485 51221 15519 51255
rect 17325 51221 17359 51255
rect 22109 51221 22143 51255
rect 25789 51221 25823 51255
rect 28733 51221 28767 51255
rect 30941 51221 30975 51255
rect 34161 51221 34195 51255
rect 36093 51221 36127 51255
rect 37933 51221 37967 51255
rect 41245 51221 41279 51255
rect 47225 51221 47259 51255
rect 52285 51221 52319 51255
rect 3433 51017 3467 51051
rect 9137 51017 9171 51051
rect 10977 51017 11011 51051
rect 13093 51017 13127 51051
rect 18061 51017 18095 51051
rect 21281 51017 21315 51051
rect 23213 51017 23247 51051
rect 25053 51017 25087 51051
rect 34621 51017 34655 51051
rect 40509 51017 40543 51051
rect 48973 51017 49007 51051
rect 57161 51017 57195 51051
rect 4712 50949 4746 50983
rect 9864 50949 9898 50983
rect 14372 50949 14406 50983
rect 22100 50949 22134 50983
rect 23940 50949 23974 50983
rect 27252 50949 27286 50983
rect 33508 50949 33542 50983
rect 35348 50949 35382 50983
rect 37556 50949 37590 50983
rect 47838 50949 47872 50983
rect 51080 50949 51114 50983
rect 2320 50881 2354 50915
rect 4445 50881 4479 50915
rect 8024 50881 8058 50915
rect 11969 50881 12003 50915
rect 16948 50881 16982 50915
rect 20168 50881 20202 50915
rect 23673 50881 23707 50915
rect 29081 50881 29115 50915
rect 33241 50881 33275 50915
rect 35081 50881 35115 50915
rect 37289 50881 37323 50915
rect 39385 50881 39419 50915
rect 42708 50881 42742 50915
rect 44281 50881 44315 50915
rect 44548 50881 44582 50915
rect 55781 50881 55815 50915
rect 56048 50881 56082 50915
rect 2053 50813 2087 50847
rect 7757 50813 7791 50847
rect 9597 50813 9631 50847
rect 11713 50813 11747 50847
rect 14105 50813 14139 50847
rect 16681 50813 16715 50847
rect 19901 50813 19935 50847
rect 21833 50813 21867 50847
rect 26985 50813 27019 50847
rect 28825 50813 28859 50847
rect 39129 50813 39163 50847
rect 42441 50813 42475 50847
rect 47593 50813 47627 50847
rect 50813 50813 50847 50847
rect 5825 50677 5859 50711
rect 15485 50677 15519 50711
rect 28365 50677 28399 50711
rect 30205 50677 30239 50711
rect 36461 50677 36495 50711
rect 38669 50677 38703 50711
rect 43821 50677 43855 50711
rect 45661 50677 45695 50711
rect 52193 50677 52227 50711
rect 3249 50473 3283 50507
rect 5457 50473 5491 50507
rect 7757 50473 7791 50507
rect 11253 50473 11287 50507
rect 15577 50473 15611 50507
rect 17417 50473 17451 50507
rect 23121 50473 23155 50507
rect 25789 50473 25823 50507
rect 30941 50473 30975 50507
rect 37933 50473 37967 50507
rect 48237 50473 48271 50507
rect 57437 50473 57471 50507
rect 6377 50337 6411 50371
rect 14197 50337 14231 50371
rect 16037 50337 16071 50371
rect 19901 50337 19935 50371
rect 21741 50337 21775 50371
rect 36553 50337 36587 50371
rect 39865 50337 39899 50371
rect 56057 50337 56091 50371
rect 1869 50269 1903 50303
rect 4169 50269 4203 50303
rect 6644 50269 6678 50303
rect 9873 50269 9907 50303
rect 12173 50269 12207 50303
rect 14464 50269 14498 50303
rect 16304 50269 16338 50303
rect 24409 50269 24443 50303
rect 24676 50269 24710 50303
rect 26985 50269 27019 50303
rect 27252 50269 27286 50303
rect 29561 50269 29595 50303
rect 29828 50269 29862 50303
rect 31401 50269 31435 50303
rect 34713 50269 34747 50303
rect 34980 50269 35014 50303
rect 36809 50269 36843 50303
rect 40132 50269 40166 50303
rect 41705 50269 41739 50303
rect 41961 50269 41995 50303
rect 45017 50269 45051 50303
rect 46857 50269 46891 50303
rect 50721 50269 50755 50303
rect 50988 50269 51022 50303
rect 2136 50201 2170 50235
rect 10140 50201 10174 50235
rect 12440 50201 12474 50235
rect 20168 50201 20202 50235
rect 21986 50201 22020 50235
rect 31646 50201 31680 50235
rect 45284 50201 45318 50235
rect 47102 50201 47136 50235
rect 56324 50201 56358 50235
rect 13553 50133 13587 50167
rect 21281 50133 21315 50167
rect 28365 50133 28399 50167
rect 32781 50133 32815 50167
rect 36093 50133 36127 50167
rect 41245 50133 41279 50167
rect 43085 50133 43119 50167
rect 46397 50133 46431 50167
rect 52101 50133 52135 50167
rect 16129 49929 16163 49963
rect 21097 49929 21131 49963
rect 24501 49929 24535 49963
rect 26341 49929 26375 49963
rect 30205 49929 30239 49963
rect 33793 49929 33827 49963
rect 44465 49929 44499 49963
rect 52009 49929 52043 49963
rect 54493 49929 54527 49963
rect 6622 49861 6656 49895
rect 13176 49861 13210 49895
rect 18797 49861 18831 49895
rect 23388 49861 23422 49895
rect 27252 49861 27286 49895
rect 29092 49861 29126 49895
rect 32505 49861 32539 49895
rect 34980 49861 35014 49895
rect 37556 49861 37590 49895
rect 39396 49861 39430 49895
rect 43177 49861 43211 49895
rect 45630 49861 45664 49895
rect 49056 49861 49090 49895
rect 50896 49861 50930 49895
rect 1860 49793 1894 49827
rect 4712 49793 4746 49827
rect 9312 49793 9346 49827
rect 12909 49793 12943 49827
rect 15005 49793 15039 49827
rect 17049 49793 17083 49827
rect 19717 49793 19751 49827
rect 19984 49793 20018 49827
rect 24961 49793 24995 49827
rect 25228 49793 25262 49827
rect 26985 49793 27019 49827
rect 28825 49793 28859 49827
rect 34713 49793 34747 49827
rect 37289 49793 37323 49827
rect 39129 49793 39163 49827
rect 48789 49793 48823 49827
rect 53380 49793 53414 49827
rect 54953 49793 54987 49827
rect 55220 49793 55254 49827
rect 1593 49725 1627 49759
rect 4445 49725 4479 49759
rect 6377 49725 6411 49759
rect 9045 49725 9079 49759
rect 14749 49725 14783 49759
rect 23121 49725 23155 49759
rect 45385 49725 45419 49759
rect 50629 49725 50663 49759
rect 53113 49725 53147 49759
rect 28365 49657 28399 49691
rect 36093 49657 36127 49691
rect 38669 49657 38703 49691
rect 2973 49589 3007 49623
rect 5825 49589 5859 49623
rect 7757 49589 7791 49623
rect 10425 49589 10459 49623
rect 14289 49589 14323 49623
rect 40509 49589 40543 49623
rect 46765 49589 46799 49623
rect 50169 49589 50203 49623
rect 56333 49589 56367 49623
rect 2973 49385 3007 49419
rect 6837 49385 6871 49419
rect 13553 49385 13587 49419
rect 21097 49385 21131 49419
rect 26433 49385 26467 49419
rect 31309 49385 31343 49419
rect 36829 49385 36863 49419
rect 41245 49385 41279 49419
rect 46397 49385 46431 49419
rect 58541 49385 58575 49419
rect 5457 49249 5491 49283
rect 14105 49249 14139 49283
rect 17233 49249 17267 49283
rect 19717 49249 19751 49283
rect 22477 49249 22511 49283
rect 25053 49249 25087 49283
rect 29929 49249 29963 49283
rect 39865 49249 39899 49283
rect 48237 49249 48271 49283
rect 55321 49249 55355 49283
rect 57161 49249 57195 49283
rect 1593 49181 1627 49215
rect 1860 49181 1894 49215
rect 5724 49181 5758 49215
rect 8953 49181 8987 49215
rect 12173 49181 12207 49215
rect 14372 49181 14406 49215
rect 17500 49181 17534 49215
rect 31769 49181 31803 49215
rect 32036 49181 32070 49215
rect 35541 49181 35575 49215
rect 40132 49181 40166 49215
rect 41705 49181 41739 49215
rect 45017 49181 45051 49215
rect 45284 49181 45318 49215
rect 48504 49181 48538 49215
rect 50169 49181 50203 49215
rect 52745 49181 52779 49215
rect 55588 49181 55622 49215
rect 57428 49181 57462 49215
rect 59461 49181 59495 49215
rect 9220 49113 9254 49147
rect 12440 49113 12474 49147
rect 19984 49113 20018 49147
rect 22744 49113 22778 49147
rect 25320 49113 25354 49147
rect 30196 49113 30230 49147
rect 41950 49113 41984 49147
rect 50414 49113 50448 49147
rect 53012 49113 53046 49147
rect 10333 49045 10367 49079
rect 15485 49045 15519 49079
rect 18613 49045 18647 49079
rect 23857 49045 23891 49079
rect 33149 49045 33183 49079
rect 43085 49045 43119 49079
rect 49617 49045 49651 49079
rect 51549 49045 51583 49079
rect 54125 49045 54159 49079
rect 56701 49045 56735 49079
rect 3525 48841 3559 48875
rect 5365 48841 5399 48875
rect 10425 48841 10459 48875
rect 21005 48841 21039 48875
rect 26433 48841 26467 48875
rect 41797 48841 41831 48875
rect 46397 48841 46431 48875
rect 56793 48841 56827 48875
rect 2412 48773 2446 48807
rect 4252 48773 4286 48807
rect 9312 48773 9346 48807
rect 17224 48773 17258 48807
rect 32404 48773 32438 48807
rect 40684 48773 40718 48807
rect 43422 48773 43456 48807
rect 49056 48773 49090 48807
rect 55658 48773 55692 48807
rect 2145 48705 2179 48739
rect 6837 48705 6871 48739
rect 8585 48705 8619 48739
rect 9045 48705 9079 48739
rect 11713 48705 11747 48739
rect 11980 48705 12014 48739
rect 13553 48705 13587 48739
rect 13820 48705 13854 48739
rect 16957 48705 16991 48739
rect 19625 48705 19659 48739
rect 19892 48705 19926 48739
rect 22477 48705 22511 48739
rect 22744 48705 22778 48739
rect 25053 48705 25087 48739
rect 25320 48705 25354 48739
rect 30472 48705 30506 48739
rect 33977 48705 34011 48739
rect 34244 48705 34278 48739
rect 37289 48705 37323 48739
rect 37556 48705 37590 48739
rect 43177 48705 43211 48739
rect 45273 48705 45307 48739
rect 48789 48705 48823 48739
rect 53205 48705 53239 48739
rect 3985 48637 4019 48671
rect 30205 48637 30239 48671
rect 32137 48637 32171 48671
rect 40417 48637 40451 48671
rect 45017 48637 45051 48671
rect 55413 48637 55447 48671
rect 50169 48569 50203 48603
rect 13093 48501 13127 48535
rect 14933 48501 14967 48535
rect 18337 48501 18371 48535
rect 23857 48501 23891 48535
rect 31585 48501 31619 48535
rect 33517 48501 33551 48535
rect 35357 48501 35391 48535
rect 38669 48501 38703 48535
rect 44557 48501 44591 48535
rect 54493 48501 54527 48535
rect 22569 48297 22603 48331
rect 53389 48297 53423 48331
rect 10793 48229 10827 48263
rect 12909 48229 12943 48263
rect 16037 48229 16071 48263
rect 20821 48229 20855 48263
rect 26985 48229 27019 48263
rect 33609 48229 33643 48263
rect 43821 48229 43855 48263
rect 56701 48229 56735 48263
rect 4997 48161 5031 48195
rect 17049 48161 17083 48195
rect 19441 48161 19475 48195
rect 36553 48161 36587 48195
rect 42441 48161 42475 48195
rect 45109 48161 45143 48195
rect 48237 48161 48271 48195
rect 50169 48161 50203 48195
rect 9413 48093 9447 48127
rect 9680 48093 9714 48127
rect 11529 48093 11563 48127
rect 14657 48093 14691 48127
rect 14924 48093 14958 48127
rect 17316 48093 17350 48127
rect 21281 48093 21315 48127
rect 25697 48093 25731 48127
rect 30389 48093 30423 48127
rect 30656 48093 30690 48127
rect 32229 48093 32263 48127
rect 32496 48093 32530 48127
rect 34713 48093 34747 48127
rect 39865 48093 39899 48127
rect 42708 48093 42742 48127
rect 48504 48093 48538 48127
rect 52009 48093 52043 48127
rect 55321 48093 55355 48127
rect 55588 48093 55622 48127
rect 5264 48025 5298 48059
rect 11796 48025 11830 48059
rect 19708 48025 19742 48059
rect 34980 48025 35014 48059
rect 36798 48025 36832 48059
rect 40132 48025 40166 48059
rect 45376 48025 45410 48059
rect 50414 48025 50448 48059
rect 52276 48025 52310 48059
rect 6377 47957 6411 47991
rect 18429 47957 18463 47991
rect 31769 47957 31803 47991
rect 36093 47957 36127 47991
rect 37933 47957 37967 47991
rect 41245 47957 41279 47991
rect 46489 47957 46523 47991
rect 49617 47957 49651 47991
rect 51549 47957 51583 47991
rect 15485 47753 15519 47787
rect 20913 47753 20947 47787
rect 24409 47753 24443 47787
rect 26433 47753 26467 47787
rect 35633 47753 35667 47787
rect 44465 47753 44499 47787
rect 50077 47753 50111 47787
rect 54125 47753 54159 47787
rect 11897 47685 11931 47719
rect 17224 47685 17258 47719
rect 23296 47685 23330 47719
rect 28908 47685 28942 47719
rect 32658 47685 32692 47719
rect 39681 47685 39715 47719
rect 43352 47685 43386 47719
rect 48789 47685 48823 47719
rect 3525 47617 3559 47651
rect 3792 47617 3826 47651
rect 6644 47617 6678 47651
rect 14361 47617 14395 47651
rect 16957 47617 16991 47651
rect 19533 47617 19567 47651
rect 19800 47617 19834 47651
rect 23029 47617 23063 47651
rect 25053 47617 25087 47651
rect 25320 47617 25354 47651
rect 32413 47617 32447 47651
rect 34253 47617 34287 47651
rect 34520 47617 34554 47651
rect 37289 47617 37323 47651
rect 37545 47617 37579 47651
rect 43085 47617 43119 47651
rect 44925 47617 44959 47651
rect 45192 47617 45226 47651
rect 53001 47617 53035 47651
rect 6377 47549 6411 47583
rect 13645 47549 13679 47583
rect 14105 47549 14139 47583
rect 28641 47549 28675 47583
rect 41337 47549 41371 47583
rect 52745 47549 52779 47583
rect 4905 47413 4939 47447
rect 7757 47413 7791 47447
rect 18337 47413 18371 47447
rect 30021 47413 30055 47447
rect 33793 47413 33827 47447
rect 38669 47413 38703 47447
rect 46305 47413 46339 47447
rect 5181 47209 5215 47243
rect 7021 47209 7055 47243
rect 20913 47209 20947 47243
rect 26801 47209 26835 47243
rect 36093 47209 36127 47243
rect 46397 47209 46431 47243
rect 49617 47209 49651 47243
rect 53941 47209 53975 47243
rect 29009 47141 29043 47175
rect 5641 47073 5675 47107
rect 19533 47073 19567 47107
rect 22477 47073 22511 47107
rect 25421 47073 25455 47107
rect 27629 47073 27663 47107
rect 48237 47073 48271 47107
rect 3801 47005 3835 47039
rect 5897 47005 5931 47039
rect 10609 47005 10643 47039
rect 14841 47005 14875 47039
rect 16865 47005 16899 47039
rect 17132 47005 17166 47039
rect 22744 47005 22778 47039
rect 27896 47005 27930 47039
rect 31125 47005 31159 47039
rect 31392 47005 31426 47039
rect 34713 47005 34747 47039
rect 36553 47005 36587 47039
rect 36820 47005 36854 47039
rect 39865 47005 39899 47039
rect 41705 47005 41739 47039
rect 41961 47005 41995 47039
rect 45017 47005 45051 47039
rect 48504 47005 48538 47039
rect 50629 47005 50663 47039
rect 50896 47005 50930 47039
rect 52561 47005 52595 47039
rect 52828 47005 52862 47039
rect 4068 46937 4102 46971
rect 10876 46937 10910 46971
rect 15108 46937 15142 46971
rect 19800 46937 19834 46971
rect 25688 46937 25722 46971
rect 34980 46937 35014 46971
rect 40132 46937 40166 46971
rect 45284 46937 45318 46971
rect 11989 46869 12023 46903
rect 16221 46869 16255 46903
rect 18245 46869 18279 46903
rect 23857 46869 23891 46903
rect 32505 46869 32539 46903
rect 37933 46869 37967 46903
rect 41245 46869 41279 46903
rect 43085 46869 43119 46903
rect 52009 46869 52043 46903
rect 3801 46665 3835 46699
rect 5641 46665 5675 46699
rect 7757 46665 7791 46699
rect 12909 46665 12943 46699
rect 21005 46665 21039 46699
rect 24041 46665 24075 46699
rect 26433 46665 26467 46699
rect 35357 46665 35391 46699
rect 45661 46665 45695 46699
rect 4506 46597 4540 46631
rect 6622 46597 6656 46631
rect 11796 46597 11830 46631
rect 15016 46597 15050 46631
rect 17040 46597 17074 46631
rect 22928 46597 22962 46631
rect 32404 46597 32438 46631
rect 34244 46597 34278 46631
rect 37556 46597 37590 46631
rect 39396 46597 39430 46631
rect 47860 46597 47894 46631
rect 50436 46597 50470 46631
rect 2688 46529 2722 46563
rect 4261 46529 4295 46563
rect 8473 46529 8507 46563
rect 14749 46529 14783 46563
rect 16773 46529 16807 46563
rect 19625 46529 19659 46563
rect 19892 46529 19926 46563
rect 22661 46529 22695 46563
rect 25053 46529 25087 46563
rect 25320 46529 25354 46563
rect 29092 46529 29126 46563
rect 32137 46529 32171 46563
rect 33977 46529 34011 46563
rect 37289 46529 37323 46563
rect 39129 46529 39163 46563
rect 42441 46529 42475 46563
rect 42708 46529 42742 46563
rect 44537 46529 44571 46563
rect 47593 46529 47627 46563
rect 50169 46529 50203 46563
rect 53665 46529 53699 46563
rect 53932 46529 53966 46563
rect 55864 46529 55898 46563
rect 2421 46461 2455 46495
rect 6377 46461 6411 46495
rect 8217 46461 8251 46495
rect 11529 46461 11563 46495
rect 28825 46461 28859 46495
rect 44281 46461 44315 46495
rect 55597 46461 55631 46495
rect 38669 46393 38703 46427
rect 9597 46325 9631 46359
rect 16129 46325 16163 46359
rect 18153 46325 18187 46359
rect 30205 46325 30239 46359
rect 33517 46325 33551 46359
rect 40509 46325 40543 46359
rect 43821 46325 43855 46359
rect 48973 46325 49007 46359
rect 51549 46325 51583 46359
rect 55045 46325 55079 46359
rect 56977 46325 57011 46359
rect 3249 46121 3283 46155
rect 5917 46121 5951 46155
rect 7849 46121 7883 46155
rect 12173 46121 12207 46155
rect 21097 46121 21131 46155
rect 23857 46121 23891 46155
rect 26249 46121 26283 46155
rect 29009 46121 29043 46155
rect 33517 46121 33551 46155
rect 37013 46121 37047 46155
rect 38853 46121 38887 46155
rect 43821 46121 43855 46155
rect 46397 46121 46431 46155
rect 51917 46121 51951 46155
rect 56701 46121 56735 46155
rect 1869 45985 1903 46019
rect 4537 45985 4571 46019
rect 6469 45985 6503 46019
rect 16681 45985 16715 46019
rect 19717 45985 19751 46019
rect 24869 45985 24903 46019
rect 27629 45985 27663 46019
rect 30297 45985 30331 46019
rect 35633 45985 35667 46019
rect 37473 45985 37507 46019
rect 45017 45985 45051 46019
rect 50537 45985 50571 46019
rect 55321 45985 55355 46019
rect 4804 45917 4838 45951
rect 6736 45917 6770 45951
rect 8953 45917 8987 45951
rect 10793 45917 10827 45951
rect 14381 45917 14415 45951
rect 14648 45917 14682 45951
rect 16948 45917 16982 45951
rect 22477 45917 22511 45951
rect 22744 45917 22778 45951
rect 27896 45917 27930 45951
rect 32137 45917 32171 45951
rect 32404 45917 32438 45951
rect 35900 45917 35934 45951
rect 37740 45917 37774 45951
rect 40601 45917 40635 45951
rect 40857 45917 40891 45951
rect 42441 45917 42475 45951
rect 42708 45917 42742 45951
rect 46857 45917 46891 45951
rect 47124 45917 47158 45951
rect 50804 45917 50838 45951
rect 52377 45917 52411 45951
rect 2136 45849 2170 45883
rect 9198 45849 9232 45883
rect 11060 45849 11094 45883
rect 19984 45849 20018 45883
rect 25114 45849 25148 45883
rect 30564 45849 30598 45883
rect 45284 45849 45318 45883
rect 52644 45849 52678 45883
rect 55588 45849 55622 45883
rect 10333 45781 10367 45815
rect 15761 45781 15795 45815
rect 18061 45781 18095 45815
rect 31677 45781 31711 45815
rect 41981 45781 42015 45815
rect 48237 45781 48271 45815
rect 53757 45781 53791 45815
rect 5089 45577 5123 45611
rect 8585 45577 8619 45611
rect 12909 45577 12943 45611
rect 21281 45577 21315 45611
rect 45661 45577 45695 45611
rect 55965 45577 55999 45611
rect 9312 45509 9346 45543
rect 14372 45509 14406 45543
rect 16948 45509 16982 45543
rect 42708 45509 42742 45543
rect 44548 45509 44582 45543
rect 47860 45509 47894 45543
rect 2136 45441 2170 45475
rect 3965 45441 3999 45475
rect 7472 45441 7506 45475
rect 11529 45441 11563 45475
rect 11796 45441 11830 45475
rect 14105 45441 14139 45475
rect 19901 45441 19935 45475
rect 20168 45441 20202 45475
rect 22100 45441 22134 45475
rect 24317 45441 24351 45475
rect 24584 45441 24618 45475
rect 28632 45441 28666 45475
rect 30472 45441 30506 45475
rect 33784 45441 33818 45475
rect 35357 45441 35391 45475
rect 35624 45441 35658 45475
rect 38292 45441 38326 45475
rect 39865 45441 39899 45475
rect 40132 45441 40166 45475
rect 42441 45441 42475 45475
rect 44281 45441 44315 45475
rect 47593 45441 47627 45475
rect 50528 45441 50562 45475
rect 53012 45441 53046 45475
rect 54841 45441 54875 45475
rect 1869 45373 1903 45407
rect 3709 45373 3743 45407
rect 7205 45373 7239 45407
rect 9045 45373 9079 45407
rect 16681 45373 16715 45407
rect 21833 45373 21867 45407
rect 28365 45373 28399 45407
rect 30205 45373 30239 45407
rect 33517 45373 33551 45407
rect 38025 45373 38059 45407
rect 50261 45373 50295 45407
rect 52745 45373 52779 45407
rect 54585 45373 54619 45407
rect 3249 45305 3283 45339
rect 18061 45305 18095 45339
rect 41245 45305 41279 45339
rect 43821 45305 43855 45339
rect 54125 45305 54159 45339
rect 10425 45237 10459 45271
rect 15485 45237 15519 45271
rect 23213 45237 23247 45271
rect 25697 45237 25731 45271
rect 29745 45237 29779 45271
rect 31585 45237 31619 45271
rect 34897 45237 34931 45271
rect 36737 45237 36771 45271
rect 39405 45237 39439 45271
rect 48973 45237 49007 45271
rect 51641 45237 51675 45271
rect 3157 45033 3191 45067
rect 21373 45033 21407 45067
rect 23213 45033 23247 45067
rect 29009 45033 29043 45067
rect 31677 45033 31711 45067
rect 51549 45033 51583 45067
rect 53389 45033 53423 45067
rect 56701 45033 56735 45067
rect 16865 44897 16899 44931
rect 19993 44897 20027 44931
rect 45753 44897 45787 44931
rect 47593 44897 47627 44931
rect 57161 44897 57195 44931
rect 1777 44829 1811 44863
rect 6377 44829 6411 44863
rect 8953 44829 8987 44863
rect 10793 44829 10827 44863
rect 14105 44829 14139 44863
rect 14372 44829 14406 44863
rect 20260 44829 20294 44863
rect 21833 44829 21867 44863
rect 25789 44829 25823 44863
rect 27629 44829 27663 44863
rect 27896 44829 27930 44863
rect 30297 44829 30331 44863
rect 32137 44829 32171 44863
rect 36093 44829 36127 44863
rect 37933 44829 37967 44863
rect 40601 44829 40635 44863
rect 42441 44829 42475 44863
rect 47860 44829 47894 44863
rect 50169 44829 50203 44863
rect 52009 44829 52043 44863
rect 55321 44829 55355 44863
rect 57417 44829 57451 44863
rect 2044 44761 2078 44795
rect 6644 44761 6678 44795
rect 9220 44761 9254 44795
rect 11038 44761 11072 44795
rect 17132 44761 17166 44795
rect 22100 44761 22134 44795
rect 26056 44761 26090 44795
rect 30564 44761 30598 44795
rect 32404 44761 32438 44795
rect 36360 44761 36394 44795
rect 38200 44761 38234 44795
rect 40868 44761 40902 44795
rect 42708 44761 42742 44795
rect 46020 44761 46054 44795
rect 50436 44761 50470 44795
rect 52276 44761 52310 44795
rect 55588 44761 55622 44795
rect 7757 44693 7791 44727
rect 10333 44693 10367 44727
rect 12173 44693 12207 44727
rect 15485 44693 15519 44727
rect 18245 44693 18279 44727
rect 27169 44693 27203 44727
rect 33517 44693 33551 44727
rect 37473 44693 37507 44727
rect 39313 44693 39347 44727
rect 41981 44693 42015 44727
rect 43821 44693 43855 44727
rect 47133 44693 47167 44727
rect 48973 44693 49007 44727
rect 58541 44693 58575 44727
rect 3065 44489 3099 44523
rect 7757 44489 7791 44523
rect 9597 44489 9631 44523
rect 12909 44489 12943 44523
rect 23213 44489 23247 44523
rect 31585 44489 31619 44523
rect 54125 44489 54159 44523
rect 55965 44489 55999 44523
rect 8484 44421 8518 44455
rect 11796 44421 11830 44455
rect 13912 44421 13946 44455
rect 17224 44421 17258 44455
rect 28632 44421 28666 44455
rect 33784 44421 33818 44455
rect 40776 44421 40810 44455
rect 47860 44421 47894 44455
rect 53012 44421 53046 44455
rect 54852 44421 54886 44455
rect 1685 44353 1719 44387
rect 1952 44353 1986 44387
rect 4353 44353 4387 44387
rect 4620 44353 4654 44387
rect 6644 44353 6678 44387
rect 8217 44353 8251 44387
rect 13645 44353 13679 44387
rect 16957 44353 16991 44387
rect 21833 44353 21867 44387
rect 22100 44353 22134 44387
rect 25053 44353 25087 44387
rect 25320 44353 25354 44387
rect 30205 44353 30239 44387
rect 30472 44353 30506 44387
rect 35357 44353 35391 44387
rect 35624 44353 35658 44387
rect 38936 44353 38970 44387
rect 43085 44353 43119 44387
rect 43352 44353 43386 44387
rect 45652 44353 45686 44387
rect 47593 44353 47627 44387
rect 49689 44353 49723 44387
rect 52745 44353 52779 44387
rect 54585 44353 54619 44387
rect 6377 44285 6411 44319
rect 11529 44285 11563 44319
rect 28365 44285 28399 44319
rect 33517 44285 33551 44319
rect 38669 44285 38703 44319
rect 40509 44285 40543 44319
rect 45385 44285 45419 44319
rect 49433 44285 49467 44319
rect 48973 44217 49007 44251
rect 5733 44149 5767 44183
rect 15025 44149 15059 44183
rect 18337 44149 18371 44183
rect 26433 44149 26467 44183
rect 29745 44149 29779 44183
rect 34897 44149 34931 44183
rect 36737 44149 36771 44183
rect 40049 44149 40083 44183
rect 41889 44149 41923 44183
rect 44465 44149 44499 44183
rect 46765 44149 46799 44183
rect 50813 44149 50847 44183
rect 6929 43945 6963 43979
rect 23857 43945 23891 43979
rect 27077 43945 27111 43979
rect 28917 43945 28951 43979
rect 32229 43945 32263 43979
rect 36369 43945 36403 43979
rect 39313 43945 39347 43979
rect 42625 43945 42659 43979
rect 46673 43945 46707 43979
rect 53389 43945 53423 43979
rect 44465 43877 44499 43911
rect 1869 43809 1903 43843
rect 14105 43809 14139 43843
rect 17141 43809 17175 43843
rect 25697 43809 25731 43843
rect 30849 43809 30883 43843
rect 43085 43809 43119 43843
rect 56517 43809 56551 43843
rect 2136 43741 2170 43775
rect 9597 43741 9631 43775
rect 12173 43741 12207 43775
rect 14372 43741 14406 43775
rect 17408 43741 17442 43775
rect 22477 43741 22511 43775
rect 25964 43741 25998 43775
rect 27537 43741 27571 43775
rect 27804 43741 27838 43775
rect 31116 43741 31150 43775
rect 32781 43741 32815 43775
rect 33048 43741 33082 43775
rect 37933 43741 37967 43775
rect 38200 43741 38234 43775
rect 41245 43741 41279 43775
rect 41512 43741 41546 43775
rect 45293 43741 45327 43775
rect 50169 43741 50203 43775
rect 52009 43741 52043 43775
rect 52265 43741 52299 43775
rect 56784 43741 56818 43775
rect 5641 43673 5675 43707
rect 9864 43673 9898 43707
rect 12440 43673 12474 43707
rect 20269 43673 20303 43707
rect 22744 43673 22778 43707
rect 35081 43673 35115 43707
rect 43352 43673 43386 43707
rect 45560 43673 45594 43707
rect 47869 43673 47903 43707
rect 50414 43673 50448 43707
rect 3249 43605 3283 43639
rect 10977 43605 11011 43639
rect 13553 43605 13587 43639
rect 15485 43605 15519 43639
rect 18521 43605 18555 43639
rect 21557 43605 21591 43639
rect 34161 43605 34195 43639
rect 49157 43605 49191 43639
rect 51549 43605 51583 43639
rect 57897 43605 57931 43639
rect 3065 43401 3099 43435
rect 5365 43401 5399 43435
rect 7757 43401 7791 43435
rect 14841 43401 14875 43435
rect 23213 43401 23247 43435
rect 25789 43401 25823 43435
rect 30481 43401 30515 43435
rect 34897 43401 34931 43435
rect 38761 43401 38795 43435
rect 46489 43401 46523 43435
rect 49617 43401 49651 43435
rect 54585 43401 54619 43435
rect 1952 43333 1986 43367
rect 6622 43333 6656 43367
rect 13728 43333 13762 43367
rect 17500 43333 17534 43367
rect 24501 43333 24535 43367
rect 29368 43333 29402 43367
rect 33784 43333 33818 43367
rect 35624 43333 35658 43367
rect 37648 43333 37682 43367
rect 42708 43333 42742 43367
rect 48504 43333 48538 43367
rect 50344 43333 50378 43367
rect 1685 43265 1719 43299
rect 4252 43265 4286 43299
rect 6377 43265 6411 43299
rect 9864 43265 9898 43299
rect 11888 43265 11922 43299
rect 13461 43265 13495 43299
rect 17233 43265 17267 43299
rect 19257 43265 19291 43299
rect 19513 43265 19547 43299
rect 21833 43265 21867 43299
rect 22100 43265 22134 43299
rect 27261 43265 27295 43299
rect 27528 43265 27562 43299
rect 29101 43265 29135 43299
rect 33517 43265 33551 43299
rect 35357 43265 35391 43299
rect 39221 43265 39255 43299
rect 45109 43265 45143 43299
rect 45376 43265 45410 43299
rect 48237 43265 48271 43299
rect 50077 43265 50111 43299
rect 53113 43265 53147 43299
rect 55965 43265 55999 43299
rect 56232 43265 56266 43299
rect 3985 43197 4019 43231
rect 9597 43197 9631 43231
rect 11621 43197 11655 43231
rect 37381 43197 37415 43231
rect 42441 43197 42475 43231
rect 36737 43129 36771 43163
rect 10977 43061 11011 43095
rect 13001 43061 13035 43095
rect 18613 43061 18647 43095
rect 20637 43061 20671 43095
rect 28641 43061 28675 43095
rect 40509 43061 40543 43095
rect 43821 43061 43855 43095
rect 51457 43061 51491 43095
rect 57345 43061 57379 43095
rect 5181 42857 5215 42891
rect 11529 42857 11563 42891
rect 23673 42857 23707 42891
rect 46397 42857 46431 42891
rect 58173 42857 58207 42891
rect 7021 42721 7055 42755
rect 17325 42721 17359 42755
rect 20453 42721 20487 42755
rect 47593 42721 47627 42755
rect 50169 42721 50203 42755
rect 53389 42721 53423 42755
rect 56793 42721 56827 42755
rect 3801 42653 3835 42687
rect 10241 42653 10275 42687
rect 15485 42653 15519 42687
rect 17592 42653 17626 42687
rect 22293 42653 22327 42687
rect 24409 42653 24443 42687
rect 24676 42653 24710 42687
rect 30849 42653 30883 42687
rect 31116 42653 31150 42687
rect 32689 42653 32723 42687
rect 32956 42653 32990 42687
rect 35357 42653 35391 42687
rect 35624 42653 35658 42687
rect 37933 42653 37967 42687
rect 38200 42653 38234 42687
rect 40509 42653 40543 42687
rect 40776 42653 40810 42687
rect 42349 42653 42383 42687
rect 45017 42653 45051 42687
rect 47860 42653 47894 42687
rect 50436 42653 50470 42687
rect 57060 42653 57094 42687
rect 4068 42585 4102 42619
rect 7288 42585 7322 42619
rect 15752 42585 15786 42619
rect 20720 42585 20754 42619
rect 22538 42585 22572 42619
rect 27261 42585 27295 42619
rect 42616 42585 42650 42619
rect 45284 42585 45318 42619
rect 53656 42585 53690 42619
rect 8401 42517 8435 42551
rect 16865 42517 16899 42551
rect 18705 42517 18739 42551
rect 21833 42517 21867 42551
rect 25789 42517 25823 42551
rect 28549 42517 28583 42551
rect 32229 42517 32263 42551
rect 34069 42517 34103 42551
rect 36737 42517 36771 42551
rect 39313 42517 39347 42551
rect 41889 42517 41923 42551
rect 43729 42517 43763 42551
rect 48973 42517 49007 42551
rect 51549 42517 51583 42551
rect 54769 42517 54803 42551
rect 10977 42313 11011 42347
rect 14289 42313 14323 42347
rect 18797 42313 18831 42347
rect 21281 42313 21315 42347
rect 24041 42313 24075 42347
rect 29101 42313 29135 42347
rect 44465 42313 44499 42347
rect 46765 42313 46799 42347
rect 55137 42313 55171 42347
rect 56885 42313 56919 42347
rect 7472 42245 7506 42279
rect 13176 42245 13210 42279
rect 17684 42245 17718 42279
rect 22928 42245 22962 42279
rect 55597 42245 55631 42279
rect 3148 42177 3182 42211
rect 7205 42177 7239 42211
rect 9864 42177 9898 42211
rect 12909 42177 12943 42211
rect 14749 42177 14783 42211
rect 15016 42177 15050 42211
rect 19901 42177 19935 42211
rect 20168 42177 20202 42211
rect 22661 42177 22695 42211
rect 24501 42177 24535 42211
rect 24768 42177 24802 42211
rect 27988 42177 28022 42211
rect 34969 42177 35003 42211
rect 38761 42177 38795 42211
rect 39028 42177 39062 42211
rect 43177 42177 43211 42211
rect 45385 42177 45419 42211
rect 45652 42177 45686 42211
rect 48973 42177 49007 42211
rect 49240 42177 49274 42211
rect 50813 42177 50847 42211
rect 51080 42177 51114 42211
rect 54024 42177 54058 42211
rect 2881 42109 2915 42143
rect 9597 42109 9631 42143
rect 17417 42109 17451 42143
rect 27721 42109 27755 42143
rect 34713 42109 34747 42143
rect 53757 42109 53791 42143
rect 4261 41973 4295 42007
rect 8585 41973 8619 42007
rect 16129 41973 16163 42007
rect 25881 41973 25915 42007
rect 36093 41973 36127 42007
rect 40141 41973 40175 42007
rect 50353 41973 50387 42007
rect 52193 41973 52227 42007
rect 5181 41769 5215 41803
rect 8401 41769 8435 41803
rect 11621 41769 11655 41803
rect 21557 41769 21591 41803
rect 29009 41769 29043 41803
rect 41889 41769 41923 41803
rect 43821 41769 43855 41803
rect 46397 41769 46431 41803
rect 7021 41633 7055 41667
rect 12081 41633 12115 41667
rect 20177 41633 20211 41667
rect 22477 41633 22511 41667
rect 35357 41633 35391 41667
rect 45017 41633 45051 41667
rect 3801 41565 3835 41599
rect 4068 41565 4102 41599
rect 7288 41565 7322 41599
rect 10241 41565 10275 41599
rect 12348 41565 12382 41599
rect 14473 41565 14507 41599
rect 17325 41565 17359 41599
rect 17592 41565 17626 41599
rect 25789 41565 25823 41599
rect 26056 41565 26090 41599
rect 27629 41565 27663 41599
rect 29561 41565 29595 41599
rect 32137 41565 32171 41599
rect 37841 41565 37875 41599
rect 40509 41565 40543 41599
rect 40776 41565 40810 41599
rect 42441 41565 42475 41599
rect 47685 41565 47719 41599
rect 51549 41565 51583 41599
rect 53389 41565 53423 41599
rect 53656 41565 53690 41599
rect 55965 41565 55999 41599
rect 56232 41565 56266 41599
rect 10508 41497 10542 41531
rect 20444 41497 20478 41531
rect 22744 41497 22778 41531
rect 27896 41497 27930 41531
rect 29828 41497 29862 41531
rect 32404 41497 32438 41531
rect 35624 41497 35658 41531
rect 38108 41497 38142 41531
rect 42708 41497 42742 41531
rect 45284 41497 45318 41531
rect 47952 41497 47986 41531
rect 51816 41497 51850 41531
rect 13461 41429 13495 41463
rect 15761 41429 15795 41463
rect 18705 41429 18739 41463
rect 23857 41429 23891 41463
rect 27169 41429 27203 41463
rect 30941 41429 30975 41463
rect 33517 41429 33551 41463
rect 36737 41429 36771 41463
rect 39221 41429 39255 41463
rect 49065 41429 49099 41463
rect 52929 41429 52963 41463
rect 54769 41429 54803 41463
rect 57345 41429 57379 41463
rect 3617 41225 3651 41259
rect 5457 41225 5491 41259
rect 21281 41225 21315 41259
rect 29653 41225 29687 41259
rect 36737 41225 36771 41259
rect 43821 41225 43855 41259
rect 46581 41225 46615 41259
rect 50353 41225 50387 41259
rect 54401 41225 54435 41259
rect 4322 41157 4356 41191
rect 6736 41157 6770 41191
rect 9496 41157 9530 41191
rect 15016 41157 15050 41191
rect 17960 41157 17994 41191
rect 23480 41157 23514 41191
rect 51080 41157 51114 41191
rect 53288 41157 53322 41191
rect 55956 41157 55990 41191
rect 2237 41089 2271 41123
rect 2504 41089 2538 41123
rect 12909 41089 12943 41123
rect 13176 41089 13210 41123
rect 19901 41089 19935 41123
rect 20168 41089 20202 41123
rect 23213 41089 23247 41123
rect 25320 41089 25354 41123
rect 28540 41089 28574 41123
rect 30472 41089 30506 41123
rect 32772 41089 32806 41123
rect 35357 41089 35391 41123
rect 35624 41089 35658 41123
rect 38936 41089 38970 41123
rect 40776 41089 40810 41123
rect 42708 41089 42742 41123
rect 45201 41089 45235 41123
rect 45468 41089 45502 41123
rect 48973 41089 49007 41123
rect 49240 41089 49274 41123
rect 55689 41089 55723 41123
rect 4077 41021 4111 41055
rect 6469 41021 6503 41055
rect 9229 41021 9263 41055
rect 14749 41021 14783 41055
rect 17693 41021 17727 41055
rect 25053 41021 25087 41055
rect 28273 41021 28307 41055
rect 30205 41021 30239 41055
rect 32505 41021 32539 41055
rect 38669 41021 38703 41055
rect 40509 41021 40543 41055
rect 42441 41021 42475 41055
rect 50813 41021 50847 41055
rect 53021 41021 53055 41055
rect 16129 40953 16163 40987
rect 7849 40885 7883 40919
rect 10609 40885 10643 40919
rect 14289 40885 14323 40919
rect 19073 40885 19107 40919
rect 24593 40885 24627 40919
rect 26433 40885 26467 40919
rect 31585 40885 31619 40919
rect 33885 40885 33919 40919
rect 40049 40885 40083 40919
rect 41889 40885 41923 40919
rect 52193 40885 52227 40919
rect 57069 40885 57103 40919
rect 3249 40681 3283 40715
rect 10977 40681 11011 40715
rect 12817 40681 12851 40715
rect 18705 40681 18739 40715
rect 23857 40681 23891 40715
rect 27169 40681 27203 40715
rect 29009 40681 29043 40715
rect 41797 40681 41831 40715
rect 43821 40681 43855 40715
rect 46397 40681 46431 40715
rect 53665 40681 53699 40715
rect 56701 40681 56735 40715
rect 15301 40545 15335 40579
rect 25789 40545 25823 40579
rect 30573 40545 30607 40579
rect 37933 40545 37967 40579
rect 40417 40545 40451 40579
rect 45017 40545 45051 40579
rect 50445 40545 50479 40579
rect 52285 40545 52319 40579
rect 55321 40545 55355 40579
rect 1869 40477 1903 40511
rect 6193 40477 6227 40511
rect 6460 40477 6494 40511
rect 9597 40477 9631 40511
rect 9864 40477 9898 40511
rect 11437 40477 11471 40511
rect 11693 40477 11727 40511
rect 15568 40477 15602 40511
rect 17325 40477 17359 40511
rect 17592 40477 17626 40511
rect 22477 40477 22511 40511
rect 22744 40477 22778 40511
rect 26056 40477 26090 40511
rect 27629 40477 27663 40511
rect 30840 40477 30874 40511
rect 36093 40477 36127 40511
rect 36360 40477 36394 40511
rect 38200 40477 38234 40511
rect 42441 40477 42475 40511
rect 45273 40477 45307 40511
rect 48237 40477 48271 40511
rect 48504 40477 48538 40511
rect 50712 40477 50746 40511
rect 52552 40477 52586 40511
rect 55588 40477 55622 40511
rect 2136 40409 2170 40443
rect 19625 40409 19659 40443
rect 27896 40409 27930 40443
rect 32413 40409 32447 40443
rect 34161 40409 34195 40443
rect 40684 40409 40718 40443
rect 42708 40409 42742 40443
rect 7573 40341 7607 40375
rect 16681 40341 16715 40375
rect 21097 40341 21131 40375
rect 31953 40341 31987 40375
rect 37473 40341 37507 40375
rect 39313 40341 39347 40375
rect 49617 40341 49651 40375
rect 51825 40341 51859 40375
rect 18061 40137 18095 40171
rect 21281 40137 21315 40171
rect 26157 40137 26191 40171
rect 29745 40137 29779 40171
rect 31585 40137 31619 40171
rect 36737 40137 36771 40171
rect 40785 40137 40819 40171
rect 43821 40137 43855 40171
rect 51549 40137 51583 40171
rect 4077 40069 4111 40103
rect 47961 40069 47995 40103
rect 2237 40001 2271 40035
rect 2504 40001 2538 40035
rect 6377 40001 6411 40035
rect 6644 40001 6678 40035
rect 8473 40001 8507 40035
rect 12173 40001 12207 40035
rect 12440 40001 12474 40035
rect 14749 40001 14783 40035
rect 15016 40001 15050 40035
rect 16681 40001 16715 40035
rect 16948 40001 16982 40035
rect 19901 40001 19935 40035
rect 20168 40001 20202 40035
rect 23204 40001 23238 40035
rect 24777 40001 24811 40035
rect 25044 40001 25078 40035
rect 28365 40001 28399 40035
rect 28632 40001 28666 40035
rect 30472 40001 30506 40035
rect 32781 40001 32815 40035
rect 33048 40001 33082 40035
rect 35357 40001 35391 40035
rect 35624 40001 35658 40035
rect 37832 40001 37866 40035
rect 39405 40001 39439 40035
rect 39672 40001 39706 40035
rect 42441 40001 42475 40035
rect 42708 40001 42742 40035
rect 45661 40001 45695 40035
rect 45928 40001 45962 40035
rect 50169 40001 50203 40035
rect 50436 40001 50470 40035
rect 5825 39933 5859 39967
rect 8217 39933 8251 39967
rect 22937 39933 22971 39967
rect 30205 39933 30239 39967
rect 37565 39933 37599 39967
rect 3617 39797 3651 39831
rect 7757 39797 7791 39831
rect 9597 39797 9631 39831
rect 13553 39797 13587 39831
rect 16129 39797 16163 39831
rect 24317 39797 24351 39831
rect 34161 39797 34195 39831
rect 38945 39797 38979 39831
rect 47041 39797 47075 39831
rect 49249 39797 49283 39831
rect 3249 39593 3283 39627
rect 5181 39593 5215 39627
rect 7757 39593 7791 39627
rect 11529 39593 11563 39627
rect 18061 39593 18095 39627
rect 27169 39593 27203 39627
rect 32321 39593 32355 39627
rect 34161 39593 34195 39627
rect 37473 39593 37507 39627
rect 39313 39593 39347 39627
rect 40325 39593 40359 39627
rect 43821 39593 43855 39627
rect 47777 39593 47811 39627
rect 8953 39457 8987 39491
rect 12173 39457 12207 39491
rect 32781 39457 32815 39491
rect 36093 39457 36127 39491
rect 37933 39457 37967 39491
rect 42441 39457 42475 39491
rect 48237 39457 48271 39491
rect 1869 39389 1903 39423
rect 2136 39389 2170 39423
rect 3801 39389 3835 39423
rect 6377 39389 6411 39423
rect 6644 39389 6678 39423
rect 11713 39389 11747 39423
rect 12440 39389 12474 39423
rect 14197 39389 14231 39423
rect 14464 39389 14498 39423
rect 16681 39389 16715 39423
rect 19257 39389 19291 39423
rect 19513 39389 19547 39423
rect 22477 39389 22511 39423
rect 22744 39389 22778 39423
rect 25789 39389 25823 39423
rect 27629 39389 27663 39423
rect 30941 39389 30975 39423
rect 31208 39389 31242 39423
rect 33048 39389 33082 39423
rect 36360 39389 36394 39423
rect 38200 39389 38234 39423
rect 40509 39389 40543 39423
rect 46397 39389 46431 39423
rect 48504 39389 48538 39423
rect 50905 39389 50939 39423
rect 52745 39389 52779 39423
rect 4068 39321 4102 39355
rect 9198 39321 9232 39355
rect 16948 39321 16982 39355
rect 26056 39321 26090 39355
rect 27896 39321 27930 39355
rect 42708 39321 42742 39355
rect 46664 39321 46698 39355
rect 51172 39321 51206 39355
rect 53012 39321 53046 39355
rect 10333 39253 10367 39287
rect 13553 39253 13587 39287
rect 15577 39253 15611 39287
rect 20637 39253 20671 39287
rect 23857 39253 23891 39287
rect 29009 39253 29043 39287
rect 49617 39253 49651 39287
rect 52285 39253 52319 39287
rect 54125 39253 54159 39287
rect 8493 39049 8527 39083
rect 18337 39049 18371 39083
rect 24225 39049 24259 39083
rect 28365 39049 28399 39083
rect 31585 39049 31619 39083
rect 34253 39049 34287 39083
rect 40233 39049 40267 39083
rect 43821 39049 43855 39083
rect 49341 39049 49375 39083
rect 56701 39049 56735 39083
rect 7380 38981 7414 39015
rect 9220 38981 9254 39015
rect 12440 38981 12474 39015
rect 19064 38981 19098 39015
rect 23112 38981 23146 39015
rect 30472 38981 30506 39015
rect 33140 38981 33174 39015
rect 39120 38981 39154 39015
rect 45652 38981 45686 39015
rect 48228 38981 48262 39015
rect 53748 38981 53782 39015
rect 4068 38913 4102 38947
rect 7113 38913 7147 38947
rect 8953 38913 8987 38947
rect 12173 38913 12207 38947
rect 17224 38913 17258 38947
rect 20821 38913 20855 38947
rect 22845 38913 22879 38947
rect 26985 38913 27019 38947
rect 27252 38913 27286 38947
rect 30205 38913 30239 38947
rect 32873 38913 32907 38947
rect 34980 38913 35014 38947
rect 38853 38913 38887 38947
rect 42708 38913 42742 38947
rect 45385 38913 45419 38947
rect 49985 38913 50019 38947
rect 50537 38913 50571 38947
rect 50804 38913 50838 38947
rect 53481 38913 53515 38947
rect 55588 38913 55622 38947
rect 3801 38845 3835 38879
rect 16957 38845 16991 38879
rect 18797 38845 18831 38879
rect 34713 38845 34747 38879
rect 42441 38845 42475 38879
rect 47961 38845 47995 38879
rect 55321 38845 55355 38879
rect 5181 38709 5215 38743
rect 10333 38709 10367 38743
rect 13553 38709 13587 38743
rect 20177 38709 20211 38743
rect 20637 38709 20671 38743
rect 36093 38709 36127 38743
rect 46765 38709 46799 38743
rect 49801 38709 49835 38743
rect 51917 38709 51951 38743
rect 54861 38709 54895 38743
rect 27629 38505 27663 38539
rect 31125 38505 31159 38539
rect 36093 38505 36127 38539
rect 46857 38505 46891 38539
rect 52929 38505 52963 38539
rect 56701 38505 56735 38539
rect 47501 38369 47535 38403
rect 53389 38369 53423 38403
rect 4997 38301 5031 38335
rect 8953 38301 8987 38335
rect 9220 38301 9254 38335
rect 12081 38301 12115 38335
rect 12348 38301 12382 38335
rect 14657 38301 14691 38335
rect 16497 38301 16531 38335
rect 19257 38301 19291 38335
rect 19524 38301 19558 38335
rect 21097 38301 21131 38335
rect 24409 38301 24443 38335
rect 26249 38301 26283 38335
rect 29745 38301 29779 38335
rect 30012 38301 30046 38335
rect 32505 38301 32539 38335
rect 34713 38301 34747 38335
rect 36553 38301 36587 38335
rect 42901 38301 42935 38335
rect 45477 38301 45511 38335
rect 45744 38301 45778 38335
rect 51549 38301 51583 38335
rect 53656 38301 53690 38335
rect 55321 38301 55355 38335
rect 5264 38233 5298 38267
rect 14924 38233 14958 38267
rect 16764 38233 16798 38267
rect 21364 38233 21398 38267
rect 24676 38233 24710 38267
rect 26516 38233 26550 38267
rect 32772 38233 32806 38267
rect 34980 38233 35014 38267
rect 36820 38233 36854 38267
rect 43168 38233 43202 38267
rect 47768 38233 47802 38267
rect 51816 38233 51850 38267
rect 55588 38233 55622 38267
rect 6377 38165 6411 38199
rect 10333 38165 10367 38199
rect 13461 38165 13495 38199
rect 16037 38165 16071 38199
rect 17877 38165 17911 38199
rect 20637 38165 20671 38199
rect 22477 38165 22511 38199
rect 25789 38165 25823 38199
rect 33885 38165 33919 38199
rect 37933 38165 37967 38199
rect 44281 38165 44315 38199
rect 48881 38165 48915 38199
rect 54769 38165 54803 38199
rect 3985 37961 4019 37995
rect 5825 37961 5859 37995
rect 15853 37961 15887 37995
rect 18061 37961 18095 37995
rect 28549 37961 28583 37995
rect 30481 37961 30515 37995
rect 33517 37961 33551 37995
rect 35357 37961 35391 37995
rect 44465 37961 44499 37995
rect 4712 37893 4746 37927
rect 8668 37893 8702 37927
rect 12072 37893 12106 37927
rect 16948 37893 16982 37927
rect 18788 37893 18822 37927
rect 27436 37893 27470 37927
rect 49240 37893 49274 37927
rect 51080 37893 51114 37927
rect 54769 37893 54803 37927
rect 2872 37825 2906 37859
rect 14473 37825 14507 37859
rect 14740 37825 14774 37859
rect 18521 37825 18555 37859
rect 21833 37825 21867 37859
rect 22100 37825 22134 37859
rect 23673 37825 23707 37859
rect 23940 37825 23974 37859
rect 29368 37825 29402 37859
rect 32404 37825 32438 37859
rect 33977 37825 34011 37859
rect 34244 37825 34278 37859
rect 37289 37825 37323 37859
rect 37556 37825 37590 37859
rect 39129 37825 39163 37859
rect 39396 37825 39430 37859
rect 43085 37825 43119 37859
rect 43352 37825 43386 37859
rect 45836 37825 45870 37859
rect 48973 37825 49007 37859
rect 2605 37757 2639 37791
rect 4445 37757 4479 37791
rect 8401 37757 8435 37791
rect 11805 37757 11839 37791
rect 16681 37757 16715 37791
rect 27169 37757 27203 37791
rect 29101 37757 29135 37791
rect 32137 37757 32171 37791
rect 45569 37757 45603 37791
rect 50813 37757 50847 37791
rect 9781 37621 9815 37655
rect 13185 37621 13219 37655
rect 19901 37621 19935 37655
rect 23213 37621 23247 37655
rect 25053 37621 25087 37655
rect 38669 37621 38703 37655
rect 40509 37621 40543 37655
rect 46949 37621 46983 37655
rect 50353 37621 50387 37655
rect 52193 37621 52227 37655
rect 56057 37621 56091 37655
rect 18061 37417 18095 37451
rect 22477 37417 22511 37451
rect 27629 37417 27663 37451
rect 30941 37417 30975 37451
rect 33149 37417 33183 37451
rect 37933 37417 37967 37451
rect 42533 37417 42567 37451
rect 56701 37417 56735 37451
rect 8953 37281 8987 37315
rect 14841 37281 14875 37315
rect 34713 37281 34747 37315
rect 48237 37281 48271 37315
rect 5181 37213 5215 37247
rect 7021 37213 7055 37247
rect 9220 37213 9254 37247
rect 11529 37213 11563 37247
rect 11796 37213 11830 37247
rect 16681 37213 16715 37247
rect 16948 37213 16982 37247
rect 19257 37213 19291 37247
rect 19524 37213 19558 37247
rect 21097 37213 21131 37247
rect 24409 37213 24443 37247
rect 24676 37213 24710 37247
rect 26238 37213 26272 37247
rect 26505 37213 26539 37247
rect 29561 37213 29595 37247
rect 29817 37213 29851 37247
rect 31769 37213 31803 37247
rect 34969 37213 35003 37247
rect 36553 37213 36587 37247
rect 36809 37213 36843 37247
rect 41245 37213 41279 37247
rect 46397 37213 46431 37247
rect 46664 37213 46698 37247
rect 51549 37213 51583 37247
rect 53389 37213 53423 37247
rect 55321 37213 55355 37247
rect 5448 37145 5482 37179
rect 7288 37145 7322 37179
rect 15108 37145 15142 37179
rect 21342 37145 21376 37179
rect 32036 37145 32070 37179
rect 48504 37145 48538 37179
rect 51816 37145 51850 37179
rect 53656 37145 53690 37179
rect 55588 37145 55622 37179
rect 6561 37077 6595 37111
rect 8401 37077 8435 37111
rect 10333 37077 10367 37111
rect 12909 37077 12943 37111
rect 16221 37077 16255 37111
rect 20637 37077 20671 37111
rect 25789 37077 25823 37111
rect 36093 37077 36127 37111
rect 47777 37077 47811 37111
rect 49617 37077 49651 37111
rect 52929 37077 52963 37111
rect 54769 37077 54803 37111
rect 5825 36873 5859 36907
rect 9781 36873 9815 36907
rect 14841 36873 14875 36907
rect 18061 36873 18095 36907
rect 20269 36873 20303 36907
rect 23213 36873 23247 36907
rect 25053 36873 25087 36907
rect 33517 36873 33551 36907
rect 38669 36873 38703 36907
rect 50353 36873 50387 36907
rect 56425 36873 56459 36907
rect 4712 36805 4746 36839
rect 6828 36805 6862 36839
rect 8668 36805 8702 36839
rect 11796 36805 11830 36839
rect 13553 36805 13587 36839
rect 19156 36805 19190 36839
rect 27353 36805 27387 36839
rect 35624 36805 35658 36839
rect 37556 36805 37590 36839
rect 45928 36805 45962 36839
rect 49240 36805 49274 36839
rect 51080 36805 51114 36839
rect 4445 36737 4479 36771
rect 11529 36737 11563 36771
rect 16681 36737 16715 36771
rect 16948 36737 16982 36771
rect 18889 36737 18923 36771
rect 21833 36737 21867 36771
rect 22100 36737 22134 36771
rect 23940 36737 23974 36771
rect 29561 36737 29595 36771
rect 29828 36737 29862 36771
rect 32404 36737 32438 36771
rect 35357 36737 35391 36771
rect 37289 36737 37323 36771
rect 39385 36737 39419 36771
rect 43821 36737 43855 36771
rect 44088 36737 44122 36771
rect 50813 36737 50847 36771
rect 55045 36737 55079 36771
rect 55312 36737 55346 36771
rect 6561 36669 6595 36703
rect 8401 36669 8435 36703
rect 23673 36669 23707 36703
rect 32137 36669 32171 36703
rect 39129 36669 39163 36703
rect 45661 36669 45695 36703
rect 48973 36669 49007 36703
rect 52193 36601 52227 36635
rect 7941 36533 7975 36567
rect 12909 36533 12943 36567
rect 28825 36533 28859 36567
rect 30941 36533 30975 36567
rect 36737 36533 36771 36567
rect 40509 36533 40543 36567
rect 45201 36533 45235 36567
rect 47041 36533 47075 36567
rect 10333 36329 10367 36363
rect 18061 36329 18095 36363
rect 22477 36329 22511 36363
rect 27629 36329 27663 36363
rect 30941 36329 30975 36363
rect 33609 36329 33643 36363
rect 38669 36329 38703 36363
rect 51549 36329 51583 36363
rect 56701 36329 56735 36363
rect 8953 36193 8987 36227
rect 11529 36193 11563 36227
rect 16681 36193 16715 36227
rect 21097 36193 21131 36227
rect 29561 36193 29595 36227
rect 39865 36193 39899 36227
rect 48237 36193 48271 36227
rect 6561 36125 6595 36159
rect 6828 36125 6862 36159
rect 9209 36125 9243 36159
rect 11796 36125 11830 36159
rect 14105 36125 14139 36159
rect 19257 36125 19291 36159
rect 21364 36125 21398 36159
rect 24409 36125 24443 36159
rect 24676 36125 24710 36159
rect 26249 36125 26283 36159
rect 34897 36125 34931 36159
rect 37289 36125 37323 36159
rect 37556 36125 37590 36159
rect 40132 36125 40166 36159
rect 41705 36125 41739 36159
rect 50176 36125 50210 36159
rect 52009 36125 52043 36159
rect 55321 36125 55355 36159
rect 14350 36057 14384 36091
rect 16948 36057 16982 36091
rect 19524 36057 19558 36091
rect 26494 36057 26528 36091
rect 29828 36057 29862 36091
rect 32321 36057 32355 36091
rect 35164 36057 35198 36091
rect 41950 36057 41984 36091
rect 46489 36057 46523 36091
rect 50414 36057 50448 36091
rect 52254 36057 52288 36091
rect 55588 36057 55622 36091
rect 7941 35989 7975 36023
rect 12909 35989 12943 36023
rect 15485 35989 15519 36023
rect 20637 35989 20671 36023
rect 25789 35989 25823 36023
rect 36277 35989 36311 36023
rect 41245 35989 41279 36023
rect 43085 35989 43119 36023
rect 53389 35989 53423 36023
rect 7757 35785 7791 35819
rect 23213 35785 23247 35819
rect 25053 35785 25087 35819
rect 33517 35785 33551 35819
rect 36093 35785 36127 35819
rect 39405 35785 39439 35819
rect 41337 35785 41371 35819
rect 6644 35717 6678 35751
rect 11796 35717 11830 35751
rect 22100 35717 22134 35751
rect 23918 35717 23952 35751
rect 32404 35717 32438 35751
rect 38292 35717 38326 35751
rect 40224 35717 40258 35751
rect 42686 35717 42720 35751
rect 45928 35717 45962 35751
rect 3985 35649 4019 35683
rect 11529 35649 11563 35683
rect 13625 35649 13659 35683
rect 18245 35649 18279 35683
rect 21833 35649 21867 35683
rect 23673 35649 23707 35683
rect 27344 35649 27378 35683
rect 29184 35649 29218 35683
rect 32137 35649 32171 35683
rect 34980 35649 35014 35683
rect 42441 35649 42475 35683
rect 49332 35649 49366 35683
rect 53012 35649 53046 35683
rect 54585 35649 54619 35683
rect 54852 35649 54886 35683
rect 6377 35581 6411 35615
rect 13369 35581 13403 35615
rect 27077 35581 27111 35615
rect 28917 35581 28951 35615
rect 34713 35581 34747 35615
rect 38025 35581 38059 35615
rect 39957 35581 39991 35615
rect 45661 35581 45695 35615
rect 49065 35581 49099 35615
rect 52745 35581 52779 35615
rect 5273 35445 5307 35479
rect 12909 35445 12943 35479
rect 14749 35445 14783 35479
rect 19533 35445 19567 35479
rect 28457 35445 28491 35479
rect 30297 35445 30331 35479
rect 43821 35445 43855 35479
rect 47041 35445 47075 35479
rect 50445 35445 50479 35479
rect 54125 35445 54159 35479
rect 55965 35445 55999 35479
rect 12909 35241 12943 35275
rect 17785 35241 17819 35275
rect 28457 35241 28491 35275
rect 31033 35241 31067 35275
rect 44465 35241 44499 35275
rect 47041 35241 47075 35275
rect 6929 35105 6963 35139
rect 11529 35105 11563 35139
rect 16405 35105 16439 35139
rect 19257 35105 19291 35139
rect 21097 35105 21131 35139
rect 29653 35105 29687 35139
rect 31493 35105 31527 35139
rect 37749 35105 37783 35139
rect 40417 35105 40451 35139
rect 45661 35105 45695 35139
rect 47685 35105 47719 35139
rect 55321 35105 55355 35139
rect 11796 35037 11830 35071
rect 14105 35037 14139 35071
rect 19524 35037 19558 35071
rect 25237 35037 25271 35071
rect 27077 35037 27111 35071
rect 29920 35037 29954 35071
rect 40684 35037 40718 35071
rect 43085 35037 43119 35071
rect 45928 35037 45962 35071
rect 50169 35037 50203 35071
rect 52009 35037 52043 35071
rect 55588 35037 55622 35071
rect 57161 35037 57195 35071
rect 7196 34969 7230 35003
rect 14372 34969 14406 35003
rect 16672 34969 16706 35003
rect 21364 34969 21398 35003
rect 25504 34969 25538 35003
rect 27344 34969 27378 35003
rect 31760 34969 31794 35003
rect 36001 34969 36035 35003
rect 43352 34969 43386 35003
rect 47952 34969 47986 35003
rect 50436 34969 50470 35003
rect 52276 34969 52310 35003
rect 57406 34969 57440 35003
rect 8309 34901 8343 34935
rect 15485 34901 15519 34935
rect 20637 34901 20671 34935
rect 22477 34901 22511 34935
rect 26617 34901 26651 34935
rect 32873 34901 32907 34935
rect 41797 34901 41831 34935
rect 49065 34901 49099 34935
rect 51549 34901 51583 34935
rect 53389 34901 53423 34935
rect 56701 34901 56735 34935
rect 58541 34901 58575 34935
rect 59461 34901 59495 34935
rect 10333 34697 10367 34731
rect 12909 34697 12943 34731
rect 14749 34697 14783 34731
rect 18245 34697 18279 34731
rect 23213 34697 23247 34731
rect 25145 34697 25179 34731
rect 28365 34697 28399 34731
rect 30205 34697 30239 34731
rect 36369 34697 36403 34731
rect 38669 34697 38703 34731
rect 40509 34697 40543 34731
rect 46857 34697 46891 34731
rect 48973 34697 49007 34731
rect 6745 34629 6779 34663
rect 13636 34629 13670 34663
rect 19524 34629 19558 34663
rect 29070 34629 29104 34663
rect 37534 34629 37568 34663
rect 39396 34629 39430 34663
rect 45744 34629 45778 34663
rect 49525 34629 49559 34663
rect 54830 34629 54864 34663
rect 8953 34561 8987 34595
rect 9220 34561 9254 34595
rect 11796 34561 11830 34595
rect 16865 34561 16899 34595
rect 17132 34561 17166 34595
rect 21833 34561 21867 34595
rect 22100 34561 22134 34595
rect 24032 34561 24066 34595
rect 27252 34561 27286 34595
rect 28825 34561 28859 34595
rect 33149 34561 33183 34595
rect 33416 34561 33450 34595
rect 35256 34561 35290 34595
rect 37289 34561 37323 34595
rect 43637 34561 43671 34595
rect 43904 34561 43938 34595
rect 47860 34561 47894 34595
rect 53012 34561 53046 34595
rect 54585 34561 54619 34595
rect 11529 34493 11563 34527
rect 13369 34493 13403 34527
rect 19257 34493 19291 34527
rect 23765 34493 23799 34527
rect 26985 34493 27019 34527
rect 34989 34493 35023 34527
rect 39129 34493 39163 34527
rect 45477 34493 45511 34527
rect 47593 34493 47627 34527
rect 52745 34493 52779 34527
rect 8033 34425 8067 34459
rect 54125 34425 54159 34459
rect 20637 34357 20671 34391
rect 34529 34357 34563 34391
rect 45017 34357 45051 34391
rect 50813 34357 50847 34391
rect 55965 34357 55999 34391
rect 10333 34153 10367 34187
rect 15485 34153 15519 34187
rect 18521 34153 18555 34187
rect 22385 34153 22419 34187
rect 27629 34153 27663 34187
rect 30941 34153 30975 34187
rect 36093 34153 36127 34187
rect 51549 34153 51583 34187
rect 53389 34153 53423 34187
rect 56701 34153 56735 34187
rect 8953 34017 8987 34051
rect 17141 34017 17175 34051
rect 26249 34017 26283 34051
rect 29561 34017 29595 34051
rect 39865 34017 39899 34051
rect 57161 34017 57195 34051
rect 4905 33949 4939 33983
rect 6745 33949 6779 33983
rect 10793 33949 10827 33983
rect 14105 33949 14139 33983
rect 14372 33949 14406 33983
rect 19257 33949 19291 33983
rect 19524 33949 19558 33983
rect 24409 33949 24443 33983
rect 29828 33949 29862 33983
rect 31677 33949 31711 33983
rect 34713 33949 34747 33983
rect 34969 33949 35003 33983
rect 37933 33949 37967 33983
rect 38200 33949 38234 33983
rect 42533 33949 42567 33983
rect 45017 33949 45051 33983
rect 46857 33949 46891 33983
rect 50169 33949 50203 33983
rect 52009 33949 52043 33983
rect 52265 33949 52299 33983
rect 55321 33949 55355 33983
rect 55588 33949 55622 33983
rect 5172 33881 5206 33915
rect 7012 33881 7046 33915
rect 9220 33881 9254 33915
rect 11060 33881 11094 33915
rect 17408 33881 17442 33915
rect 21097 33881 21131 33915
rect 24676 33881 24710 33915
rect 26494 33881 26528 33915
rect 31944 33881 31978 33915
rect 40110 33881 40144 33915
rect 42800 33881 42834 33915
rect 45284 33881 45318 33915
rect 47124 33881 47158 33915
rect 50436 33881 50470 33915
rect 57428 33881 57462 33915
rect 6285 33813 6319 33847
rect 8125 33813 8159 33847
rect 12173 33813 12207 33847
rect 20637 33813 20671 33847
rect 25789 33813 25823 33847
rect 33057 33813 33091 33847
rect 39313 33813 39347 33847
rect 41245 33813 41279 33847
rect 43913 33813 43947 33847
rect 46397 33813 46431 33847
rect 48237 33813 48271 33847
rect 58541 33813 58575 33847
rect 7757 33609 7791 33643
rect 9597 33609 9631 33643
rect 18429 33609 18463 33643
rect 25053 33609 25087 33643
rect 28365 33609 28399 33643
rect 33517 33609 33551 33643
rect 35357 33609 35391 33643
rect 39681 33609 39715 33643
rect 43821 33609 43855 33643
rect 48973 33609 49007 33643
rect 50813 33609 50847 33643
rect 54125 33609 54159 33643
rect 6622 33541 6656 33575
rect 8484 33541 8518 33575
rect 11897 33541 11931 33575
rect 19524 33541 19558 33575
rect 23940 33541 23974 33575
rect 27230 33541 27264 33575
rect 30104 33541 30138 33575
rect 38568 33541 38602 33575
rect 40141 33541 40175 33575
rect 44526 33541 44560 33575
rect 47860 33541 47894 33575
rect 49700 33541 49734 33575
rect 53012 33541 53046 33575
rect 54769 33541 54803 33575
rect 56517 33541 56551 33575
rect 4344 33473 4378 33507
rect 6377 33473 6411 33507
rect 8217 33473 8251 33507
rect 14372 33473 14406 33507
rect 17049 33473 17083 33507
rect 17316 33473 17350 33507
rect 21833 33473 21867 33507
rect 22100 33473 22134 33507
rect 23673 33473 23707 33507
rect 29837 33473 29871 33507
rect 32393 33473 32427 33507
rect 34233 33473 34267 33507
rect 42708 33473 42742 33507
rect 49433 33473 49467 33507
rect 4077 33405 4111 33439
rect 14105 33405 14139 33439
rect 19257 33405 19291 33439
rect 26985 33405 27019 33439
rect 32137 33405 32171 33439
rect 33977 33405 34011 33439
rect 38301 33405 38335 33439
rect 42441 33405 42475 33439
rect 44281 33405 44315 33439
rect 47593 33405 47627 33439
rect 52745 33405 52779 33439
rect 20637 33337 20671 33371
rect 5457 33269 5491 33303
rect 13185 33269 13219 33303
rect 15485 33269 15519 33303
rect 23213 33269 23247 33303
rect 31217 33269 31251 33303
rect 41429 33269 41463 33303
rect 45661 33269 45695 33303
rect 5181 33065 5215 33099
rect 7021 33065 7055 33099
rect 10333 33065 10367 33099
rect 12173 33065 12207 33099
rect 21005 33065 21039 33099
rect 22845 33065 22879 33099
rect 25789 33065 25823 33099
rect 36185 33065 36219 33099
rect 46397 33065 46431 33099
rect 52285 33065 52319 33099
rect 56701 33065 56735 33099
rect 58541 33065 58575 33099
rect 8953 32929 8987 32963
rect 14841 32929 14875 32963
rect 16681 32929 16715 32963
rect 29929 32929 29963 32963
rect 40325 32929 40359 32963
rect 42165 32929 42199 32963
rect 53389 32929 53423 32963
rect 57161 32929 57195 32963
rect 3801 32861 3835 32895
rect 5641 32861 5675 32895
rect 10793 32861 10827 32895
rect 11060 32861 11094 32895
rect 19625 32861 19659 32895
rect 19892 32861 19926 32895
rect 21465 32861 21499 32895
rect 21732 32861 21766 32895
rect 24409 32861 24443 32895
rect 24676 32861 24710 32895
rect 26985 32861 27019 32895
rect 30196 32861 30230 32895
rect 31953 32861 31987 32895
rect 32220 32861 32254 32895
rect 34805 32861 34839 32895
rect 36645 32861 36679 32895
rect 40592 32861 40626 32895
rect 45017 32861 45051 32895
rect 45284 32861 45318 32895
rect 46857 32861 46891 32895
rect 50905 32861 50939 32895
rect 51172 32861 51206 32895
rect 55321 32861 55355 32895
rect 55588 32861 55622 32895
rect 59461 32861 59495 32895
rect 4068 32793 4102 32827
rect 5908 32793 5942 32827
rect 9220 32793 9254 32827
rect 15108 32793 15142 32827
rect 16948 32793 16982 32827
rect 27252 32793 27286 32827
rect 35050 32793 35084 32827
rect 36912 32793 36946 32827
rect 42410 32793 42444 32827
rect 47102 32793 47136 32827
rect 53656 32793 53690 32827
rect 57428 32793 57462 32827
rect 16221 32725 16255 32759
rect 18061 32725 18095 32759
rect 28365 32725 28399 32759
rect 31309 32725 31343 32759
rect 33333 32725 33367 32759
rect 38025 32725 38059 32759
rect 41705 32725 41739 32759
rect 43545 32725 43579 32759
rect 48237 32725 48271 32759
rect 54769 32725 54803 32759
rect 4721 32521 4755 32555
rect 7757 32521 7791 32555
rect 9597 32521 9631 32555
rect 19901 32521 19935 32555
rect 23949 32521 23983 32555
rect 25789 32521 25823 32555
rect 31493 32521 31527 32555
rect 38669 32521 38703 32555
rect 43821 32521 43855 32555
rect 45661 32521 45695 32555
rect 48973 32521 49007 32555
rect 57345 32521 57379 32555
rect 6644 32453 6678 32487
rect 8462 32453 8496 32487
rect 12532 32453 12566 32487
rect 18766 32453 18800 32487
rect 22814 32453 22848 32487
rect 30380 32453 30414 32487
rect 32404 32453 32438 32487
rect 40132 32453 40166 32487
rect 44548 32453 44582 32487
rect 47860 32453 47894 32487
rect 54392 32453 54426 32487
rect 3341 32385 3375 32419
rect 3608 32385 3642 32419
rect 6377 32385 6411 32419
rect 8217 32385 8251 32419
rect 14361 32385 14395 32419
rect 16681 32385 16715 32419
rect 16948 32385 16982 32419
rect 18521 32385 18555 32419
rect 22569 32385 22603 32419
rect 24409 32385 24443 32419
rect 24665 32385 24699 32419
rect 28172 32385 28206 32419
rect 30113 32385 30147 32419
rect 32137 32385 32171 32419
rect 34621 32385 34655 32419
rect 34888 32385 34922 32419
rect 37556 32385 37590 32419
rect 39865 32385 39899 32419
rect 42441 32385 42475 32419
rect 42708 32385 42742 32419
rect 44281 32385 44315 32419
rect 47593 32385 47627 32419
rect 51080 32385 51114 32419
rect 54125 32385 54159 32419
rect 55965 32385 55999 32419
rect 56232 32385 56266 32419
rect 12265 32317 12299 32351
rect 14105 32317 14139 32351
rect 27905 32317 27939 32351
rect 37289 32317 37323 32351
rect 50813 32317 50847 32351
rect 18061 32249 18095 32283
rect 13645 32181 13679 32215
rect 15485 32181 15519 32215
rect 29285 32181 29319 32215
rect 33517 32181 33551 32215
rect 36001 32181 36035 32215
rect 41245 32181 41279 32215
rect 52193 32181 52227 32215
rect 55505 32181 55539 32215
rect 5181 31977 5215 32011
rect 17325 31977 17359 32011
rect 27537 31977 27571 32011
rect 33517 31977 33551 32011
rect 39313 31977 39347 32011
rect 41797 31977 41831 32011
rect 43637 31977 43671 32011
rect 46397 31977 46431 32011
rect 54769 31977 54803 32011
rect 57897 31977 57931 32011
rect 11621 31909 11655 31943
rect 31585 31909 31619 31943
rect 10241 31841 10275 31875
rect 14105 31841 14139 31875
rect 19625 31841 19659 31875
rect 35909 31841 35943 31875
rect 37933 31841 37967 31875
rect 40417 31841 40451 31875
rect 42257 31841 42291 31875
rect 45017 31841 45051 31875
rect 48237 31841 48271 31875
rect 51549 31841 51583 31875
rect 53389 31841 53423 31875
rect 3801 31773 3835 31807
rect 4068 31773 4102 31807
rect 10508 31773 10542 31807
rect 12081 31773 12115 31807
rect 12337 31773 12371 31807
rect 14372 31773 14406 31807
rect 15945 31773 15979 31807
rect 19892 31773 19926 31807
rect 22385 31773 22419 31807
rect 22652 31773 22686 31807
rect 26065 31773 26099 31807
rect 30205 31773 30239 31807
rect 30472 31773 30506 31807
rect 32137 31773 32171 31807
rect 32404 31773 32438 31807
rect 36176 31773 36210 31807
rect 38200 31773 38234 31807
rect 40684 31773 40718 31807
rect 42524 31773 42558 31807
rect 45284 31773 45318 31807
rect 48504 31773 48538 31807
rect 51816 31773 51850 31807
rect 53656 31773 53690 31807
rect 56517 31773 56551 31807
rect 56784 31773 56818 31807
rect 16190 31705 16224 31739
rect 13461 31637 13495 31671
rect 15485 31637 15519 31671
rect 21005 31637 21039 31671
rect 23765 31637 23799 31671
rect 37289 31637 37323 31671
rect 49617 31637 49651 31671
rect 52929 31637 52963 31671
rect 4261 31433 4295 31467
rect 14749 31433 14783 31467
rect 21281 31433 21315 31467
rect 31125 31433 31159 31467
rect 34621 31433 34655 31467
rect 36461 31433 36495 31467
rect 44005 31433 44039 31467
rect 50353 31433 50387 31467
rect 52193 31433 52227 31467
rect 29837 31365 29871 31399
rect 33508 31365 33542 31399
rect 35348 31365 35382 31399
rect 42892 31365 42926 31399
rect 49240 31365 49274 31399
rect 2881 31297 2915 31331
rect 3148 31297 3182 31331
rect 11529 31297 11563 31331
rect 11796 31297 11830 31331
rect 13636 31297 13670 31331
rect 18061 31297 18095 31331
rect 18328 31297 18362 31331
rect 20168 31297 20202 31331
rect 23213 31297 23247 31331
rect 23480 31297 23514 31331
rect 25320 31297 25354 31331
rect 28264 31297 28298 31331
rect 35081 31297 35115 31331
rect 38301 31297 38335 31331
rect 38568 31297 38602 31331
rect 40776 31297 40810 31331
rect 42625 31297 42659 31331
rect 45661 31297 45695 31331
rect 45928 31297 45962 31331
rect 48973 31297 49007 31331
rect 50813 31297 50847 31331
rect 51080 31297 51114 31331
rect 54484 31297 54518 31331
rect 13369 31229 13403 31263
rect 19901 31229 19935 31263
rect 25053 31229 25087 31263
rect 27997 31229 28031 31263
rect 33241 31229 33275 31263
rect 40509 31229 40543 31263
rect 54217 31229 54251 31263
rect 12909 31093 12943 31127
rect 19441 31093 19475 31127
rect 24593 31093 24627 31127
rect 26433 31093 26467 31127
rect 29377 31093 29411 31127
rect 39681 31093 39715 31127
rect 41889 31093 41923 31127
rect 47041 31093 47075 31127
rect 55597 31093 55631 31127
rect 13461 30889 13495 30923
rect 15485 30889 15519 30923
rect 17325 30889 17359 30923
rect 39313 30889 39347 30923
rect 52285 30889 52319 30923
rect 58541 30889 58575 30923
rect 12081 30753 12115 30787
rect 22477 30753 22511 30787
rect 43085 30753 43119 30787
rect 48237 30753 48271 30787
rect 3893 30685 3927 30719
rect 6469 30685 6503 30719
rect 9321 30685 9355 30719
rect 12348 30685 12382 30719
rect 14105 30685 14139 30719
rect 14372 30685 14406 30719
rect 15945 30685 15979 30719
rect 16212 30685 16246 30719
rect 20637 30685 20671 30719
rect 25789 30685 25823 30719
rect 27629 30685 27663 30719
rect 27896 30685 27930 30719
rect 31125 30685 31159 30719
rect 34713 30685 34747 30719
rect 34980 30685 35014 30719
rect 37933 30685 37967 30719
rect 38200 30685 38234 30719
rect 41245 30685 41279 30719
rect 46397 30685 46431 30719
rect 48504 30685 48538 30719
rect 50905 30685 50939 30719
rect 51172 30685 51206 30719
rect 52745 30685 52779 30719
rect 55321 30685 55355 30719
rect 55588 30685 55622 30719
rect 57161 30685 57195 30719
rect 4160 30617 4194 30651
rect 6736 30617 6770 30651
rect 9588 30617 9622 30651
rect 20904 30617 20938 30651
rect 22744 30617 22778 30651
rect 26056 30617 26090 30651
rect 31392 30617 31426 30651
rect 41512 30617 41546 30651
rect 43352 30617 43386 30651
rect 46664 30617 46698 30651
rect 53012 30617 53046 30651
rect 57406 30617 57440 30651
rect 5273 30549 5307 30583
rect 7849 30549 7883 30583
rect 10701 30549 10735 30583
rect 22017 30549 22051 30583
rect 23857 30549 23891 30583
rect 27169 30549 27203 30583
rect 29009 30549 29043 30583
rect 32505 30549 32539 30583
rect 36093 30549 36127 30583
rect 42625 30549 42659 30583
rect 44465 30549 44499 30583
rect 47777 30549 47811 30583
rect 49617 30549 49651 30583
rect 54125 30549 54159 30583
rect 56701 30549 56735 30583
rect 3985 30345 4019 30379
rect 5825 30345 5859 30379
rect 10977 30345 11011 30379
rect 19441 30345 19475 30379
rect 21281 30345 21315 30379
rect 24593 30345 24627 30379
rect 29745 30345 29779 30379
rect 33517 30345 33551 30379
rect 40969 30345 41003 30379
rect 52193 30345 52227 30379
rect 56701 30345 56735 30379
rect 14372 30277 14406 30311
rect 25320 30277 25354 30311
rect 28632 30277 28666 30311
rect 45928 30277 45962 30311
rect 51080 30277 51114 30311
rect 2605 30209 2639 30243
rect 2872 30209 2906 30243
rect 4445 30209 4479 30243
rect 4712 30209 4746 30243
rect 8024 30209 8058 30243
rect 9864 30209 9898 30243
rect 11529 30209 11563 30243
rect 11796 30209 11830 30243
rect 14105 30209 14139 30243
rect 18328 30209 18362 30243
rect 20168 30209 20202 30243
rect 23480 30209 23514 30243
rect 28365 30209 28399 30243
rect 30205 30209 30239 30243
rect 30472 30209 30506 30243
rect 32393 30209 32427 30243
rect 34253 30209 34287 30243
rect 37749 30209 37783 30243
rect 38016 30209 38050 30243
rect 39845 30209 39879 30243
rect 44088 30209 44122 30243
rect 49240 30209 49274 30243
rect 53012 30209 53046 30243
rect 55588 30209 55622 30243
rect 7757 30141 7791 30175
rect 9597 30141 9631 30175
rect 18061 30141 18095 30175
rect 19901 30141 19935 30175
rect 23213 30141 23247 30175
rect 25053 30141 25087 30175
rect 32137 30141 32171 30175
rect 39589 30141 39623 30175
rect 43821 30141 43855 30175
rect 45661 30141 45695 30175
rect 48973 30141 49007 30175
rect 50813 30141 50847 30175
rect 52745 30141 52779 30175
rect 55321 30141 55355 30175
rect 15485 30073 15519 30107
rect 26433 30073 26467 30107
rect 31585 30073 31619 30107
rect 39129 30073 39163 30107
rect 50353 30073 50387 30107
rect 9137 30005 9171 30039
rect 12909 30005 12943 30039
rect 35541 30005 35575 30039
rect 45201 30005 45235 30039
rect 47041 30005 47075 30039
rect 54125 30005 54159 30039
rect 13277 29801 13311 29835
rect 22017 29801 22051 29835
rect 27169 29801 27203 29835
rect 29009 29801 29043 29835
rect 31401 29801 31435 29835
rect 38853 29801 38887 29835
rect 42625 29801 42659 29835
rect 47133 29801 47167 29835
rect 53113 29801 53147 29835
rect 56701 29801 56735 29835
rect 11897 29665 11931 29699
rect 20637 29665 20671 29699
rect 30021 29665 30055 29699
rect 37473 29665 37507 29699
rect 41245 29665 41279 29699
rect 43085 29665 43119 29699
rect 45753 29665 45787 29699
rect 51733 29665 51767 29699
rect 55321 29665 55355 29699
rect 5181 29597 5215 29631
rect 5448 29597 5482 29631
rect 7021 29597 7055 29631
rect 7288 29597 7322 29631
rect 10057 29597 10091 29631
rect 14657 29597 14691 29631
rect 17049 29597 17083 29631
rect 20904 29597 20938 29631
rect 22477 29597 22511 29631
rect 22744 29597 22778 29631
rect 25789 29597 25823 29631
rect 27629 29597 27663 29631
rect 27896 29597 27930 29631
rect 30288 29597 30322 29631
rect 31861 29597 31895 29631
rect 34713 29597 34747 29631
rect 34980 29597 35014 29631
rect 41512 29597 41546 29631
rect 46020 29597 46054 29631
rect 55577 29597 55611 29631
rect 57161 29597 57195 29631
rect 57417 29597 57451 29631
rect 10324 29529 10358 29563
rect 12164 29529 12198 29563
rect 14924 29529 14958 29563
rect 17316 29529 17350 29563
rect 26056 29529 26090 29563
rect 32128 29529 32162 29563
rect 37740 29529 37774 29563
rect 43352 29529 43386 29563
rect 47593 29529 47627 29563
rect 52000 29529 52034 29563
rect 6561 29461 6595 29495
rect 8401 29461 8435 29495
rect 11437 29461 11471 29495
rect 16037 29461 16071 29495
rect 18429 29461 18463 29495
rect 23857 29461 23891 29495
rect 33241 29461 33275 29495
rect 36093 29461 36127 29495
rect 44465 29461 44499 29495
rect 48881 29461 48915 29495
rect 58541 29461 58575 29495
rect 59553 29461 59587 29495
rect 3985 29257 4019 29291
rect 5825 29257 5859 29291
rect 10977 29257 11011 29291
rect 16129 29257 16163 29291
rect 20821 29257 20855 29291
rect 25881 29257 25915 29291
rect 28641 29257 28675 29291
rect 31585 29257 31619 29291
rect 48973 29257 49007 29291
rect 56701 29257 56735 29291
rect 2872 29189 2906 29223
rect 6745 29189 6779 29223
rect 9864 29189 9898 29223
rect 13176 29189 13210 29223
rect 22744 29189 22778 29223
rect 24746 29189 24780 29223
rect 27506 29189 27540 29223
rect 30472 29189 30506 29223
rect 33140 29189 33174 29223
rect 34980 29189 35014 29223
rect 37832 29189 37866 29223
rect 45928 29189 45962 29223
rect 53113 29189 53147 29223
rect 55566 29189 55600 29223
rect 2605 29121 2639 29155
rect 4445 29121 4479 29155
rect 4712 29121 4746 29155
rect 12909 29121 12943 29155
rect 14749 29121 14783 29155
rect 15016 29121 15050 29155
rect 17684 29121 17718 29155
rect 19533 29121 19567 29155
rect 24501 29121 24535 29155
rect 27261 29121 27295 29155
rect 32873 29121 32907 29155
rect 37565 29121 37599 29155
rect 39681 29121 39715 29155
rect 39948 29121 39982 29155
rect 43821 29121 43855 29155
rect 44088 29121 44122 29155
rect 47593 29121 47627 29155
rect 47860 29121 47894 29155
rect 49700 29121 49734 29155
rect 55321 29121 55355 29155
rect 9597 29053 9631 29087
rect 17417 29053 17451 29087
rect 22477 29053 22511 29087
rect 30205 29053 30239 29087
rect 34713 29053 34747 29087
rect 45661 29053 45695 29087
rect 49433 29053 49467 29087
rect 8033 28985 8067 29019
rect 23857 28985 23891 29019
rect 41061 28985 41095 29019
rect 47041 28985 47075 29019
rect 50813 28985 50847 29019
rect 54401 28985 54435 29019
rect 14289 28917 14323 28951
rect 18797 28917 18831 28951
rect 34253 28917 34287 28951
rect 36093 28917 36127 28951
rect 38945 28917 38979 28951
rect 45201 28917 45235 28951
rect 6377 28713 6411 28747
rect 8401 28713 8435 28747
rect 11989 28713 12023 28747
rect 18705 28713 18739 28747
rect 20637 28713 20671 28747
rect 33793 28713 33827 28747
rect 38761 28713 38795 28747
rect 41521 28713 41555 28747
rect 44465 28713 44499 28747
rect 48973 28713 49007 28747
rect 54585 28713 54619 28747
rect 4997 28577 5031 28611
rect 37381 28577 37415 28611
rect 40141 28577 40175 28611
rect 43085 28577 43119 28611
rect 53205 28577 53239 28611
rect 5264 28509 5298 28543
rect 7021 28509 7055 28543
rect 10701 28509 10735 28543
rect 15485 28509 15519 28543
rect 17325 28509 17359 28543
rect 19257 28509 19291 28543
rect 19524 28509 19558 28543
rect 21833 28509 21867 28543
rect 25145 28509 25179 28543
rect 26985 28509 27019 28543
rect 29561 28509 29595 28543
rect 32413 28509 32447 28543
rect 32680 28509 32714 28543
rect 34805 28509 34839 28543
rect 35072 28509 35106 28543
rect 37648 28509 37682 28543
rect 43352 28509 43386 28543
rect 45753 28509 45787 28543
rect 46009 28509 46043 28543
rect 47593 28509 47627 28543
rect 50169 28509 50203 28543
rect 57069 28509 57103 28543
rect 7288 28441 7322 28475
rect 15752 28441 15786 28475
rect 17592 28441 17626 28475
rect 22100 28441 22134 28475
rect 25412 28441 25446 28475
rect 27252 28441 27286 28475
rect 29806 28441 29840 28475
rect 40408 28441 40442 28475
rect 47860 28441 47894 28475
rect 50436 28441 50470 28475
rect 53472 28441 53506 28475
rect 57314 28441 57348 28475
rect 16865 28373 16899 28407
rect 23213 28373 23247 28407
rect 26525 28373 26559 28407
rect 28365 28373 28399 28407
rect 30941 28373 30975 28407
rect 36185 28373 36219 28407
rect 47133 28373 47167 28407
rect 51549 28373 51583 28407
rect 58449 28373 58483 28407
rect 59461 28373 59495 28407
rect 9137 28169 9171 28203
rect 10977 28169 11011 28203
rect 25881 28169 25915 28203
rect 30205 28169 30239 28203
rect 39957 28169 39991 28203
rect 47041 28169 47075 28203
rect 49065 28169 49099 28203
rect 50905 28169 50939 28203
rect 54769 28169 54803 28203
rect 8024 28101 8058 28135
rect 9864 28101 9898 28135
rect 12992 28101 13026 28135
rect 15016 28101 15050 28135
rect 17316 28101 17350 28135
rect 19502 28101 19536 28135
rect 29070 28101 29104 28135
rect 35072 28101 35106 28135
rect 38669 28101 38703 28135
rect 44088 28101 44122 28135
rect 45928 28101 45962 28135
rect 49792 28101 49826 28135
rect 7757 28033 7791 28067
rect 12725 28033 12759 28067
rect 14749 28033 14783 28067
rect 19257 28033 19291 28067
rect 23020 28033 23054 28067
rect 24593 28033 24627 28067
rect 26985 28033 27019 28067
rect 27252 28033 27286 28067
rect 28825 28033 28859 28067
rect 32137 28033 32171 28067
rect 32404 28033 32438 28067
rect 43821 28033 43855 28067
rect 45661 28033 45695 28067
rect 47685 28033 47719 28067
rect 47952 28033 47986 28067
rect 53389 28033 53423 28067
rect 53656 28033 53690 28067
rect 55965 28033 55999 28067
rect 56232 28033 56266 28067
rect 9597 27965 9631 27999
rect 17049 27965 17083 27999
rect 22753 27965 22787 27999
rect 34805 27965 34839 27999
rect 49525 27965 49559 27999
rect 28365 27897 28399 27931
rect 45201 27897 45235 27931
rect 14105 27829 14139 27863
rect 16129 27829 16163 27863
rect 18429 27829 18463 27863
rect 20637 27829 20671 27863
rect 24133 27829 24167 27863
rect 33517 27829 33551 27863
rect 36185 27829 36219 27863
rect 57345 27829 57379 27863
rect 8217 27557 8251 27591
rect 13553 27557 13587 27591
rect 16405 27557 16439 27591
rect 20637 27557 20671 27591
rect 28365 27557 28399 27591
rect 41889 27557 41923 27591
rect 44465 27557 44499 27591
rect 54769 27557 54803 27591
rect 19257 27489 19291 27523
rect 40509 27489 40543 27523
rect 43085 27489 43119 27523
rect 50169 27489 50203 27523
rect 6837 27421 6871 27455
rect 7104 27421 7138 27455
rect 12173 27421 12207 27455
rect 12440 27421 12474 27455
rect 15025 27421 15059 27455
rect 15292 27421 15326 27455
rect 16865 27421 16899 27455
rect 17132 27421 17166 27455
rect 19524 27421 19558 27455
rect 22477 27421 22511 27455
rect 22744 27421 22778 27455
rect 24409 27421 24443 27455
rect 26985 27421 27019 27455
rect 29561 27421 29595 27455
rect 31401 27421 31435 27455
rect 31657 27421 31691 27455
rect 34713 27421 34747 27455
rect 34980 27421 35014 27455
rect 37289 27421 37323 27455
rect 40776 27421 40810 27455
rect 43352 27421 43386 27455
rect 45017 27421 45051 27455
rect 46857 27421 46891 27455
rect 53389 27421 53423 27455
rect 56517 27421 56551 27455
rect 24676 27353 24710 27387
rect 27252 27353 27286 27387
rect 29828 27353 29862 27387
rect 37556 27353 37590 27387
rect 45284 27353 45318 27387
rect 47124 27353 47158 27387
rect 50436 27353 50470 27387
rect 53656 27353 53690 27387
rect 56784 27353 56818 27387
rect 18245 27285 18279 27319
rect 23857 27285 23891 27319
rect 25789 27285 25823 27319
rect 30941 27285 30975 27319
rect 32781 27285 32815 27319
rect 36093 27285 36127 27319
rect 38669 27285 38703 27319
rect 46397 27285 46431 27319
rect 48237 27285 48271 27319
rect 51549 27285 51583 27319
rect 57897 27285 57931 27319
rect 18061 27081 18095 27115
rect 23489 27081 23523 27115
rect 25329 27081 25363 27115
rect 45661 27081 45695 27115
rect 48973 27081 49007 27115
rect 50813 27081 50847 27115
rect 54769 27081 54803 27115
rect 57345 27081 57379 27115
rect 13553 27013 13587 27047
rect 16948 27013 16982 27047
rect 22376 27013 22410 27047
rect 32772 27013 32806 27047
rect 34980 27013 35014 27047
rect 42708 27013 42742 27047
rect 47860 27013 47894 27047
rect 49700 27013 49734 27047
rect 56232 27013 56266 27047
rect 7665 26945 7699 26979
rect 7932 26945 7966 26979
rect 11529 26945 11563 26979
rect 11796 26945 11830 26979
rect 19901 26945 19935 26979
rect 20168 26945 20202 26979
rect 24216 26945 24250 26979
rect 28733 26945 28767 26979
rect 32505 26945 32539 26979
rect 34713 26945 34747 26979
rect 37657 26945 37691 26979
rect 37924 26945 37958 26979
rect 39497 26945 39531 26979
rect 39764 26945 39798 26979
rect 42441 26945 42475 26979
rect 44281 26945 44315 26979
rect 44548 26945 44582 26979
rect 49433 26945 49467 26979
rect 53389 26945 53423 26979
rect 53656 26945 53690 26979
rect 55965 26945 55999 26979
rect 16681 26877 16715 26911
rect 22109 26877 22143 26911
rect 23949 26877 23983 26911
rect 47593 26877 47627 26911
rect 36093 26809 36127 26843
rect 9045 26741 9079 26775
rect 12909 26741 12943 26775
rect 15025 26741 15059 26775
rect 21281 26741 21315 26775
rect 30205 26741 30239 26775
rect 33885 26741 33919 26775
rect 39037 26741 39071 26775
rect 40877 26741 40911 26775
rect 43821 26741 43855 26775
rect 11713 26537 11747 26571
rect 13553 26537 13587 26571
rect 17325 26537 17359 26571
rect 23121 26537 23155 26571
rect 25789 26537 25823 26571
rect 29009 26537 29043 26571
rect 41245 26537 41279 26571
rect 43361 26537 43395 26571
rect 46397 26537 46431 26571
rect 48237 26537 48271 26571
rect 51549 26537 51583 26571
rect 54769 26537 54803 26571
rect 15485 26469 15519 26503
rect 30941 26469 30975 26503
rect 57805 26469 57839 26503
rect 6653 26401 6687 26435
rect 19901 26401 19935 26435
rect 46857 26401 46891 26435
rect 50169 26401 50203 26435
rect 6920 26333 6954 26367
rect 10333 26333 10367 26367
rect 12173 26333 12207 26367
rect 14105 26333 14139 26367
rect 15945 26333 15979 26367
rect 20168 26333 20202 26367
rect 21741 26333 21775 26367
rect 22008 26333 22042 26367
rect 24409 26333 24443 26367
rect 27629 26333 27663 26367
rect 27896 26333 27930 26367
rect 29561 26333 29595 26367
rect 31401 26333 31435 26367
rect 31668 26333 31702 26367
rect 34713 26333 34747 26367
rect 36553 26333 36587 26367
rect 39865 26333 39899 26367
rect 42073 26333 42107 26367
rect 45017 26333 45051 26367
rect 50436 26333 50470 26367
rect 53389 26333 53423 26367
rect 56517 26333 56551 26367
rect 10600 26265 10634 26299
rect 12440 26265 12474 26299
rect 14372 26265 14406 26299
rect 16212 26265 16246 26299
rect 24676 26265 24710 26299
rect 29828 26265 29862 26299
rect 34958 26265 34992 26299
rect 36798 26265 36832 26299
rect 40132 26265 40166 26299
rect 45284 26265 45318 26299
rect 47124 26265 47158 26299
rect 53656 26265 53690 26299
rect 8033 26197 8067 26231
rect 21281 26197 21315 26231
rect 32781 26197 32815 26231
rect 36093 26197 36127 26231
rect 37933 26197 37967 26231
rect 8493 25993 8527 26027
rect 13553 25993 13587 26027
rect 18061 25993 18095 26027
rect 25513 25993 25547 26027
rect 31401 25993 31435 26027
rect 38669 25993 38703 26027
rect 57345 25993 57379 26027
rect 7380 25925 7414 25959
rect 9198 25925 9232 25959
rect 14258 25925 14292 25959
rect 16948 25925 16982 25959
rect 35440 25925 35474 25959
rect 39396 25925 39430 25959
rect 44548 25925 44582 25959
rect 50436 25925 50470 25959
rect 54392 25925 54426 25959
rect 4712 25857 4746 25891
rect 7113 25857 7147 25891
rect 12440 25857 12474 25891
rect 16681 25857 16715 25891
rect 18613 25857 18647 25891
rect 22100 25857 22134 25891
rect 24133 25857 24167 25891
rect 24400 25857 24434 25891
rect 26985 25857 27019 25891
rect 27252 25857 27286 25891
rect 30021 25857 30055 25891
rect 30288 25857 30322 25891
rect 32965 25857 32999 25891
rect 37556 25857 37590 25891
rect 39129 25857 39163 25891
rect 42708 25857 42742 25891
rect 44281 25857 44315 25891
rect 47961 25857 47995 25891
rect 50169 25857 50203 25891
rect 56232 25857 56266 25891
rect 4445 25789 4479 25823
rect 8953 25789 8987 25823
rect 12173 25789 12207 25823
rect 14013 25789 14047 25823
rect 20361 25789 20395 25823
rect 21833 25789 21867 25823
rect 35173 25789 35207 25823
rect 37289 25789 37323 25823
rect 42441 25789 42475 25823
rect 54125 25789 54159 25823
rect 55965 25789 55999 25823
rect 5825 25653 5859 25687
rect 10333 25653 10367 25687
rect 15393 25653 15427 25687
rect 23213 25653 23247 25687
rect 28365 25653 28399 25687
rect 34253 25653 34287 25687
rect 36553 25653 36587 25687
rect 40509 25653 40543 25687
rect 43821 25653 43855 25687
rect 45661 25653 45695 25687
rect 49433 25653 49467 25687
rect 51549 25653 51583 25687
rect 55505 25653 55539 25687
rect 13553 25449 13587 25483
rect 16497 25449 16531 25483
rect 23121 25449 23155 25483
rect 30941 25449 30975 25483
rect 32781 25449 32815 25483
rect 43085 25449 43119 25483
rect 46397 25449 46431 25483
rect 48237 25449 48271 25483
rect 54769 25449 54803 25483
rect 58173 25449 58207 25483
rect 12173 25313 12207 25347
rect 15117 25313 15151 25347
rect 19901 25313 19935 25347
rect 29561 25313 29595 25347
rect 36553 25313 36587 25347
rect 45017 25313 45051 25347
rect 56793 25313 56827 25347
rect 4537 25245 4571 25279
rect 6377 25245 6411 25279
rect 8953 25245 8987 25279
rect 9220 25245 9254 25279
rect 15384 25245 15418 25279
rect 17325 25245 17359 25279
rect 20168 25245 20202 25279
rect 21741 25245 21775 25279
rect 24409 25245 24443 25279
rect 26249 25245 26283 25279
rect 31401 25245 31435 25279
rect 31668 25245 31702 25279
rect 34713 25245 34747 25279
rect 36820 25245 36854 25279
rect 39865 25245 39899 25279
rect 40132 25245 40166 25279
rect 41705 25245 41739 25279
rect 41961 25245 41995 25279
rect 45284 25245 45318 25279
rect 46857 25245 46891 25279
rect 47113 25245 47147 25279
rect 50169 25245 50203 25279
rect 50436 25245 50470 25279
rect 53389 25245 53423 25279
rect 4804 25177 4838 25211
rect 6622 25177 6656 25211
rect 12440 25177 12474 25211
rect 17592 25177 17626 25211
rect 22008 25177 22042 25211
rect 24676 25177 24710 25211
rect 26494 25177 26528 25211
rect 29828 25177 29862 25211
rect 34980 25177 35014 25211
rect 53656 25177 53690 25211
rect 57060 25177 57094 25211
rect 5917 25109 5951 25143
rect 7757 25109 7791 25143
rect 10333 25109 10367 25143
rect 18705 25109 18739 25143
rect 21281 25109 21315 25143
rect 25789 25109 25823 25143
rect 27629 25109 27663 25143
rect 36093 25109 36127 25143
rect 37933 25109 37967 25143
rect 41245 25109 41279 25143
rect 51549 25109 51583 25143
rect 5181 24905 5215 24939
rect 13553 24905 13587 24939
rect 23213 24905 23247 24939
rect 25513 24905 25547 24939
rect 30205 24905 30239 24939
rect 38669 24905 38703 24939
rect 57345 24905 57379 24939
rect 37556 24837 37590 24871
rect 2228 24769 2262 24803
rect 3801 24769 3835 24803
rect 4068 24769 4102 24803
rect 6377 24769 6411 24803
rect 6644 24769 6678 24803
rect 9045 24769 9079 24803
rect 9312 24769 9346 24803
rect 12173 24769 12207 24803
rect 12440 24769 12474 24803
rect 14749 24769 14783 24803
rect 15016 24769 15050 24803
rect 17592 24769 17626 24803
rect 19809 24769 19843 24803
rect 20076 24769 20110 24803
rect 21833 24769 21867 24803
rect 22100 24769 22134 24803
rect 24400 24769 24434 24803
rect 27252 24769 27286 24803
rect 28825 24769 28859 24803
rect 29092 24769 29126 24803
rect 32137 24769 32171 24803
rect 32404 24769 32438 24803
rect 34233 24769 34267 24803
rect 37289 24769 37323 24803
rect 39385 24769 39419 24803
rect 43433 24769 43467 24803
rect 45273 24769 45307 24803
rect 47593 24769 47627 24803
rect 47860 24769 47894 24803
rect 49433 24769 49467 24803
rect 49700 24769 49734 24803
rect 54392 24769 54426 24803
rect 55965 24769 55999 24803
rect 56232 24769 56266 24803
rect 1961 24701 1995 24735
rect 17325 24701 17359 24735
rect 24133 24701 24167 24735
rect 26985 24701 27019 24735
rect 33977 24701 34011 24735
rect 39129 24701 39163 24735
rect 43177 24701 43211 24735
rect 45017 24701 45051 24735
rect 54125 24701 54159 24735
rect 33517 24633 33551 24667
rect 40509 24633 40543 24667
rect 44557 24633 44591 24667
rect 46397 24633 46431 24667
rect 3341 24565 3375 24599
rect 7757 24565 7791 24599
rect 10425 24565 10459 24599
rect 16129 24565 16163 24599
rect 18705 24565 18739 24599
rect 21189 24565 21223 24599
rect 28365 24565 28399 24599
rect 35357 24565 35391 24599
rect 48973 24565 49007 24599
rect 50813 24565 50847 24599
rect 55505 24565 55539 24599
rect 6561 24361 6595 24395
rect 13461 24361 13495 24395
rect 25789 24361 25823 24395
rect 30941 24361 30975 24395
rect 32781 24361 32815 24395
rect 37933 24361 37967 24395
rect 41245 24361 41279 24395
rect 43085 24361 43119 24395
rect 48973 24361 49007 24395
rect 56701 24361 56735 24395
rect 1869 24225 1903 24259
rect 15485 24225 15519 24259
rect 31401 24225 31435 24259
rect 34713 24225 34747 24259
rect 41705 24225 41739 24259
rect 45017 24225 45051 24259
rect 53113 24225 53147 24259
rect 55321 24225 55355 24259
rect 2136 24157 2170 24191
rect 9321 24157 9355 24191
rect 9588 24157 9622 24191
rect 11621 24157 11655 24191
rect 12081 24157 12115 24191
rect 15752 24157 15786 24191
rect 17325 24157 17359 24191
rect 17592 24157 17626 24191
rect 19441 24157 19475 24191
rect 19708 24157 19742 24191
rect 21281 24157 21315 24191
rect 24409 24157 24443 24191
rect 24665 24157 24699 24191
rect 26249 24157 26283 24191
rect 26516 24157 26550 24191
rect 29561 24157 29595 24191
rect 34980 24157 35014 24191
rect 36553 24157 36587 24191
rect 36820 24157 36854 24191
rect 39865 24157 39899 24191
rect 40132 24157 40166 24191
rect 41972 24157 42006 24191
rect 47593 24157 47627 24191
rect 49617 24157 49651 24191
rect 50169 24157 50203 24191
rect 55588 24157 55622 24191
rect 57161 24157 57195 24191
rect 59553 24361 59587 24395
rect 5273 24089 5307 24123
rect 12348 24089 12382 24123
rect 21548 24089 21582 24123
rect 29828 24089 29862 24123
rect 31646 24089 31680 24123
rect 45284 24089 45318 24123
rect 47860 24089 47894 24123
rect 50436 24089 50470 24123
rect 53380 24089 53414 24123
rect 57406 24089 57440 24123
rect 59461 24089 59495 24123
rect 3249 24021 3283 24055
rect 10701 24021 10735 24055
rect 11437 24021 11471 24055
rect 16865 24021 16899 24055
rect 18705 24021 18739 24055
rect 20821 24021 20855 24055
rect 22661 24021 22695 24055
rect 27629 24021 27663 24055
rect 36093 24021 36127 24055
rect 46397 24021 46431 24055
rect 49433 24021 49467 24055
rect 51549 24021 51583 24055
rect 54493 24021 54527 24055
rect 58541 24021 58575 24055
rect 5825 23817 5859 23851
rect 13277 23817 13311 23851
rect 20637 23817 20671 23851
rect 23213 23817 23247 23851
rect 25513 23817 25547 23851
rect 28365 23817 28399 23851
rect 33517 23817 33551 23851
rect 35357 23817 35391 23851
rect 41889 23817 41923 23851
rect 48973 23817 49007 23851
rect 50813 23817 50847 23851
rect 54769 23817 54803 23851
rect 57345 23817 57379 23851
rect 2596 23749 2630 23783
rect 9680 23749 9714 23783
rect 17684 23749 17718 23783
rect 19524 23749 19558 23783
rect 22100 23749 22134 23783
rect 27252 23749 27286 23783
rect 29092 23749 29126 23783
rect 32404 23749 32438 23783
rect 34244 23749 34278 23783
rect 45928 23749 45962 23783
rect 49700 23749 49734 23783
rect 53656 23749 53690 23783
rect 56232 23749 56266 23783
rect 2329 23681 2363 23715
rect 4712 23681 4746 23715
rect 7840 23681 7874 23715
rect 12164 23681 12198 23715
rect 15016 23681 15050 23715
rect 19257 23681 19291 23715
rect 21833 23681 21867 23715
rect 24400 23681 24434 23715
rect 32137 23681 32171 23715
rect 38844 23681 38878 23715
rect 40776 23681 40810 23715
rect 44088 23681 44122 23715
rect 47593 23681 47627 23715
rect 47860 23681 47894 23715
rect 49433 23681 49467 23715
rect 53389 23681 53423 23715
rect 55965 23681 55999 23715
rect 4445 23613 4479 23647
rect 7573 23613 7607 23647
rect 9413 23613 9447 23647
rect 11897 23613 11931 23647
rect 14749 23613 14783 23647
rect 17417 23613 17451 23647
rect 24133 23613 24167 23647
rect 26985 23613 27019 23647
rect 28825 23613 28859 23647
rect 33977 23613 34011 23647
rect 38577 23613 38611 23647
rect 40509 23613 40543 23647
rect 43821 23613 43855 23647
rect 45661 23613 45695 23647
rect 3709 23477 3743 23511
rect 8953 23477 8987 23511
rect 10793 23477 10827 23511
rect 16129 23477 16163 23511
rect 18797 23477 18831 23511
rect 30205 23477 30239 23511
rect 39957 23477 39991 23511
rect 45201 23477 45235 23511
rect 47041 23477 47075 23511
rect 6561 23273 6595 23307
rect 8401 23273 8435 23307
rect 16865 23273 16899 23307
rect 18705 23273 18739 23307
rect 25789 23273 25823 23307
rect 27629 23273 27663 23307
rect 46949 23273 46983 23307
rect 49341 23273 49375 23307
rect 5181 23137 5215 23171
rect 13553 23137 13587 23171
rect 15485 23137 15519 23171
rect 17325 23137 17359 23171
rect 30941 23137 30975 23171
rect 47961 23137 47995 23171
rect 1869 23069 1903 23103
rect 2136 23069 2170 23103
rect 5448 23069 5482 23103
rect 7021 23069 7055 23103
rect 7288 23069 7322 23103
rect 9321 23069 9355 23103
rect 9588 23069 9622 23103
rect 15752 23069 15786 23103
rect 17592 23069 17626 23103
rect 19257 23069 19291 23103
rect 21097 23069 21131 23103
rect 24409 23069 24443 23103
rect 26249 23069 26283 23103
rect 26516 23069 26550 23103
rect 32781 23069 32815 23103
rect 35265 23069 35299 23103
rect 37657 23069 37691 23103
rect 40601 23069 40635 23103
rect 41245 23069 41279 23103
rect 43085 23069 43119 23103
rect 45569 23069 45603 23103
rect 45836 23069 45870 23103
rect 50169 23069 50203 23103
rect 50436 23069 50470 23103
rect 52009 23069 52043 23103
rect 57161 23069 57195 23103
rect 11805 23001 11839 23035
rect 19524 23001 19558 23035
rect 21364 23001 21398 23035
rect 24676 23001 24710 23035
rect 31208 23001 31242 23035
rect 33048 23001 33082 23035
rect 35532 23001 35566 23035
rect 37924 23001 37958 23035
rect 41512 23001 41546 23035
rect 43352 23001 43386 23035
rect 48228 23001 48262 23035
rect 52254 23001 52288 23035
rect 57428 23001 57462 23035
rect 3249 22933 3283 22967
rect 10701 22933 10735 22967
rect 20637 22933 20671 22967
rect 22477 22933 22511 22967
rect 32321 22933 32355 22967
rect 34161 22933 34195 22967
rect 36645 22933 36679 22967
rect 39037 22933 39071 22967
rect 40417 22933 40451 22967
rect 42625 22933 42659 22967
rect 44465 22933 44499 22967
rect 51549 22933 51583 22967
rect 53389 22933 53423 22967
rect 58541 22933 58575 22967
rect 10609 22729 10643 22763
rect 13093 22729 13127 22763
rect 23213 22729 23247 22763
rect 25145 22729 25179 22763
rect 30941 22729 30975 22763
rect 46213 22729 46247 22763
rect 49617 22729 49651 22763
rect 57253 22729 57287 22763
rect 2504 22661 2538 22695
rect 9496 22661 9530 22695
rect 22100 22661 22134 22695
rect 27353 22661 27387 22695
rect 29828 22661 29862 22695
rect 43260 22661 43294 22695
rect 50436 22661 50470 22695
rect 56140 22661 56174 22695
rect 2237 22593 2271 22627
rect 9229 22593 9263 22627
rect 11713 22593 11747 22627
rect 11980 22593 12014 22627
rect 14749 22593 14783 22627
rect 15016 22593 15050 22627
rect 18153 22593 18187 22627
rect 18420 22593 18454 22627
rect 21097 22593 21131 22627
rect 21833 22593 21867 22627
rect 23765 22593 23799 22627
rect 24032 22593 24066 22627
rect 33517 22593 33551 22627
rect 33784 22593 33818 22627
rect 35357 22593 35391 22627
rect 35624 22593 35658 22627
rect 38752 22593 38786 22627
rect 40325 22593 40359 22627
rect 40592 22593 40626 22627
rect 42993 22593 43027 22627
rect 45100 22593 45134 22627
rect 48237 22593 48271 22627
rect 48504 22593 48538 22627
rect 50169 22593 50203 22627
rect 53012 22593 53046 22627
rect 29561 22525 29595 22559
rect 38485 22525 38519 22559
rect 44833 22525 44867 22559
rect 52745 22525 52779 22559
rect 55873 22525 55907 22559
rect 3617 22389 3651 22423
rect 16129 22389 16163 22423
rect 19533 22389 19567 22423
rect 20913 22389 20947 22423
rect 28641 22389 28675 22423
rect 34897 22389 34931 22423
rect 36737 22389 36771 22423
rect 39865 22389 39899 22423
rect 41705 22389 41739 22423
rect 44373 22389 44407 22423
rect 51549 22389 51583 22423
rect 54125 22389 54159 22423
rect 20637 22185 20671 22219
rect 25789 22185 25823 22219
rect 32321 22185 32355 22219
rect 34161 22185 34195 22219
rect 37473 22185 37507 22219
rect 39313 22185 39347 22219
rect 42625 22185 42659 22219
rect 44465 22185 44499 22219
rect 52009 22185 52043 22219
rect 15761 22049 15795 22083
rect 30941 22049 30975 22083
rect 37933 22049 37967 22083
rect 1869 21981 1903 22015
rect 2136 21981 2170 22015
rect 3801 21981 3835 22015
rect 11621 21981 11655 22015
rect 16028 21981 16062 22015
rect 19257 21981 19291 22015
rect 21097 21981 21131 22015
rect 24409 21981 24443 22015
rect 27629 21981 27663 22015
rect 32781 21981 32815 22015
rect 36093 21981 36127 22015
rect 36360 21981 36394 22015
rect 38200 21981 38234 22015
rect 41245 21981 41279 22015
rect 43085 21981 43119 22015
rect 43352 21981 43386 22015
rect 46305 21981 46339 22015
rect 50629 21981 50663 22015
rect 50896 21981 50930 22015
rect 52469 21981 52503 22015
rect 52736 21981 52770 22015
rect 56149 21981 56183 22015
rect 4046 21913 4080 21947
rect 11888 21913 11922 21947
rect 19524 21913 19558 21947
rect 21364 21913 21398 21947
rect 24676 21913 24710 21947
rect 27896 21913 27930 21947
rect 31208 21913 31242 21947
rect 33048 21913 33082 21947
rect 41512 21913 41546 21947
rect 3249 21845 3283 21879
rect 5181 21845 5215 21879
rect 13001 21845 13035 21879
rect 17141 21845 17175 21879
rect 22477 21845 22511 21879
rect 29009 21845 29043 21879
rect 47593 21845 47627 21879
rect 53849 21845 53883 21879
rect 57437 21845 57471 21879
rect 3433 21641 3467 21675
rect 16129 21641 16163 21675
rect 23213 21641 23247 21675
rect 25145 21641 25179 21675
rect 29009 21641 29043 21675
rect 34897 21641 34931 21675
rect 36737 21641 36771 21675
rect 40049 21641 40083 21675
rect 41889 21641 41923 21675
rect 49709 21641 49743 21675
rect 51549 21641 51583 21675
rect 2320 21573 2354 21607
rect 4160 21573 4194 21607
rect 16926 21573 16960 21607
rect 22100 21573 22134 21607
rect 30472 21573 30506 21607
rect 33784 21573 33818 21607
rect 38936 21573 38970 21607
rect 40776 21573 40810 21607
rect 42809 21573 42843 21607
rect 48596 21573 48630 21607
rect 53472 21573 53506 21607
rect 2053 21505 2087 21539
rect 3893 21505 3927 21539
rect 7288 21505 7322 21539
rect 12265 21505 12299 21539
rect 12532 21505 12566 21539
rect 14749 21505 14783 21539
rect 15016 21505 15050 21539
rect 18521 21505 18555 21539
rect 18788 21505 18822 21539
rect 21833 21505 21867 21539
rect 24032 21505 24066 21539
rect 27896 21505 27930 21539
rect 30205 21505 30239 21539
rect 33517 21505 33551 21539
rect 35357 21505 35391 21539
rect 35624 21505 35658 21539
rect 38669 21505 38703 21539
rect 40509 21505 40543 21539
rect 45273 21505 45307 21539
rect 48329 21505 48363 21539
rect 50436 21505 50470 21539
rect 53205 21505 53239 21539
rect 55045 21505 55079 21539
rect 55312 21505 55346 21539
rect 7021 21437 7055 21471
rect 16681 21437 16715 21471
rect 23765 21437 23799 21471
rect 27629 21437 27663 21471
rect 45017 21437 45051 21471
rect 50169 21437 50203 21471
rect 5273 21301 5307 21335
rect 8401 21301 8435 21335
rect 13645 21301 13679 21335
rect 18061 21301 18095 21335
rect 19901 21301 19935 21335
rect 31585 21301 31619 21335
rect 44097 21301 44131 21335
rect 46397 21301 46431 21335
rect 54585 21301 54619 21335
rect 56425 21301 56459 21335
rect 5457 21097 5491 21131
rect 13277 21097 13311 21131
rect 16497 21097 16531 21131
rect 18429 21097 18463 21131
rect 20637 21097 20671 21131
rect 25789 21097 25823 21131
rect 28825 21097 28859 21131
rect 37565 21097 37599 21131
rect 41245 21097 41279 21131
rect 44097 21097 44131 21131
rect 51549 21097 51583 21131
rect 56701 21097 56735 21131
rect 58541 21097 58575 21131
rect 11897 20961 11931 20995
rect 15117 20961 15151 20995
rect 19257 20961 19291 20995
rect 30021 20961 30055 20995
rect 52009 20961 52043 20995
rect 6377 20893 6411 20927
rect 8953 20893 8987 20927
rect 12164 20893 12198 20927
rect 15384 20893 15418 20927
rect 19524 20893 19558 20927
rect 21097 20893 21131 20927
rect 24409 20893 24443 20927
rect 27445 20893 27479 20927
rect 30288 20893 30322 20927
rect 31861 20893 31895 20927
rect 36185 20893 36219 20927
rect 36452 20893 36486 20927
rect 39865 20893 39899 20927
rect 40132 20893 40166 20927
rect 42717 20893 42751 20927
rect 42984 20893 43018 20927
rect 45661 20893 45695 20927
rect 47501 20893 47535 20927
rect 50169 20893 50203 20927
rect 52276 20893 52310 20927
rect 55321 20893 55355 20927
rect 57161 20893 57195 20927
rect 4169 20825 4203 20859
rect 6644 20825 6678 20859
rect 9220 20825 9254 20859
rect 16957 20825 16991 20859
rect 21342 20825 21376 20859
rect 24676 20825 24710 20859
rect 27712 20825 27746 20859
rect 45928 20825 45962 20859
rect 47768 20825 47802 20859
rect 50436 20825 50470 20859
rect 55588 20825 55622 20859
rect 57428 20825 57462 20859
rect 7757 20757 7791 20791
rect 10333 20757 10367 20791
rect 22477 20757 22511 20791
rect 31401 20757 31435 20791
rect 33149 20757 33183 20791
rect 47041 20757 47075 20791
rect 48881 20757 48915 20791
rect 53389 20757 53423 20791
rect 3893 20553 3927 20587
rect 7757 20553 7791 20587
rect 9597 20553 9631 20587
rect 20913 20553 20947 20587
rect 23213 20553 23247 20587
rect 33885 20553 33919 20587
rect 43821 20553 43855 20587
rect 46765 20553 46799 20587
rect 51273 20553 51307 20587
rect 54125 20553 54159 20587
rect 55965 20553 55999 20587
rect 4598 20485 4632 20519
rect 11888 20485 11922 20519
rect 15016 20485 15050 20519
rect 22100 20485 22134 20519
rect 24768 20485 24802 20519
rect 32772 20485 32806 20519
rect 34989 20485 35023 20519
rect 49985 20485 50019 20519
rect 54830 20485 54864 20519
rect 2780 20417 2814 20451
rect 6633 20417 6667 20451
rect 8217 20417 8251 20451
rect 8473 20417 8507 20451
rect 14749 20417 14783 20451
rect 17960 20417 17994 20451
rect 19533 20417 19567 20451
rect 19800 20417 19834 20451
rect 21833 20417 21867 20451
rect 27620 20417 27654 20451
rect 30205 20417 30239 20451
rect 30472 20417 30506 20451
rect 37289 20417 37323 20451
rect 37556 20417 37590 20451
rect 40509 20417 40543 20451
rect 40776 20417 40810 20451
rect 42708 20417 42742 20451
rect 45652 20417 45686 20451
rect 47777 20417 47811 20451
rect 48044 20417 48078 20451
rect 53012 20417 53046 20451
rect 54585 20417 54619 20451
rect 2513 20349 2547 20383
rect 4353 20349 4387 20383
rect 6377 20349 6411 20383
rect 11621 20349 11655 20383
rect 17693 20349 17727 20383
rect 24501 20349 24535 20383
rect 27353 20349 27387 20383
rect 32505 20349 32539 20383
rect 42441 20349 42475 20383
rect 45385 20349 45419 20383
rect 52745 20349 52779 20383
rect 13001 20281 13035 20315
rect 5733 20213 5767 20247
rect 16129 20213 16163 20247
rect 19073 20213 19107 20247
rect 25881 20213 25915 20247
rect 28733 20213 28767 20247
rect 31585 20213 31619 20247
rect 36277 20213 36311 20247
rect 38669 20213 38703 20247
rect 41889 20213 41923 20247
rect 49157 20213 49191 20247
rect 16313 20009 16347 20043
rect 18705 20009 18739 20043
rect 20637 20009 20671 20043
rect 22753 20009 22787 20043
rect 25789 20009 25823 20043
rect 28549 20009 28583 20043
rect 32137 20009 32171 20043
rect 36277 20009 36311 20043
rect 43729 20009 43763 20043
rect 46581 20009 46615 20043
rect 48605 20009 48639 20043
rect 53389 20009 53423 20043
rect 56701 20009 56735 20043
rect 58541 20009 58575 20043
rect 14933 19873 14967 19907
rect 30757 19873 30791 19907
rect 32597 19873 32631 19907
rect 34897 19873 34931 19907
rect 40509 19873 40543 19907
rect 50169 19873 50203 19907
rect 52009 19873 52043 19907
rect 4353 19805 4387 19839
rect 4620 19805 4654 19839
rect 6653 19805 6687 19839
rect 8953 19805 8987 19839
rect 11529 19805 11563 19839
rect 15200 19805 15234 19839
rect 17325 19805 17359 19839
rect 19257 19805 19291 19839
rect 19513 19805 19547 19839
rect 24409 19805 24443 19839
rect 24676 19805 24710 19839
rect 27169 19805 27203 19839
rect 31024 19805 31058 19839
rect 32853 19805 32887 19839
rect 35164 19805 35198 19839
rect 37841 19805 37875 19839
rect 42349 19805 42383 19839
rect 45201 19805 45235 19839
rect 47225 19805 47259 19839
rect 47481 19805 47515 19839
rect 50425 19805 50459 19839
rect 52276 19805 52310 19839
rect 55321 19805 55355 19839
rect 55577 19805 55611 19839
rect 57161 19805 57195 19839
rect 57417 19805 57451 19839
rect 8217 19737 8251 19771
rect 9220 19737 9254 19771
rect 11796 19737 11830 19771
rect 17592 19737 17626 19771
rect 21465 19737 21499 19771
rect 27436 19737 27470 19771
rect 38108 19737 38142 19771
rect 40776 19737 40810 19771
rect 42616 19737 42650 19771
rect 45468 19737 45502 19771
rect 5733 19669 5767 19703
rect 10333 19669 10367 19703
rect 12909 19669 12943 19703
rect 33977 19669 34011 19703
rect 39221 19669 39255 19703
rect 41889 19669 41923 19703
rect 51549 19669 51583 19703
rect 9597 19465 9631 19499
rect 18705 19465 18739 19499
rect 21281 19465 21315 19499
rect 28365 19465 28399 19499
rect 31585 19465 31619 19499
rect 36553 19465 36587 19499
rect 43821 19465 43855 19499
rect 46581 19465 46615 19499
rect 48973 19465 49007 19499
rect 50813 19465 50847 19499
rect 1860 19397 1894 19431
rect 4344 19397 4378 19431
rect 6644 19397 6678 19431
rect 13614 19397 13648 19431
rect 22078 19397 22112 19431
rect 27252 19397 27286 19431
rect 32382 19397 32416 19431
rect 40776 19397 40810 19431
rect 47860 19397 47894 19431
rect 49700 19397 49734 19431
rect 54033 19397 54067 19431
rect 55781 19397 55815 19431
rect 1593 19329 1627 19363
rect 4077 19329 4111 19363
rect 8217 19329 8251 19363
rect 8484 19329 8518 19363
rect 11529 19329 11563 19363
rect 11796 19329 11830 19363
rect 13369 19329 13403 19363
rect 17325 19329 17359 19363
rect 17592 19329 17626 19363
rect 19901 19329 19935 19363
rect 20168 19329 20202 19363
rect 21833 19329 21867 19363
rect 23929 19329 23963 19363
rect 26985 19329 27019 19363
rect 30205 19329 30239 19363
rect 30472 19329 30506 19363
rect 35173 19329 35207 19363
rect 35440 19329 35474 19363
rect 38936 19329 38970 19363
rect 42441 19329 42475 19363
rect 42708 19329 42742 19363
rect 45468 19329 45502 19363
rect 47593 19329 47627 19363
rect 49433 19329 49467 19363
rect 6377 19261 6411 19295
rect 23673 19261 23707 19295
rect 32137 19261 32171 19295
rect 38669 19261 38703 19295
rect 40509 19261 40543 19295
rect 45201 19261 45235 19295
rect 5457 19193 5491 19227
rect 12909 19193 12943 19227
rect 41889 19193 41923 19227
rect 2973 19125 3007 19159
rect 7757 19125 7791 19159
rect 14749 19125 14783 19159
rect 23213 19125 23247 19159
rect 25053 19125 25087 19159
rect 33517 19125 33551 19159
rect 40049 19125 40083 19159
rect 10333 18921 10367 18955
rect 32505 18921 32539 18955
rect 41245 18921 41279 18955
rect 43729 18921 43763 18955
rect 46489 18921 46523 18955
rect 1593 18785 1627 18819
rect 39865 18785 39899 18819
rect 1860 18717 1894 18751
rect 6377 18717 6411 18751
rect 6644 18717 6678 18751
rect 8953 18717 8987 18751
rect 9220 18717 9254 18751
rect 11529 18717 11563 18751
rect 13277 18717 13311 18751
rect 14105 18717 14139 18751
rect 15945 18717 15979 18751
rect 20729 18717 20763 18751
rect 25697 18717 25731 18751
rect 31125 18717 31159 18751
rect 31392 18717 31426 18751
rect 36093 18717 36127 18751
rect 36360 18717 36394 18751
rect 37933 18717 37967 18751
rect 40132 18717 40166 18751
rect 42349 18717 42383 18751
rect 45109 18717 45143 18751
rect 51917 18717 51951 18751
rect 56701 18717 56735 18751
rect 14372 18649 14406 18683
rect 16190 18649 16224 18683
rect 20996 18649 21030 18683
rect 27445 18649 27479 18683
rect 38200 18649 38234 18683
rect 42616 18649 42650 18683
rect 45376 18649 45410 18683
rect 52184 18649 52218 18683
rect 56968 18649 57002 18683
rect 2973 18581 3007 18615
rect 7757 18581 7791 18615
rect 15485 18581 15519 18615
rect 17325 18581 17359 18615
rect 22109 18581 22143 18615
rect 37473 18581 37507 18615
rect 39313 18581 39347 18615
rect 53297 18581 53331 18615
rect 58081 18581 58115 18615
rect 3157 18377 3191 18411
rect 12909 18377 12943 18411
rect 14749 18377 14783 18411
rect 19441 18377 19475 18411
rect 21281 18377 21315 18411
rect 28917 18377 28951 18411
rect 31217 18377 31251 18411
rect 36737 18377 36771 18411
rect 39681 18377 39715 18411
rect 43821 18377 43855 18411
rect 46397 18377 46431 18411
rect 2044 18309 2078 18343
rect 3862 18309 3896 18343
rect 6644 18309 6678 18343
rect 13636 18309 13670 18343
rect 18328 18309 18362 18343
rect 22100 18309 22134 18343
rect 23940 18309 23974 18343
rect 27804 18309 27838 18343
rect 30104 18309 30138 18343
rect 33784 18309 33818 18343
rect 38568 18309 38602 18343
rect 40141 18309 40175 18343
rect 56232 18309 56266 18343
rect 1777 18241 1811 18275
rect 3617 18241 3651 18275
rect 6377 18241 6411 18275
rect 8217 18241 8251 18275
rect 8484 18241 8518 18275
rect 11529 18241 11563 18275
rect 11796 18241 11830 18275
rect 13369 18241 13403 18275
rect 20168 18241 20202 18275
rect 21833 18241 21867 18275
rect 23673 18241 23707 18275
rect 27537 18241 27571 18275
rect 29837 18241 29871 18275
rect 35357 18241 35391 18275
rect 35624 18241 35658 18275
rect 38301 18241 38335 18275
rect 41889 18241 41923 18275
rect 42441 18241 42475 18275
rect 42708 18241 42742 18275
rect 45017 18241 45051 18275
rect 45284 18241 45318 18275
rect 50721 18241 50755 18275
rect 50988 18241 51022 18275
rect 54208 18241 54242 18275
rect 55965 18241 55999 18275
rect 18061 18173 18095 18207
rect 19901 18173 19935 18207
rect 33517 18173 33551 18207
rect 53941 18173 53975 18207
rect 7757 18105 7791 18139
rect 23213 18105 23247 18139
rect 4997 18037 5031 18071
rect 9597 18037 9631 18071
rect 25053 18037 25087 18071
rect 34897 18037 34931 18071
rect 52101 18037 52135 18071
rect 55321 18037 55355 18071
rect 57345 18037 57379 18071
rect 22293 17833 22327 17867
rect 37473 17833 37507 17867
rect 39313 17833 39347 17867
rect 43545 17833 43579 17867
rect 46397 17833 46431 17867
rect 52653 17833 52687 17867
rect 3801 17697 3835 17731
rect 14105 17697 14139 17731
rect 30941 17697 30975 17731
rect 32781 17697 32815 17731
rect 37933 17697 37967 17731
rect 42165 17697 42199 17731
rect 45017 17697 45051 17731
rect 47685 17697 47719 17731
rect 51273 17697 51307 17731
rect 6285 17629 6319 17663
rect 8953 17629 8987 17663
rect 10793 17629 10827 17663
rect 14372 17629 14406 17663
rect 15945 17629 15979 17663
rect 20913 17629 20947 17663
rect 25145 17629 25179 17663
rect 25401 17629 25435 17663
rect 27629 17629 27663 17663
rect 36093 17629 36127 17663
rect 38200 17629 38234 17663
rect 53113 17629 53147 17663
rect 53380 17629 53414 17663
rect 56793 17629 56827 17663
rect 4046 17561 4080 17595
rect 6552 17561 6586 17595
rect 9220 17561 9254 17595
rect 11038 17561 11072 17595
rect 16190 17561 16224 17595
rect 21180 17561 21214 17595
rect 27896 17561 27930 17595
rect 31208 17561 31242 17595
rect 33048 17561 33082 17595
rect 36360 17561 36394 17595
rect 42432 17561 42466 17595
rect 45284 17561 45318 17595
rect 47952 17561 47986 17595
rect 51540 17561 51574 17595
rect 57060 17561 57094 17595
rect 5181 17493 5215 17527
rect 7665 17493 7699 17527
rect 10333 17493 10367 17527
rect 12173 17493 12207 17527
rect 15485 17493 15519 17527
rect 17325 17493 17359 17527
rect 26525 17493 26559 17527
rect 29009 17493 29043 17527
rect 32321 17493 32355 17527
rect 34161 17493 34195 17527
rect 49065 17493 49099 17527
rect 54493 17493 54527 17527
rect 58173 17493 58207 17527
rect 3893 17289 3927 17323
rect 7757 17289 7791 17323
rect 9597 17289 9631 17323
rect 12909 17289 12943 17323
rect 21281 17289 21315 17323
rect 23213 17289 23247 17323
rect 35357 17289 35391 17323
rect 38761 17289 38795 17323
rect 40601 17289 40635 17323
rect 43821 17289 43855 17323
rect 46397 17289 46431 17323
rect 52193 17289 52227 17323
rect 57345 17289 57379 17323
rect 2780 17221 2814 17255
rect 14372 17221 14406 17255
rect 20168 17221 20202 17255
rect 24676 17221 24710 17255
rect 30472 17221 30506 17255
rect 32382 17221 32416 17255
rect 37626 17221 37660 17255
rect 39466 17221 39500 17255
rect 54392 17221 54426 17255
rect 56232 17221 56266 17255
rect 2513 17153 2547 17187
rect 4353 17153 4387 17187
rect 4620 17153 4654 17187
rect 6377 17153 6411 17187
rect 6644 17153 6678 17187
rect 8217 17153 8251 17187
rect 8484 17153 8518 17187
rect 11529 17153 11563 17187
rect 11796 17153 11830 17187
rect 14105 17153 14139 17187
rect 17233 17153 17267 17187
rect 17500 17153 17534 17187
rect 19901 17153 19935 17187
rect 21833 17153 21867 17187
rect 22100 17153 22134 17187
rect 24409 17153 24443 17187
rect 28632 17153 28666 17187
rect 33977 17153 34011 17187
rect 34244 17153 34278 17187
rect 37381 17153 37415 17187
rect 39221 17153 39255 17187
rect 42708 17153 42742 17187
rect 45017 17153 45051 17187
rect 45284 17153 45318 17187
rect 48973 17153 49007 17187
rect 49240 17153 49274 17187
rect 51080 17153 51114 17187
rect 54125 17153 54159 17187
rect 55965 17153 55999 17187
rect 28365 17085 28399 17119
rect 30205 17085 30239 17119
rect 32137 17085 32171 17119
rect 42441 17085 42475 17119
rect 50813 17085 50847 17119
rect 29745 17017 29779 17051
rect 5733 16949 5767 16983
rect 15485 16949 15519 16983
rect 18613 16949 18647 16983
rect 25789 16949 25823 16983
rect 31585 16949 31619 16983
rect 33517 16949 33551 16983
rect 50353 16949 50387 16983
rect 55505 16949 55539 16983
rect 5181 16745 5215 16779
rect 7021 16745 7055 16779
rect 10333 16745 10367 16779
rect 12173 16745 12207 16779
rect 15485 16745 15519 16779
rect 18521 16745 18555 16779
rect 37473 16745 37507 16779
rect 43913 16745 43947 16779
rect 46397 16745 46431 16779
rect 48789 16745 48823 16779
rect 52929 16745 52963 16779
rect 8953 16609 8987 16643
rect 14105 16609 14139 16643
rect 24409 16609 24443 16643
rect 36093 16609 36127 16643
rect 37933 16609 37967 16643
rect 40693 16609 40727 16643
rect 42533 16609 42567 16643
rect 47409 16609 47443 16643
rect 53389 16609 53423 16643
rect 3801 16541 3835 16575
rect 4068 16541 4102 16575
rect 5641 16541 5675 16575
rect 9220 16541 9254 16575
rect 10793 16541 10827 16575
rect 11060 16541 11094 16575
rect 14372 16541 14406 16575
rect 17141 16541 17175 16575
rect 20913 16541 20947 16575
rect 24676 16541 24710 16575
rect 26249 16541 26283 16575
rect 31033 16541 31067 16575
rect 36360 16541 36394 16575
rect 45017 16541 45051 16575
rect 47676 16541 47710 16575
rect 51549 16541 51583 16575
rect 51816 16541 51850 16575
rect 56517 16541 56551 16575
rect 5908 16473 5942 16507
rect 17408 16473 17442 16507
rect 21180 16473 21214 16507
rect 26494 16473 26528 16507
rect 31300 16473 31334 16507
rect 38200 16473 38234 16507
rect 40960 16473 40994 16507
rect 42800 16473 42834 16507
rect 45284 16473 45318 16507
rect 53656 16473 53690 16507
rect 56784 16473 56818 16507
rect 22293 16405 22327 16439
rect 25789 16405 25823 16439
rect 27629 16405 27663 16439
rect 32413 16405 32447 16439
rect 39313 16405 39347 16439
rect 42073 16405 42107 16439
rect 54769 16405 54803 16439
rect 57897 16405 57931 16439
rect 7757 16201 7791 16235
rect 9597 16201 9631 16235
rect 20545 16201 20579 16235
rect 23213 16201 23247 16235
rect 31585 16201 31619 16235
rect 33517 16201 33551 16235
rect 43821 16201 43855 16235
rect 46397 16201 46431 16235
rect 51733 16201 51767 16235
rect 57345 16201 57379 16235
rect 3608 16133 3642 16167
rect 8484 16133 8518 16167
rect 14648 16133 14682 16167
rect 19432 16133 19466 16167
rect 22100 16133 22134 16167
rect 24676 16133 24710 16167
rect 30472 16133 30506 16167
rect 32404 16133 32438 16167
rect 34958 16133 34992 16167
rect 42686 16133 42720 16167
rect 47952 16133 47986 16167
rect 50620 16133 50654 16167
rect 54392 16133 54426 16167
rect 56232 16133 56266 16167
rect 1768 16065 1802 16099
rect 6644 16065 6678 16099
rect 8217 16065 8251 16099
rect 14381 16065 14415 16099
rect 17325 16065 17359 16099
rect 17592 16065 17626 16099
rect 19165 16065 19199 16099
rect 24409 16065 24443 16099
rect 27241 16065 27275 16099
rect 30205 16065 30239 16099
rect 32137 16065 32171 16099
rect 38108 16065 38142 16099
rect 40408 16065 40442 16099
rect 42441 16065 42475 16099
rect 45017 16065 45051 16099
rect 45284 16065 45318 16099
rect 50353 16065 50387 16099
rect 1501 15997 1535 16031
rect 3341 15997 3375 16031
rect 6377 15997 6411 16031
rect 21833 15997 21867 16031
rect 26985 15997 27019 16031
rect 34713 15997 34747 16031
rect 37841 15997 37875 16031
rect 40141 15997 40175 16031
rect 47685 15997 47719 16031
rect 54125 15997 54159 16031
rect 55965 15997 55999 16031
rect 4721 15929 4755 15963
rect 55505 15929 55539 15963
rect 2881 15861 2915 15895
rect 15761 15861 15795 15895
rect 18705 15861 18739 15895
rect 25789 15861 25823 15895
rect 28365 15861 28399 15895
rect 36093 15861 36127 15895
rect 39221 15861 39255 15895
rect 41521 15861 41555 15895
rect 49065 15861 49099 15895
rect 6929 15657 6963 15691
rect 18705 15657 18739 15691
rect 21189 15657 21223 15691
rect 23489 15657 23523 15691
rect 25789 15657 25823 15691
rect 39037 15657 39071 15691
rect 41245 15657 41279 15691
rect 43085 15657 43119 15691
rect 46397 15657 46431 15691
rect 57805 15657 57839 15691
rect 14381 15521 14415 15555
rect 22109 15521 22143 15555
rect 24409 15521 24443 15555
rect 39865 15521 39899 15555
rect 1869 15453 1903 15487
rect 2136 15453 2170 15487
rect 5549 15453 5583 15487
rect 10425 15453 10459 15487
rect 14648 15453 14682 15487
rect 17325 15453 17359 15487
rect 24676 15453 24710 15487
rect 26801 15453 26835 15487
rect 27068 15453 27102 15487
rect 30757 15453 30791 15487
rect 32781 15453 32815 15487
rect 34713 15453 34747 15487
rect 34980 15453 35014 15487
rect 37657 15453 37691 15487
rect 40121 15453 40155 15487
rect 41705 15453 41739 15487
rect 45017 15453 45051 15487
rect 47869 15453 47903 15487
rect 50169 15453 50203 15487
rect 52009 15453 52043 15487
rect 56425 15453 56459 15487
rect 5816 15385 5850 15419
rect 10692 15385 10726 15419
rect 17592 15385 17626 15419
rect 19901 15385 19935 15419
rect 22376 15385 22410 15419
rect 31024 15385 31058 15419
rect 33048 15385 33082 15419
rect 37924 15385 37958 15419
rect 41950 15385 41984 15419
rect 45284 15385 45318 15419
rect 50436 15385 50470 15419
rect 52276 15385 52310 15419
rect 56692 15385 56726 15419
rect 3249 15317 3283 15351
rect 11805 15317 11839 15351
rect 15761 15317 15795 15351
rect 28181 15317 28215 15351
rect 32137 15317 32171 15351
rect 34161 15317 34195 15351
rect 36093 15317 36127 15351
rect 49157 15317 49191 15351
rect 51549 15317 51583 15351
rect 53389 15317 53423 15351
rect 7941 15113 7975 15147
rect 18797 15113 18831 15147
rect 20637 15113 20671 15147
rect 26341 15113 26375 15147
rect 38945 15113 38979 15147
rect 40877 15113 40911 15147
rect 46397 15113 46431 15147
rect 57345 15113 57379 15147
rect 1952 15045 1986 15079
rect 12532 15045 12566 15079
rect 14556 15045 14590 15079
rect 23388 15045 23422 15079
rect 25228 15045 25262 15079
rect 27252 15045 27286 15079
rect 29092 15045 29126 15079
rect 34980 15045 35014 15079
rect 39742 15045 39776 15079
rect 47952 15045 47986 15079
rect 1685 14977 1719 15011
rect 6828 14977 6862 15011
rect 8493 14977 8527 15011
rect 8760 14977 8794 15011
rect 14289 14977 14323 15011
rect 17684 14977 17718 15011
rect 19257 14977 19291 15011
rect 19513 14977 19547 15011
rect 23121 14977 23155 15011
rect 24961 14977 24995 15011
rect 26985 14977 27019 15011
rect 33140 14977 33174 15011
rect 34713 14977 34747 15011
rect 37565 14977 37599 15011
rect 37832 14977 37866 15011
rect 39497 14977 39531 15011
rect 45017 14977 45051 15011
rect 45284 14977 45318 15011
rect 49781 14977 49815 15011
rect 52745 14977 52779 15011
rect 53012 14977 53046 15011
rect 56232 14977 56266 15011
rect 6561 14909 6595 14943
rect 12265 14909 12299 14943
rect 17417 14909 17451 14943
rect 28825 14909 28859 14943
rect 32873 14909 32907 14943
rect 47685 14909 47719 14943
rect 49525 14909 49559 14943
rect 55965 14909 55999 14943
rect 3065 14773 3099 14807
rect 9873 14773 9907 14807
rect 13645 14773 13679 14807
rect 15669 14773 15703 14807
rect 24501 14773 24535 14807
rect 28365 14773 28399 14807
rect 30205 14773 30239 14807
rect 34253 14773 34287 14807
rect 36093 14773 36127 14807
rect 49065 14773 49099 14807
rect 50905 14773 50939 14807
rect 54125 14773 54159 14807
rect 8125 14569 8159 14603
rect 18521 14569 18555 14603
rect 23673 14569 23707 14603
rect 31861 14569 31895 14603
rect 41245 14569 41279 14603
rect 46673 14569 46707 14603
rect 20453 14433 20487 14467
rect 34069 14433 34103 14467
rect 34897 14433 34931 14467
rect 39313 14433 39347 14467
rect 39865 14433 39899 14467
rect 45293 14433 45327 14467
rect 52009 14433 52043 14467
rect 1685 14365 1719 14399
rect 1952 14365 1986 14399
rect 6745 14365 6779 14399
rect 9873 14365 9907 14399
rect 12173 14365 12207 14399
rect 14105 14365 14139 14399
rect 14372 14365 14406 14399
rect 17141 14365 17175 14399
rect 22293 14365 22327 14399
rect 30481 14365 30515 14399
rect 30748 14365 30782 14399
rect 35164 14365 35198 14399
rect 40132 14365 40166 14399
rect 47593 14365 47627 14399
rect 47860 14365 47894 14399
rect 50169 14365 50203 14399
rect 52265 14365 52299 14399
rect 56701 14365 56735 14399
rect 4537 14297 4571 14331
rect 7012 14297 7046 14331
rect 12440 14297 12474 14331
rect 17408 14297 17442 14331
rect 20720 14297 20754 14331
rect 22560 14297 22594 14331
rect 25973 14297 26007 14331
rect 27537 14297 27571 14331
rect 32321 14297 32355 14331
rect 37565 14297 37599 14331
rect 45560 14297 45594 14331
rect 50414 14297 50448 14331
rect 56946 14297 56980 14331
rect 3065 14229 3099 14263
rect 5825 14229 5859 14263
rect 11161 14229 11195 14263
rect 13553 14229 13587 14263
rect 15485 14229 15519 14263
rect 21833 14229 21867 14263
rect 36277 14229 36311 14263
rect 48973 14229 49007 14263
rect 51549 14229 51583 14263
rect 53389 14229 53423 14263
rect 58081 14229 58115 14263
rect 7941 14025 7975 14059
rect 12909 14025 12943 14059
rect 18061 14025 18095 14059
rect 21281 14025 21315 14059
rect 23213 14025 23247 14059
rect 34161 14025 34195 14059
rect 38945 14025 38979 14059
rect 46121 14025 46155 14059
rect 49065 14025 49099 14059
rect 57345 14025 57379 14059
rect 1952 13957 1986 13991
rect 9864 13957 9898 13991
rect 14372 13957 14406 13991
rect 20168 13957 20202 13991
rect 22078 13957 22112 13991
rect 25320 13957 25354 13991
rect 27252 13957 27286 13991
rect 33048 13957 33082 13991
rect 35256 13957 35290 13991
rect 47952 13957 47986 13991
rect 50068 13957 50102 13991
rect 54861 13957 54895 13991
rect 56232 13957 56266 13991
rect 1685 13889 1719 13923
rect 6828 13889 6862 13923
rect 11796 13889 11830 13923
rect 14105 13889 14139 13923
rect 16681 13889 16715 13923
rect 16948 13889 16982 13923
rect 25053 13889 25087 13923
rect 26985 13889 27019 13923
rect 28825 13889 28859 13923
rect 29092 13889 29126 13923
rect 32781 13889 32815 13923
rect 34989 13889 35023 13923
rect 37565 13889 37599 13923
rect 37832 13889 37866 13923
rect 43157 13889 43191 13923
rect 44741 13889 44775 13923
rect 45008 13889 45042 13923
rect 49801 13889 49835 13923
rect 53113 13889 53147 13923
rect 6561 13821 6595 13855
rect 9597 13821 9631 13855
rect 11529 13821 11563 13855
rect 19901 13821 19935 13855
rect 21833 13821 21867 13855
rect 42901 13821 42935 13855
rect 47685 13821 47719 13855
rect 55965 13821 55999 13855
rect 3065 13685 3099 13719
rect 10977 13685 11011 13719
rect 15485 13685 15519 13719
rect 26433 13685 26467 13719
rect 28365 13685 28399 13719
rect 30205 13685 30239 13719
rect 36369 13685 36403 13719
rect 44281 13685 44315 13719
rect 51181 13685 51215 13719
rect 8217 13481 8251 13515
rect 12173 13481 12207 13515
rect 26709 13481 26743 13515
rect 36369 13481 36403 13515
rect 38945 13481 38979 13515
rect 42809 13481 42843 13515
rect 46397 13481 46431 13515
rect 49341 13481 49375 13515
rect 51549 13481 51583 13515
rect 53389 13481 53423 13515
rect 25329 13345 25363 13379
rect 27169 13345 27203 13379
rect 34989 13345 35023 13379
rect 37565 13345 37599 13379
rect 52009 13345 52043 13379
rect 1869 13277 1903 13311
rect 2136 13277 2170 13311
rect 4997 13277 5031 13311
rect 6837 13277 6871 13311
rect 8953 13277 8987 13311
rect 10793 13277 10827 13311
rect 11060 13277 11094 13311
rect 20729 13277 20763 13311
rect 25596 13277 25630 13311
rect 27436 13277 27470 13311
rect 30941 13277 30975 13311
rect 32781 13277 32815 13311
rect 35256 13277 35290 13311
rect 41429 13277 41463 13311
rect 45017 13277 45051 13311
rect 47961 13277 47995 13311
rect 48228 13277 48262 13311
rect 50169 13277 50203 13311
rect 50436 13277 50470 13311
rect 52276 13277 52310 13311
rect 56701 13277 56735 13311
rect 5264 13209 5298 13243
rect 7104 13209 7138 13243
rect 9220 13209 9254 13243
rect 15577 13209 15611 13243
rect 20996 13209 21030 13243
rect 31208 13209 31242 13243
rect 33048 13209 33082 13243
rect 37832 13209 37866 13243
rect 41696 13209 41730 13243
rect 45284 13209 45318 13243
rect 3249 13141 3283 13175
rect 6377 13141 6411 13175
rect 10333 13141 10367 13175
rect 16865 13141 16899 13175
rect 22109 13141 22143 13175
rect 28549 13141 28583 13175
rect 32321 13141 32355 13175
rect 34161 13141 34195 13175
rect 57989 13141 58023 13175
rect 3525 12937 3559 12971
rect 7757 12937 7791 12971
rect 10977 12937 11011 12971
rect 15209 12937 15243 12971
rect 21281 12937 21315 12971
rect 36093 12937 36127 12971
rect 38945 12937 38979 12971
rect 46765 12937 46799 12971
rect 51917 12937 51951 12971
rect 54861 12937 54895 12971
rect 2412 12869 2446 12903
rect 4230 12869 4264 12903
rect 9864 12869 9898 12903
rect 14096 12869 14130 12903
rect 20168 12869 20202 12903
rect 24032 12869 24066 12903
rect 27528 12869 27562 12903
rect 34958 12869 34992 12903
rect 44925 12869 44959 12903
rect 48964 12869 48998 12903
rect 53748 12869 53782 12903
rect 2145 12801 2179 12835
rect 6644 12801 6678 12835
rect 9597 12801 9631 12835
rect 16681 12801 16715 12835
rect 16948 12801 16982 12835
rect 19901 12801 19935 12835
rect 23765 12801 23799 12835
rect 27261 12801 27295 12835
rect 29357 12801 29391 12835
rect 32137 12801 32171 12835
rect 32404 12801 32438 12835
rect 37565 12801 37599 12835
rect 37832 12801 37866 12835
rect 43177 12801 43211 12835
rect 45385 12801 45419 12835
rect 45652 12801 45686 12835
rect 48697 12801 48731 12835
rect 50793 12801 50827 12835
rect 53481 12801 53515 12835
rect 56221 12801 56255 12835
rect 3985 12733 4019 12767
rect 6377 12733 6411 12767
rect 13829 12733 13863 12767
rect 29101 12733 29135 12767
rect 34713 12733 34747 12767
rect 50537 12733 50571 12767
rect 55965 12733 55999 12767
rect 5365 12597 5399 12631
rect 18061 12597 18095 12631
rect 25145 12597 25179 12631
rect 28641 12597 28675 12631
rect 30481 12597 30515 12631
rect 33517 12597 33551 12631
rect 50077 12597 50111 12631
rect 57345 12597 57379 12631
rect 15485 12393 15519 12427
rect 22293 12393 22327 12427
rect 28825 12393 28859 12427
rect 38945 12393 38979 12427
rect 43913 12393 43947 12427
rect 5641 12257 5675 12291
rect 9413 12257 9447 12291
rect 24409 12257 24443 12291
rect 37565 12257 37599 12291
rect 46397 12257 46431 12291
rect 48237 12257 48271 12291
rect 53021 12257 53055 12291
rect 57253 12257 57287 12291
rect 3801 12189 3835 12223
rect 9680 12189 9714 12223
rect 14105 12189 14139 12223
rect 14361 12189 14395 12223
rect 15945 12189 15979 12223
rect 20913 12189 20947 12223
rect 24676 12189 24710 12223
rect 27445 12189 27479 12223
rect 27712 12189 27746 12223
rect 29561 12189 29595 12223
rect 29828 12189 29862 12223
rect 31401 12189 31435 12223
rect 34713 12189 34747 12223
rect 40693 12189 40727 12223
rect 42533 12189 42567 12223
rect 51181 12189 51215 12223
rect 53288 12189 53322 12223
rect 55413 12189 55447 12223
rect 55680 12189 55714 12223
rect 57520 12189 57554 12223
rect 4068 12121 4102 12155
rect 5886 12121 5920 12155
rect 16212 12121 16246 12155
rect 21180 12121 21214 12155
rect 31646 12121 31680 12155
rect 34980 12121 35014 12155
rect 37832 12121 37866 12155
rect 40960 12121 40994 12155
rect 42778 12121 42812 12155
rect 46664 12121 46698 12155
rect 48504 12121 48538 12155
rect 51448 12121 51482 12155
rect 5181 12053 5215 12087
rect 7021 12053 7055 12087
rect 10793 12053 10827 12087
rect 17325 12053 17359 12087
rect 25789 12053 25823 12087
rect 30941 12053 30975 12087
rect 32781 12053 32815 12087
rect 36093 12053 36127 12087
rect 42073 12053 42107 12087
rect 47777 12053 47811 12087
rect 49617 12053 49651 12087
rect 52561 12053 52595 12087
rect 54401 12053 54435 12087
rect 56793 12053 56827 12087
rect 58633 12053 58667 12087
rect 4261 11849 4295 11883
rect 7757 11849 7791 11883
rect 13553 11849 13587 11883
rect 23213 11849 23247 11883
rect 29285 11849 29319 11883
rect 31125 11849 31159 11883
rect 33517 11849 33551 11883
rect 38853 11849 38887 11883
rect 41889 11849 41923 11883
rect 43821 11849 43855 11883
rect 45661 11849 45695 11883
rect 50353 11849 50387 11883
rect 55505 11849 55539 11883
rect 3148 11781 3182 11815
rect 6622 11781 6656 11815
rect 9680 11781 9714 11815
rect 14258 11781 14292 11815
rect 16948 11781 16982 11815
rect 22100 11781 22134 11815
rect 24400 11781 24434 11815
rect 28172 11781 28206 11815
rect 30012 11781 30046 11815
rect 42708 11781 42742 11815
rect 44548 11781 44582 11815
rect 54392 11781 54426 11815
rect 58449 11781 58483 11815
rect 2881 11713 2915 11747
rect 9413 11713 9447 11747
rect 12440 11713 12474 11747
rect 20168 11713 20202 11747
rect 21833 11713 21867 11747
rect 24133 11713 24167 11747
rect 27905 11713 27939 11747
rect 32137 11713 32171 11747
rect 32404 11713 32438 11747
rect 34244 11713 34278 11747
rect 37473 11713 37507 11747
rect 37740 11713 37774 11747
rect 40509 11713 40543 11747
rect 40776 11713 40810 11747
rect 42441 11713 42475 11747
rect 49240 11713 49274 11747
rect 50813 11713 50847 11747
rect 51080 11713 51114 11747
rect 55965 11713 55999 11747
rect 56232 11713 56266 11747
rect 58633 11713 58667 11747
rect 6377 11645 6411 11679
rect 12173 11645 12207 11679
rect 14013 11645 14047 11679
rect 16681 11645 16715 11679
rect 19901 11645 19935 11679
rect 29745 11645 29779 11679
rect 33977 11645 34011 11679
rect 44281 11645 44315 11679
rect 48973 11645 49007 11679
rect 54125 11645 54159 11679
rect 10793 11509 10827 11543
rect 15393 11509 15427 11543
rect 18061 11509 18095 11543
rect 21281 11509 21315 11543
rect 25513 11509 25547 11543
rect 35357 11509 35391 11543
rect 52193 11509 52227 11543
rect 57345 11509 57379 11543
rect 5825 11305 5859 11339
rect 11529 11305 11563 11339
rect 15485 11305 15519 11339
rect 17325 11305 17359 11339
rect 21281 11305 21315 11339
rect 23489 11305 23523 11339
rect 31953 11305 31987 11339
rect 33793 11305 33827 11339
rect 36093 11305 36127 11339
rect 38761 11305 38795 11339
rect 39865 11305 39899 11339
rect 41889 11305 41923 11339
rect 49617 11305 49651 11339
rect 52929 11305 52963 11339
rect 13553 11237 13587 11271
rect 12173 11169 12207 11203
rect 15945 11169 15979 11203
rect 40509 11169 40543 11203
rect 46397 11169 46431 11203
rect 53389 11169 53423 11203
rect 56885 11169 56919 11203
rect 4445 11101 4479 11135
rect 4712 11101 4746 11135
rect 9413 11101 9447 11135
rect 9680 11101 9714 11135
rect 11713 11101 11747 11135
rect 14105 11101 14139 11135
rect 16201 11101 16235 11135
rect 19901 11101 19935 11135
rect 22109 11101 22143 11135
rect 24409 11101 24443 11135
rect 24676 11101 24710 11135
rect 30573 11101 30607 11135
rect 30840 11101 30874 11135
rect 32413 11101 32447 11135
rect 32680 11101 32714 11135
rect 34713 11101 34747 11135
rect 34980 11101 35014 11135
rect 37381 11101 37415 11135
rect 40049 11101 40083 11135
rect 46664 11101 46698 11135
rect 48237 11101 48271 11135
rect 48504 11101 48538 11135
rect 51549 11101 51583 11135
rect 53656 11101 53690 11135
rect 12440 11033 12474 11067
rect 14372 11033 14406 11067
rect 20168 11033 20202 11067
rect 22376 11033 22410 11067
rect 37648 11033 37682 11067
rect 40776 11033 40810 11067
rect 51816 11033 51850 11067
rect 57152 11033 57186 11067
rect 10793 10965 10827 10999
rect 25789 10965 25823 10999
rect 47777 10965 47811 10999
rect 54769 10965 54803 10999
rect 58265 10965 58299 10999
rect 15485 10761 15519 10795
rect 21005 10761 21039 10795
rect 23213 10761 23247 10795
rect 33793 10761 33827 10795
rect 38669 10761 38703 10795
rect 41889 10761 41923 10795
rect 47041 10761 47075 10795
rect 48237 10761 48271 10795
rect 50353 10761 50387 10795
rect 55505 10761 55539 10795
rect 57345 10761 57379 10795
rect 9588 10693 9622 10727
rect 14350 10693 14384 10727
rect 16948 10693 16982 10727
rect 22100 10693 22134 10727
rect 24308 10693 24342 10727
rect 32680 10693 32714 10727
rect 34520 10693 34554 10727
rect 44088 10693 44122 10727
rect 45928 10693 45962 10727
rect 54392 10693 54426 10727
rect 56232 10693 56266 10727
rect 9321 10625 9355 10659
rect 11796 10625 11830 10659
rect 16681 10625 16715 10659
rect 19173 10625 19207 10659
rect 19892 10625 19926 10659
rect 24041 10625 24075 10659
rect 27629 10625 27663 10659
rect 27896 10625 27930 10659
rect 32413 10625 32447 10659
rect 37556 10625 37590 10659
rect 40509 10625 40543 10659
rect 40776 10625 40810 10659
rect 43821 10625 43855 10659
rect 45661 10625 45695 10659
rect 48421 10625 48455 10659
rect 49240 10625 49274 10659
rect 50813 10625 50847 10659
rect 51080 10625 51114 10659
rect 54125 10625 54159 10659
rect 11529 10557 11563 10591
rect 14105 10557 14139 10591
rect 19625 10557 19659 10591
rect 21833 10557 21867 10591
rect 34253 10557 34287 10591
rect 37289 10557 37323 10591
rect 48973 10557 49007 10591
rect 55965 10557 55999 10591
rect 10701 10421 10735 10455
rect 12909 10421 12943 10455
rect 18061 10421 18095 10455
rect 18981 10421 19015 10455
rect 25421 10421 25455 10455
rect 29009 10421 29043 10455
rect 35633 10421 35667 10455
rect 45201 10421 45235 10455
rect 52193 10421 52227 10455
rect 16129 10217 16163 10251
rect 17969 10217 18003 10251
rect 20913 10217 20947 10251
rect 38577 10217 38611 10251
rect 44465 10217 44499 10251
rect 48605 10217 48639 10251
rect 52929 10217 52963 10251
rect 54769 10217 54803 10251
rect 6101 10081 6135 10115
rect 9137 10081 9171 10115
rect 10977 10081 11011 10115
rect 28457 10081 28491 10115
rect 29561 10081 29595 10115
rect 37197 10081 37231 10115
rect 53389 10081 53423 10115
rect 56885 10081 56919 10115
rect 9404 10013 9438 10047
rect 14749 10013 14783 10047
rect 16589 10013 16623 10047
rect 16856 10013 16890 10047
rect 19625 10013 19659 10047
rect 24409 10013 24443 10047
rect 24676 10013 24710 10047
rect 26709 10013 26743 10047
rect 32781 10013 32815 10047
rect 43085 10013 43119 10047
rect 45017 10013 45051 10047
rect 47317 10013 47351 10047
rect 51549 10013 51583 10047
rect 53656 10013 53690 10047
rect 6368 9945 6402 9979
rect 11222 9945 11256 9979
rect 15016 9945 15050 9979
rect 29828 9945 29862 9979
rect 33048 9945 33082 9979
rect 37464 9945 37498 9979
rect 43352 9945 43386 9979
rect 45284 9945 45318 9979
rect 51816 9945 51850 9979
rect 57152 9945 57186 9979
rect 59461 9945 59495 9979
rect 7481 9877 7515 9911
rect 10517 9877 10551 9911
rect 12357 9877 12391 9911
rect 25789 9877 25823 9911
rect 30941 9877 30975 9911
rect 34161 9877 34195 9911
rect 46397 9877 46431 9911
rect 58265 9877 58299 9911
rect 20729 9673 20763 9707
rect 30205 9673 30239 9707
rect 38669 9673 38703 9707
rect 41889 9673 41923 9707
rect 45661 9673 45695 9707
rect 50353 9673 50387 9707
rect 6644 9605 6678 9639
rect 9312 9605 9346 9639
rect 12909 9605 12943 9639
rect 16948 9605 16982 9639
rect 34060 9605 34094 9639
rect 49240 9605 49274 9639
rect 53656 9605 53690 9639
rect 56232 9605 56266 9639
rect 16681 9537 16715 9571
rect 19616 9537 19650 9571
rect 23213 9537 23247 9571
rect 23480 9537 23514 9571
rect 25053 9537 25087 9571
rect 25320 9537 25354 9571
rect 26985 9537 27019 9571
rect 27252 9537 27286 9571
rect 29092 9537 29126 9571
rect 37289 9537 37323 9571
rect 37545 9537 37579 9571
rect 40509 9537 40543 9571
rect 40776 9537 40810 9571
rect 42441 9537 42475 9571
rect 42708 9537 42742 9571
rect 44281 9537 44315 9571
rect 44548 9537 44582 9571
rect 48973 9537 49007 9571
rect 50813 9537 50847 9571
rect 51080 9537 51114 9571
rect 6377 9469 6411 9503
rect 9045 9469 9079 9503
rect 19349 9469 19383 9503
rect 28825 9469 28859 9503
rect 33793 9469 33827 9503
rect 53389 9469 53423 9503
rect 55965 9469 55999 9503
rect 18061 9401 18095 9435
rect 52193 9401 52227 9435
rect 57345 9401 57379 9435
rect 7757 9333 7791 9367
rect 10425 9333 10459 9367
rect 14197 9333 14231 9367
rect 24593 9333 24627 9367
rect 26433 9333 26467 9367
rect 28365 9333 28399 9367
rect 35173 9333 35207 9367
rect 43821 9333 43855 9367
rect 54769 9333 54803 9367
rect 7297 9129 7331 9163
rect 10333 9129 10367 9163
rect 15485 9129 15519 9163
rect 25789 9129 25823 9163
rect 27629 9129 27663 9163
rect 42073 9129 42107 9163
rect 43913 9129 43947 9163
rect 52561 9129 52595 9163
rect 5917 8993 5951 9027
rect 20361 8993 20395 9027
rect 26249 8993 26283 9027
rect 40693 8993 40727 9027
rect 51181 8993 51215 9027
rect 4077 8925 4111 8959
rect 6184 8925 6218 8959
rect 8953 8925 8987 8959
rect 9220 8925 9254 8959
rect 10793 8925 10827 8959
rect 14105 8925 14139 8959
rect 14372 8925 14406 8959
rect 22201 8925 22235 8959
rect 24409 8925 24443 8959
rect 24676 8925 24710 8959
rect 26516 8925 26550 8959
rect 29561 8925 29595 8959
rect 32413 8925 32447 8959
rect 34713 8925 34747 8959
rect 36553 8925 36587 8959
rect 42533 8925 42567 8959
rect 45017 8925 45051 8959
rect 46857 8925 46891 8959
rect 51448 8925 51482 8959
rect 53021 8925 53055 8959
rect 55321 8925 55355 8959
rect 57161 8925 57195 8959
rect 4344 8857 4378 8891
rect 11038 8857 11072 8891
rect 20628 8857 20662 8891
rect 22468 8857 22502 8891
rect 29828 8857 29862 8891
rect 34958 8857 34992 8891
rect 36798 8857 36832 8891
rect 40960 8857 40994 8891
rect 42778 8857 42812 8891
rect 45262 8857 45296 8891
rect 47124 8857 47158 8891
rect 53288 8857 53322 8891
rect 55588 8857 55622 8891
rect 57428 8857 57462 8891
rect 5457 8789 5491 8823
rect 12173 8789 12207 8823
rect 21741 8789 21775 8823
rect 23581 8789 23615 8823
rect 30941 8789 30975 8823
rect 33701 8789 33735 8823
rect 36093 8789 36127 8823
rect 37933 8789 37967 8823
rect 46397 8789 46431 8823
rect 48237 8789 48271 8823
rect 54401 8789 54435 8823
rect 56701 8789 56735 8823
rect 58541 8789 58575 8823
rect 10425 8585 10459 8619
rect 13645 8585 13679 8619
rect 20545 8585 20579 8619
rect 23397 8585 23431 8619
rect 25237 8585 25271 8619
rect 28365 8585 28399 8619
rect 30205 8585 30239 8619
rect 34805 8585 34839 8619
rect 36645 8585 36679 8619
rect 45661 8585 45695 8619
rect 48973 8585 49007 8619
rect 54125 8585 54159 8619
rect 4712 8517 4746 8551
rect 6644 8517 6678 8551
rect 9312 8517 9346 8551
rect 12510 8517 12544 8551
rect 19432 8517 19466 8551
rect 22284 8517 22318 8551
rect 29070 8517 29104 8551
rect 33692 8517 33726 8551
rect 37556 8517 37590 8551
rect 44548 8517 44582 8551
rect 49678 8517 49712 8551
rect 54861 8517 54895 8551
rect 4445 8449 4479 8483
rect 14556 8449 14590 8483
rect 24124 8449 24158 8483
rect 26985 8449 27019 8483
rect 27252 8449 27286 8483
rect 35265 8449 35299 8483
rect 35532 8449 35566 8483
rect 37289 8449 37323 8483
rect 39385 8449 39419 8483
rect 42697 8449 42731 8483
rect 44281 8449 44315 8483
rect 47593 8449 47627 8483
rect 47860 8449 47894 8483
rect 49433 8449 49467 8483
rect 52745 8449 52779 8483
rect 53012 8449 53046 8483
rect 6377 8381 6411 8415
rect 9045 8381 9079 8415
rect 12265 8381 12299 8415
rect 14289 8381 14323 8415
rect 19165 8381 19199 8415
rect 22017 8381 22051 8415
rect 23857 8381 23891 8415
rect 28825 8381 28859 8415
rect 33425 8381 33459 8415
rect 39129 8381 39163 8415
rect 42441 8381 42475 8415
rect 5825 8313 5859 8347
rect 15669 8313 15703 8347
rect 43821 8313 43855 8347
rect 7757 8245 7791 8279
rect 38669 8245 38703 8279
rect 40509 8245 40543 8279
rect 50813 8245 50847 8279
rect 56149 8245 56183 8279
rect 7297 8041 7331 8075
rect 11713 8041 11747 8075
rect 23029 8041 23063 8075
rect 25789 8041 25823 8075
rect 27629 8041 27663 8075
rect 30941 8041 30975 8075
rect 36093 8041 36127 8075
rect 38853 8041 38887 8075
rect 43085 8041 43119 8075
rect 46397 8041 46431 8075
rect 48237 8041 48271 8075
rect 54125 8041 54159 8075
rect 56701 8041 56735 8075
rect 58541 8041 58575 8075
rect 26249 7905 26283 7939
rect 46857 7905 46891 7939
rect 50169 7905 50203 7939
rect 52745 7905 52779 7939
rect 1869 7837 1903 7871
rect 4077 7837 4111 7871
rect 5917 7837 5951 7871
rect 6184 7837 6218 7871
rect 10333 7837 10367 7871
rect 12173 7837 12207 7871
rect 14473 7837 14507 7871
rect 16313 7837 16347 7871
rect 19349 7837 19383 7871
rect 21649 7837 21683 7871
rect 21916 7837 21950 7871
rect 24409 7837 24443 7871
rect 26516 7837 26550 7871
rect 29561 7837 29595 7871
rect 29828 7837 29862 7871
rect 32137 7837 32171 7871
rect 32393 7837 32427 7871
rect 34713 7837 34747 7871
rect 34980 7837 35014 7871
rect 37473 7837 37507 7871
rect 37740 7837 37774 7871
rect 41797 7837 41831 7871
rect 45017 7837 45051 7871
rect 47124 7837 47158 7871
rect 55321 7837 55355 7871
rect 57161 7837 57195 7871
rect 2136 7769 2170 7803
rect 4344 7769 4378 7803
rect 10600 7769 10634 7803
rect 12440 7769 12474 7803
rect 14740 7769 14774 7803
rect 16580 7769 16614 7803
rect 19616 7769 19650 7803
rect 24676 7769 24710 7803
rect 45284 7769 45318 7803
rect 50436 7769 50470 7803
rect 53012 7769 53046 7803
rect 55588 7769 55622 7803
rect 57406 7769 57440 7803
rect 3249 7701 3283 7735
rect 5457 7701 5491 7735
rect 13553 7701 13587 7735
rect 15853 7701 15887 7735
rect 17693 7701 17727 7735
rect 20729 7701 20763 7735
rect 33517 7701 33551 7735
rect 51549 7701 51583 7735
rect 5365 7497 5399 7531
rect 21097 7497 21131 7531
rect 25237 7497 25271 7531
rect 28365 7497 28399 7531
rect 36737 7497 36771 7531
rect 40049 7497 40083 7531
rect 41889 7497 41923 7531
rect 44189 7497 44223 7531
rect 50353 7497 50387 7531
rect 54125 7497 54159 7531
rect 55965 7497 55999 7531
rect 2320 7429 2354 7463
rect 4077 7429 4111 7463
rect 13176 7429 13210 7463
rect 15016 7429 15050 7463
rect 18144 7429 18178 7463
rect 27252 7429 27286 7463
rect 29828 7429 29862 7463
rect 32404 7429 32438 7463
rect 38936 7429 38970 7463
rect 43076 7429 43110 7463
rect 49240 7429 49274 7463
rect 54830 7429 54864 7463
rect 2053 7361 2087 7395
rect 7012 7361 7046 7395
rect 8585 7361 8619 7395
rect 8852 7361 8886 7395
rect 14749 7361 14783 7395
rect 17877 7361 17911 7395
rect 19984 7361 20018 7395
rect 24124 7361 24158 7395
rect 26985 7361 27019 7395
rect 35357 7361 35391 7395
rect 35624 7361 35658 7395
rect 40776 7361 40810 7395
rect 45928 7361 45962 7395
rect 51080 7361 51114 7395
rect 52745 7361 52779 7395
rect 53012 7361 53046 7395
rect 54585 7361 54619 7395
rect 6745 7293 6779 7327
rect 12909 7293 12943 7327
rect 19717 7293 19751 7327
rect 23857 7293 23891 7327
rect 29561 7293 29595 7327
rect 32137 7293 32171 7327
rect 38669 7293 38703 7327
rect 40509 7293 40543 7327
rect 42809 7293 42843 7327
rect 45661 7293 45695 7327
rect 48973 7293 49007 7327
rect 50813 7293 50847 7327
rect 30941 7225 30975 7259
rect 3433 7157 3467 7191
rect 8125 7157 8159 7191
rect 9965 7157 9999 7191
rect 14289 7157 14323 7191
rect 16129 7157 16163 7191
rect 19257 7157 19291 7191
rect 33517 7157 33551 7191
rect 47041 7157 47075 7191
rect 52193 7157 52227 7191
rect 6561 6953 6595 6987
rect 8401 6953 8435 6987
rect 13553 6953 13587 6987
rect 21189 6953 21223 6987
rect 25789 6953 25823 6987
rect 39221 6953 39255 6987
rect 47133 6953 47167 6987
rect 51549 6953 51583 6987
rect 54217 6953 54251 6987
rect 56701 6953 56735 6987
rect 58541 6953 58575 6987
rect 59461 6953 59495 6987
rect 15117 6817 15151 6851
rect 17325 6817 17359 6851
rect 24409 6817 24443 6851
rect 32689 6817 32723 6851
rect 40601 6817 40635 6851
rect 52837 6817 52871 6851
rect 1869 6749 1903 6783
rect 5181 6749 5215 6783
rect 5448 6749 5482 6783
rect 7021 6749 7055 6783
rect 8953 6749 8987 6783
rect 12173 6749 12207 6783
rect 12440 6749 12474 6783
rect 15384 6749 15418 6783
rect 17592 6749 17626 6783
rect 19809 6749 19843 6783
rect 22477 6749 22511 6783
rect 27629 6749 27663 6783
rect 30849 6749 30883 6783
rect 31116 6749 31150 6783
rect 36001 6749 36035 6783
rect 37841 6749 37875 6783
rect 43085 6749 43119 6783
rect 45753 6749 45787 6783
rect 47593 6749 47627 6783
rect 47860 6749 47894 6783
rect 50169 6749 50203 6783
rect 50436 6749 50470 6783
rect 55321 6749 55355 6783
rect 55588 6749 55622 6783
rect 57161 6749 57195 6783
rect 57428 6749 57462 6783
rect 2136 6681 2170 6715
rect 7288 6681 7322 6715
rect 9220 6681 9254 6715
rect 20076 6681 20110 6715
rect 22744 6681 22778 6715
rect 24676 6681 24710 6715
rect 27896 6681 27930 6715
rect 32934 6681 32968 6715
rect 36268 6681 36302 6715
rect 38086 6681 38120 6715
rect 40868 6681 40902 6715
rect 43352 6681 43386 6715
rect 46020 6681 46054 6715
rect 53104 6681 53138 6715
rect 3249 6613 3283 6647
rect 10333 6613 10367 6647
rect 16497 6613 16531 6647
rect 18705 6613 18739 6647
rect 23857 6613 23891 6647
rect 29009 6613 29043 6647
rect 32229 6613 32263 6647
rect 34069 6613 34103 6647
rect 37381 6613 37415 6647
rect 41981 6613 42015 6647
rect 44465 6613 44499 6647
rect 48973 6613 49007 6647
rect 5273 6409 5307 6443
rect 8677 6409 8711 6443
rect 10793 6409 10827 6443
rect 13277 6409 13311 6443
rect 16129 6409 16163 6443
rect 18337 6409 18371 6443
rect 20913 6409 20947 6443
rect 23489 6409 23523 6443
rect 25789 6409 25823 6443
rect 36737 6409 36771 6443
rect 41245 6409 41279 6443
rect 49341 6409 49375 6443
rect 54677 6409 54711 6443
rect 2320 6341 2354 6375
rect 4160 6341 4194 6375
rect 9658 6341 9692 6375
rect 12164 6341 12198 6375
rect 15016 6341 15050 6375
rect 17224 6341 17258 6375
rect 24654 6341 24688 6375
rect 32404 6341 32438 6375
rect 38292 6341 38326 6375
rect 48228 6341 48262 6375
rect 50068 6341 50102 6375
rect 2053 6273 2087 6307
rect 3893 6273 3927 6307
rect 7205 6273 7239 6307
rect 11897 6273 11931 6307
rect 14749 6273 14783 6307
rect 19800 6273 19834 6307
rect 22109 6273 22143 6307
rect 22376 6273 22410 6307
rect 27252 6273 27286 6307
rect 29745 6273 29779 6307
rect 30012 6273 30046 6307
rect 35624 6273 35658 6307
rect 40132 6273 40166 6307
rect 43821 6273 43855 6307
rect 44088 6273 44122 6307
rect 45928 6273 45962 6307
rect 47961 6273 47995 6307
rect 49801 6273 49835 6307
rect 53564 6273 53598 6307
rect 9413 6205 9447 6239
rect 16957 6205 16991 6239
rect 19533 6205 19567 6239
rect 24409 6205 24443 6239
rect 26985 6205 27019 6239
rect 32137 6205 32171 6239
rect 35357 6205 35391 6239
rect 38025 6205 38059 6239
rect 39865 6205 39899 6239
rect 45661 6205 45695 6239
rect 53297 6205 53331 6239
rect 3433 6069 3467 6103
rect 28365 6069 28399 6103
rect 31125 6069 31159 6103
rect 33517 6069 33551 6103
rect 39405 6069 39439 6103
rect 45201 6069 45235 6103
rect 47041 6069 47075 6103
rect 51181 6069 51215 6103
rect 10333 5865 10367 5899
rect 17693 5865 17727 5899
rect 20637 5865 20671 5899
rect 23213 5865 23247 5899
rect 29009 5865 29043 5899
rect 30941 5865 30975 5899
rect 36369 5865 36403 5899
rect 41705 5865 41739 5899
rect 52745 5865 52779 5899
rect 3985 5729 4019 5763
rect 5825 5729 5859 5763
rect 8953 5729 8987 5763
rect 10793 5729 10827 5763
rect 16313 5729 16347 5763
rect 27629 5729 27663 5763
rect 29561 5729 29595 5763
rect 32689 5729 32723 5763
rect 40325 5729 40359 5763
rect 4241 5661 4275 5695
rect 9220 5661 9254 5695
rect 14473 5661 14507 5695
rect 16580 5661 16614 5695
rect 19257 5661 19291 5695
rect 21833 5661 21867 5695
rect 25789 5661 25823 5695
rect 26056 5661 26090 5695
rect 27896 5661 27930 5695
rect 32956 5661 32990 5695
rect 37933 5661 37967 5695
rect 38200 5661 38234 5695
rect 43085 5661 43119 5695
rect 43352 5661 43386 5695
rect 45017 5661 45051 5695
rect 45284 5661 45318 5695
rect 51457 5661 51491 5695
rect 6092 5593 6126 5627
rect 11060 5593 11094 5627
rect 14740 5593 14774 5627
rect 19524 5593 19558 5627
rect 22100 5593 22134 5627
rect 29828 5593 29862 5627
rect 35081 5593 35115 5627
rect 40592 5593 40626 5627
rect 46857 5593 46891 5627
rect 5365 5525 5399 5559
rect 7205 5525 7239 5559
rect 12173 5525 12207 5559
rect 15853 5525 15887 5559
rect 27169 5525 27203 5559
rect 34069 5525 34103 5559
rect 39313 5525 39347 5559
rect 44465 5525 44499 5559
rect 46397 5525 46431 5559
rect 48145 5525 48179 5559
rect 3801 5321 3835 5355
rect 10609 5321 10643 5355
rect 45385 5321 45419 5355
rect 51549 5321 51583 5355
rect 54217 5321 54251 5355
rect 4506 5253 4540 5287
rect 6644 5253 6678 5287
rect 9496 5253 9530 5287
rect 11989 5253 12023 5287
rect 20168 5253 20202 5287
rect 29745 5253 29779 5287
rect 32772 5253 32806 5287
rect 35440 5253 35474 5287
rect 39589 5253 39623 5287
rect 44272 5253 44306 5287
rect 48596 5253 48630 5287
rect 50436 5253 50470 5287
rect 2421 5185 2455 5219
rect 2688 5185 2722 5219
rect 6377 5185 6411 5219
rect 9229 5185 9263 5219
rect 14464 5185 14498 5219
rect 23397 5185 23431 5219
rect 28181 5185 28215 5219
rect 32505 5185 32539 5219
rect 38016 5185 38050 5219
rect 44005 5185 44039 5219
rect 48329 5185 48363 5219
rect 52837 5185 52871 5219
rect 53104 5185 53138 5219
rect 4261 5117 4295 5151
rect 14197 5117 14231 5151
rect 19901 5117 19935 5151
rect 35173 5117 35207 5151
rect 37749 5117 37783 5151
rect 41337 5117 41371 5151
rect 50169 5117 50203 5151
rect 5641 4981 5675 5015
rect 7757 4981 7791 5015
rect 13277 4981 13311 5015
rect 15577 4981 15611 5015
rect 21281 4981 21315 5015
rect 24685 4981 24719 5015
rect 33885 4981 33919 5015
rect 36553 4981 36587 5015
rect 39129 4981 39163 5015
rect 49709 4981 49743 5015
rect 15485 4777 15519 4811
rect 21465 4777 21499 4811
rect 23305 4777 23339 4811
rect 36737 4777 36771 4811
rect 41245 4777 41279 4811
rect 48973 4777 49007 4811
rect 9781 4641 9815 4675
rect 11621 4641 11655 4675
rect 15945 4641 15979 4675
rect 26985 4641 27019 4675
rect 30021 4641 30055 4675
rect 3801 4573 3835 4607
rect 4068 4573 4102 4607
rect 5641 4573 5675 4607
rect 10048 4573 10082 4607
rect 14105 4573 14139 4607
rect 20085 4573 20119 4607
rect 21925 4573 21959 4607
rect 25145 4573 25179 4607
rect 27252 4573 27286 4607
rect 30288 4573 30322 4607
rect 32781 4573 32815 4607
rect 33048 4573 33082 4607
rect 35357 4573 35391 4607
rect 35624 4573 35658 4607
rect 37197 4573 37231 4607
rect 39865 4573 39899 4607
rect 40121 4573 40155 4607
rect 41705 4573 41739 4607
rect 47593 4573 47627 4607
rect 47849 4573 47883 4607
rect 50169 4573 50203 4607
rect 50436 4573 50470 4607
rect 52009 4573 52043 4607
rect 5886 4505 5920 4539
rect 11866 4505 11900 4539
rect 14372 4505 14406 4539
rect 16212 4505 16246 4539
rect 20352 4505 20386 4539
rect 22192 4505 22226 4539
rect 25412 4505 25446 4539
rect 37464 4505 37498 4539
rect 41950 4505 41984 4539
rect 52276 4505 52310 4539
rect 5181 4437 5215 4471
rect 7021 4437 7055 4471
rect 11161 4437 11195 4471
rect 13001 4437 13035 4471
rect 17325 4437 17359 4471
rect 26525 4437 26559 4471
rect 28365 4437 28399 4471
rect 31401 4437 31435 4471
rect 34161 4437 34195 4471
rect 38577 4437 38611 4471
rect 43085 4437 43119 4471
rect 51549 4437 51583 4471
rect 53389 4437 53423 4471
rect 14749 4233 14783 4267
rect 23213 4233 23247 4267
rect 18613 4165 18647 4199
rect 27230 4165 27264 4199
rect 53012 4165 53046 4199
rect 3709 4097 3743 4131
rect 3976 4097 4010 4131
rect 6377 4097 6411 4131
rect 6644 4097 6678 4131
rect 11529 4097 11563 4131
rect 11796 4097 11830 4131
rect 13625 4097 13659 4131
rect 16681 4097 16715 4131
rect 16937 4097 16971 4131
rect 21833 4097 21867 4131
rect 22100 4097 22134 4131
rect 24308 4097 24342 4131
rect 26985 4097 27019 4131
rect 30012 4097 30046 4131
rect 33048 4097 33082 4131
rect 34877 4097 34911 4131
rect 37289 4097 37323 4131
rect 37556 4097 37590 4131
rect 39129 4097 39163 4131
rect 39396 4097 39430 4131
rect 44272 4097 44306 4131
rect 47849 4097 47883 4131
rect 49893 4097 49927 4131
rect 50160 4097 50194 4131
rect 52745 4097 52779 4131
rect 13369 4029 13403 4063
rect 20361 4029 20395 4063
rect 24041 4029 24075 4063
rect 29745 4029 29779 4063
rect 32781 4029 32815 4063
rect 34621 4029 34655 4063
rect 44005 4029 44039 4063
rect 47593 4029 47627 4063
rect 5089 3961 5123 3995
rect 7757 3961 7791 3995
rect 34161 3961 34195 3995
rect 36001 3961 36035 3995
rect 45385 3961 45419 3995
rect 12909 3893 12943 3927
rect 18061 3893 18095 3927
rect 25421 3893 25455 3927
rect 28365 3893 28399 3927
rect 31125 3893 31159 3927
rect 38669 3893 38703 3927
rect 40509 3893 40543 3927
rect 48973 3893 49007 3927
rect 51273 3893 51307 3927
rect 54125 3893 54159 3927
rect 6009 3689 6043 3723
rect 11805 3689 11839 3723
rect 15485 3689 15519 3723
rect 17325 3689 17359 3723
rect 22477 3689 22511 3723
rect 31033 3689 31067 3723
rect 41245 3689 41279 3723
rect 43821 3689 43855 3723
rect 49617 3689 49651 3723
rect 53573 3689 53607 3723
rect 4629 3553 4663 3587
rect 10425 3553 10459 3587
rect 14105 3553 14139 3587
rect 15945 3553 15979 3587
rect 26709 3553 26743 3587
rect 32597 3553 32631 3587
rect 34713 3553 34747 3587
rect 39865 3553 39899 3587
rect 42441 3553 42475 3587
rect 4896 3485 4930 3519
rect 10692 3485 10726 3519
rect 16212 3485 16246 3519
rect 19257 3485 19291 3519
rect 21097 3485 21131 3519
rect 24869 3485 24903 3519
rect 26976 3485 27010 3519
rect 29653 3485 29687 3519
rect 29920 3485 29954 3519
rect 36553 3485 36587 3519
rect 40132 3485 40166 3519
rect 42708 3485 42742 3519
rect 48237 3485 48271 3519
rect 48504 3485 48538 3519
rect 50353 3485 50387 3519
rect 50620 3485 50654 3519
rect 52193 3485 52227 3519
rect 14372 3417 14406 3451
rect 19502 3417 19536 3451
rect 21364 3417 21398 3451
rect 25136 3417 25170 3451
rect 32864 3417 32898 3451
rect 34958 3417 34992 3451
rect 36798 3417 36832 3451
rect 52438 3417 52472 3451
rect 20637 3349 20671 3383
rect 26249 3349 26283 3383
rect 28089 3349 28123 3383
rect 33977 3349 34011 3383
rect 36093 3349 36127 3383
rect 37933 3349 37967 3383
rect 51733 3349 51767 3383
rect 14749 3145 14783 3179
rect 18061 3145 18095 3179
rect 23857 3145 23891 3179
rect 25697 3145 25731 3179
rect 30205 3145 30239 3179
rect 34069 3145 34103 3179
rect 35909 3145 35943 3179
rect 40509 3145 40543 3179
rect 43821 3145 43855 3179
rect 52193 3145 52227 3179
rect 11796 3077 11830 3111
rect 13636 3077 13670 3111
rect 16948 3077 16982 3111
rect 22744 3077 22778 3111
rect 24584 3077 24618 3111
rect 27252 3077 27286 3111
rect 32956 3077 32990 3111
rect 34796 3077 34830 3111
rect 39374 3077 39408 3111
rect 42708 3077 42742 3111
rect 51080 3077 51114 3111
rect 53012 3077 53046 3111
rect 11529 3009 11563 3043
rect 13369 3009 13403 3043
rect 16681 3009 16715 3043
rect 18521 3009 18555 3043
rect 18777 3009 18811 3043
rect 22477 3009 22511 3043
rect 29081 3009 29115 3043
rect 32689 3009 32723 3043
rect 34529 3009 34563 3043
rect 37289 3009 37323 3043
rect 37556 3009 37590 3043
rect 39129 3009 39163 3043
rect 42441 3009 42475 3043
rect 50813 3009 50847 3043
rect 52745 3009 52779 3043
rect 24317 2941 24351 2975
rect 26985 2941 27019 2975
rect 28825 2941 28859 2975
rect 38669 2873 38703 2907
rect 54125 2873 54159 2907
rect 12909 2805 12943 2839
rect 19901 2805 19935 2839
rect 28365 2805 28399 2839
rect 18613 2601 18647 2635
rect 23213 2601 23247 2635
rect 25789 2601 25823 2635
rect 28365 2601 28399 2635
rect 33977 2601 34011 2635
rect 36093 2601 36127 2635
rect 38669 2601 38703 2635
rect 13093 2533 13127 2567
rect 11713 2465 11747 2499
rect 17233 2465 17267 2499
rect 24409 2465 24443 2499
rect 26985 2465 27019 2499
rect 34713 2465 34747 2499
rect 37289 2465 37323 2499
rect 1685 2397 1719 2431
rect 1961 2397 1995 2431
rect 11980 2397 12014 2431
rect 17500 2397 17534 2431
rect 19901 2397 19935 2431
rect 20157 2397 20191 2431
rect 21833 2397 21867 2431
rect 24676 2397 24710 2431
rect 27252 2397 27286 2431
rect 34161 2397 34195 2431
rect 34980 2397 35014 2431
rect 37556 2397 37590 2431
rect 1777 2329 1811 2363
rect 22078 2329 22112 2363
rect 21281 2261 21315 2295
<< metal1 >>
rect 1104 60410 59340 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 34934 60410
rect 34986 60358 34998 60410
rect 35050 60358 35062 60410
rect 35114 60358 35126 60410
rect 35178 60358 35190 60410
rect 35242 60358 59340 60410
rect 1104 60336 59340 60358
rect 26234 60188 26240 60240
rect 26292 60228 26298 60240
rect 27341 60231 27399 60237
rect 27341 60228 27353 60231
rect 26292 60200 27353 60228
rect 26292 60188 26298 60200
rect 27341 60197 27353 60200
rect 27387 60197 27399 60231
rect 27341 60191 27399 60197
rect 38841 60231 38899 60237
rect 38841 60197 38853 60231
rect 38887 60228 38899 60231
rect 39669 60231 39727 60237
rect 39669 60228 39681 60231
rect 38887 60200 39681 60228
rect 38887 60197 38899 60200
rect 38841 60191 38899 60197
rect 39669 60197 39681 60200
rect 39715 60197 39727 60231
rect 39669 60191 39727 60197
rect 58621 60231 58679 60237
rect 58621 60197 58633 60231
rect 58667 60228 58679 60231
rect 60366 60228 60372 60240
rect 58667 60200 60372 60228
rect 58667 60197 58679 60200
rect 58621 60191 58679 60197
rect 60366 60188 60372 60200
rect 60424 60188 60430 60240
rect 30944 60132 32260 60160
rect 6457 60095 6515 60101
rect 6457 60061 6469 60095
rect 6503 60061 6515 60095
rect 6457 60055 6515 60061
rect 6472 59956 6500 60055
rect 11514 60052 11520 60104
rect 11572 60092 11578 60104
rect 11701 60095 11759 60101
rect 11701 60092 11713 60095
rect 11572 60064 11713 60092
rect 11572 60052 11578 60064
rect 11701 60061 11713 60064
rect 11747 60061 11759 60095
rect 29914 60092 29920 60104
rect 29875 60064 29920 60092
rect 11701 60055 11759 60061
rect 29914 60052 29920 60064
rect 29972 60052 29978 60104
rect 30944 60092 30972 60132
rect 32122 60092 32128 60104
rect 30024 60064 30972 60092
rect 32083 60064 32128 60092
rect 6724 60027 6782 60033
rect 6724 59993 6736 60027
rect 6770 60024 6782 60027
rect 7742 60024 7748 60036
rect 6770 59996 7748 60024
rect 6770 59993 6782 59996
rect 6724 59987 6782 59993
rect 7742 59984 7748 59996
rect 7800 59984 7806 60036
rect 11968 60027 12026 60033
rect 11968 59993 11980 60027
rect 12014 60024 12026 60027
rect 12894 60024 12900 60036
rect 12014 59996 12900 60024
rect 12014 59993 12026 59996
rect 11968 59987 12026 59993
rect 12894 59984 12900 59996
rect 12952 59984 12958 60036
rect 27249 60027 27307 60033
rect 27249 59993 27261 60027
rect 27295 60024 27307 60027
rect 27525 60027 27583 60033
rect 27525 60024 27537 60027
rect 27295 59996 27537 60024
rect 27295 59993 27307 59996
rect 27249 59987 27307 59993
rect 27525 59993 27537 59996
rect 27571 60024 27583 60027
rect 28442 60024 28448 60036
rect 27571 59996 28448 60024
rect 27571 59993 27583 59996
rect 27525 59987 27583 59993
rect 28442 59984 28448 59996
rect 28500 60024 28506 60036
rect 30024 60024 30052 60064
rect 32122 60052 32128 60064
rect 32180 60052 32186 60104
rect 32232 60092 32260 60132
rect 34054 60092 34060 60104
rect 32232 60064 34060 60092
rect 34054 60052 34060 60064
rect 34112 60052 34118 60104
rect 35345 60095 35403 60101
rect 35345 60061 35357 60095
rect 35391 60092 35403 60095
rect 37461 60095 37519 60101
rect 37461 60092 37473 60095
rect 35391 60064 37473 60092
rect 35391 60061 35403 60064
rect 35345 60055 35403 60061
rect 37461 60061 37473 60064
rect 37507 60092 37519 60095
rect 37550 60092 37556 60104
rect 37507 60064 37556 60092
rect 37507 60061 37519 60064
rect 37461 60055 37519 60061
rect 37550 60052 37556 60064
rect 37608 60092 37614 60104
rect 39853 60095 39911 60101
rect 39853 60092 39865 60095
rect 37608 60064 39865 60092
rect 37608 60052 37614 60064
rect 39853 60061 39865 60064
rect 39899 60092 39911 60095
rect 40402 60092 40408 60104
rect 39899 60064 40408 60092
rect 39899 60061 39911 60064
rect 39853 60055 39911 60061
rect 40402 60052 40408 60064
rect 40460 60052 40466 60104
rect 43622 60052 43628 60104
rect 43680 60092 43686 60104
rect 45005 60095 45063 60101
rect 45005 60092 45017 60095
rect 43680 60064 45017 60092
rect 43680 60052 43686 60064
rect 45005 60061 45017 60064
rect 45051 60092 45063 60095
rect 45554 60092 45560 60104
rect 45051 60064 45560 60092
rect 45051 60061 45063 60064
rect 45005 60055 45063 60061
rect 45554 60052 45560 60064
rect 45612 60092 45618 60104
rect 47765 60095 47823 60101
rect 47765 60092 47777 60095
rect 45612 60064 47777 60092
rect 45612 60052 45618 60064
rect 47765 60061 47777 60064
rect 47811 60092 47823 60095
rect 48958 60092 48964 60104
rect 47811 60064 48964 60092
rect 47811 60061 47823 60064
rect 47765 60055 47823 60061
rect 48958 60052 48964 60064
rect 49016 60052 49022 60104
rect 50157 60095 50215 60101
rect 50157 60061 50169 60095
rect 50203 60092 50215 60095
rect 50798 60092 50804 60104
rect 50203 60064 50804 60092
rect 50203 60061 50215 60064
rect 50157 60055 50215 60061
rect 50798 60052 50804 60064
rect 50856 60052 50862 60104
rect 53377 60095 53435 60101
rect 53377 60061 53389 60095
rect 53423 60092 53435 60095
rect 54110 60092 54116 60104
rect 53423 60064 54116 60092
rect 53423 60061 53435 60064
rect 53377 60055 53435 60061
rect 54110 60052 54116 60064
rect 54168 60052 54174 60104
rect 28500 59996 30052 60024
rect 30184 60027 30242 60033
rect 28500 59984 28506 59996
rect 30184 59993 30196 60027
rect 30230 60024 30242 60027
rect 30230 59996 31524 60024
rect 30230 59993 30242 59996
rect 30184 59987 30242 59993
rect 6914 59956 6920 59968
rect 6472 59928 6920 59956
rect 6914 59916 6920 59928
rect 6972 59916 6978 59968
rect 7837 59959 7895 59965
rect 7837 59925 7849 59959
rect 7883 59956 7895 59959
rect 8478 59956 8484 59968
rect 7883 59928 8484 59956
rect 7883 59925 7895 59928
rect 7837 59919 7895 59925
rect 8478 59916 8484 59928
rect 8536 59916 8542 59968
rect 13078 59956 13084 59968
rect 13039 59928 13084 59956
rect 13078 59916 13084 59928
rect 13136 59916 13142 59968
rect 29362 59916 29368 59968
rect 29420 59956 29426 59968
rect 31297 59959 31355 59965
rect 31297 59956 31309 59959
rect 29420 59928 31309 59956
rect 29420 59916 29426 59928
rect 31297 59925 31309 59928
rect 31343 59925 31355 59959
rect 31496 59956 31524 59996
rect 31570 59984 31576 60036
rect 31628 60024 31634 60036
rect 32370 60027 32428 60033
rect 32370 60024 32382 60027
rect 31628 59996 32382 60024
rect 31628 59984 31634 59996
rect 32370 59993 32382 59996
rect 32416 59993 32428 60027
rect 32370 59987 32428 59993
rect 35612 60027 35670 60033
rect 35612 59993 35624 60027
rect 35658 60024 35670 60027
rect 37728 60027 37786 60033
rect 35658 59996 37688 60024
rect 35658 59993 35670 59996
rect 35612 59987 35670 59993
rect 33505 59959 33563 59965
rect 33505 59956 33517 59959
rect 31496 59928 33517 59956
rect 31297 59919 31355 59925
rect 33505 59925 33517 59928
rect 33551 59925 33563 59959
rect 36722 59956 36728 59968
rect 36683 59928 36728 59956
rect 33505 59919 33563 59925
rect 36722 59916 36728 59928
rect 36780 59916 36786 59968
rect 37660 59956 37688 59996
rect 37728 59993 37740 60027
rect 37774 60024 37786 60027
rect 38746 60024 38752 60036
rect 37774 59996 38752 60024
rect 37774 59993 37786 59996
rect 37728 59987 37786 59993
rect 38746 59984 38752 59996
rect 38804 59984 38810 60036
rect 39669 60027 39727 60033
rect 39669 59993 39681 60027
rect 39715 60024 39727 60027
rect 40098 60027 40156 60033
rect 40098 60024 40110 60027
rect 39715 59996 40110 60024
rect 39715 59993 39727 59996
rect 39669 59987 39727 59993
rect 40098 59993 40110 59996
rect 40144 59993 40156 60027
rect 40098 59987 40156 59993
rect 45272 60027 45330 60033
rect 45272 59993 45284 60027
rect 45318 60024 45330 60027
rect 46934 60024 46940 60036
rect 45318 59996 46940 60024
rect 45318 59993 45330 59996
rect 45272 59987 45330 59993
rect 46934 59984 46940 59996
rect 46992 59984 46998 60036
rect 48032 60027 48090 60033
rect 48032 59993 48044 60027
rect 48078 60024 48090 60027
rect 49326 60024 49332 60036
rect 48078 59996 49332 60024
rect 48078 59993 48090 59996
rect 48032 59987 48090 59993
rect 49326 59984 49332 59996
rect 49384 59984 49390 60036
rect 50424 60027 50482 60033
rect 50424 59993 50436 60027
rect 50470 60024 50482 60027
rect 50614 60024 50620 60036
rect 50470 59996 50620 60024
rect 50470 59993 50482 59996
rect 50424 59987 50482 59993
rect 50614 59984 50620 59996
rect 50672 59984 50678 60036
rect 53644 60027 53702 60033
rect 53644 59993 53656 60027
rect 53690 60024 53702 60027
rect 54938 60024 54944 60036
rect 53690 59996 54944 60024
rect 53690 59993 53702 59996
rect 53644 59987 53702 59993
rect 54938 59984 54944 59996
rect 54996 59984 55002 60036
rect 58434 60024 58440 60036
rect 58395 59996 58440 60024
rect 58434 59984 58440 59996
rect 58492 59984 58498 60036
rect 41233 59959 41291 59965
rect 41233 59956 41245 59959
rect 37660 59928 41245 59956
rect 41233 59925 41245 59928
rect 41279 59925 41291 59959
rect 41233 59919 41291 59925
rect 44174 59916 44180 59968
rect 44232 59956 44238 59968
rect 46385 59959 46443 59965
rect 46385 59956 46397 59959
rect 44232 59928 46397 59956
rect 44232 59916 44238 59928
rect 46385 59925 46397 59928
rect 46431 59925 46443 59959
rect 46385 59919 46443 59925
rect 48774 59916 48780 59968
rect 48832 59956 48838 59968
rect 49145 59959 49203 59965
rect 49145 59956 49157 59959
rect 48832 59928 49157 59956
rect 48832 59916 48838 59928
rect 49145 59925 49157 59928
rect 49191 59925 49203 59959
rect 51534 59956 51540 59968
rect 51495 59928 51540 59956
rect 49145 59919 49203 59925
rect 51534 59916 51540 59928
rect 51592 59916 51598 59968
rect 53190 59916 53196 59968
rect 53248 59956 53254 59968
rect 54757 59959 54815 59965
rect 54757 59956 54769 59959
rect 53248 59928 54769 59956
rect 53248 59916 53254 59928
rect 54757 59925 54769 59928
rect 54803 59925 54815 59959
rect 54757 59919 54815 59925
rect 1104 59866 59340 59888
rect 1104 59814 19574 59866
rect 19626 59814 19638 59866
rect 19690 59814 19702 59866
rect 19754 59814 19766 59866
rect 19818 59814 19830 59866
rect 19882 59814 50294 59866
rect 50346 59814 50358 59866
rect 50410 59814 50422 59866
rect 50474 59814 50486 59866
rect 50538 59814 50550 59866
rect 50602 59814 59340 59866
rect 1104 59792 59340 59814
rect 7742 59752 7748 59764
rect 7703 59724 7748 59752
rect 7742 59712 7748 59724
rect 7800 59712 7806 59764
rect 12894 59752 12900 59764
rect 12855 59724 12900 59752
rect 12894 59712 12900 59724
rect 12952 59712 12958 59764
rect 31570 59752 31576 59764
rect 31531 59724 31576 59752
rect 31570 59712 31576 59724
rect 31628 59712 31634 59764
rect 33965 59755 34023 59761
rect 33965 59721 33977 59755
rect 34011 59721 34023 59755
rect 33965 59715 34023 59721
rect 6914 59684 6920 59696
rect 6380 59656 6920 59684
rect 6380 59625 6408 59656
rect 6914 59644 6920 59656
rect 6972 59684 6978 59696
rect 27522 59684 27528 59696
rect 6972 59656 8248 59684
rect 6972 59644 6978 59656
rect 6365 59619 6423 59625
rect 6365 59585 6377 59619
rect 6411 59585 6423 59619
rect 6365 59579 6423 59585
rect 6632 59619 6690 59625
rect 6632 59585 6644 59619
rect 6678 59616 6690 59619
rect 8110 59616 8116 59628
rect 6678 59588 8116 59616
rect 6678 59585 6690 59588
rect 6632 59579 6690 59585
rect 8110 59576 8116 59588
rect 8168 59576 8174 59628
rect 8220 59625 8248 59656
rect 11532 59656 12434 59684
rect 8205 59619 8263 59625
rect 8205 59585 8217 59619
rect 8251 59585 8263 59619
rect 8205 59579 8263 59585
rect 8472 59619 8530 59625
rect 8472 59585 8484 59619
rect 8518 59616 8530 59619
rect 9490 59616 9496 59628
rect 8518 59588 9496 59616
rect 8518 59585 8530 59588
rect 8472 59579 8530 59585
rect 9490 59576 9496 59588
rect 9548 59576 9554 59628
rect 11532 59560 11560 59656
rect 11784 59619 11842 59625
rect 11784 59585 11796 59619
rect 11830 59616 11842 59619
rect 12250 59616 12256 59628
rect 11830 59588 12256 59616
rect 11830 59585 11842 59588
rect 11784 59579 11842 59585
rect 12250 59576 12256 59588
rect 12308 59576 12314 59628
rect 12406 59616 12434 59656
rect 22480 59656 24348 59684
rect 13357 59619 13415 59625
rect 13357 59616 13369 59619
rect 12406 59588 13369 59616
rect 13357 59585 13369 59588
rect 13403 59585 13415 59619
rect 13357 59579 13415 59585
rect 13624 59619 13682 59625
rect 13624 59585 13636 59619
rect 13670 59616 13682 59619
rect 14642 59616 14648 59628
rect 13670 59588 14648 59616
rect 13670 59585 13682 59588
rect 13624 59579 13682 59585
rect 14642 59576 14648 59588
rect 14700 59576 14706 59628
rect 19889 59619 19947 59625
rect 19889 59585 19901 59619
rect 19935 59616 19947 59619
rect 19978 59616 19984 59628
rect 19935 59588 19984 59616
rect 19935 59585 19947 59588
rect 19889 59579 19947 59585
rect 19978 59576 19984 59588
rect 20036 59576 20042 59628
rect 20156 59619 20214 59625
rect 20156 59585 20168 59619
rect 20202 59616 20214 59619
rect 21174 59616 21180 59628
rect 20202 59588 21180 59616
rect 20202 59585 20214 59588
rect 20156 59579 20214 59585
rect 21174 59576 21180 59588
rect 21232 59576 21238 59628
rect 22480 59560 22508 59656
rect 22732 59619 22790 59625
rect 22732 59585 22744 59619
rect 22778 59616 22790 59619
rect 23842 59616 23848 59628
rect 22778 59588 23848 59616
rect 22778 59585 22790 59588
rect 22732 59579 22790 59585
rect 23842 59576 23848 59588
rect 23900 59576 23906 59628
rect 24320 59625 24348 59656
rect 26988 59656 27528 59684
rect 24305 59619 24363 59625
rect 24305 59585 24317 59619
rect 24351 59585 24363 59619
rect 24305 59579 24363 59585
rect 24572 59619 24630 59625
rect 24572 59585 24584 59619
rect 24618 59616 24630 59619
rect 25958 59616 25964 59628
rect 24618 59588 25964 59616
rect 24618 59585 24630 59588
rect 24572 59579 24630 59585
rect 25958 59576 25964 59588
rect 26016 59576 26022 59628
rect 26988 59625 27016 59656
rect 27522 59644 27528 59656
rect 27580 59644 27586 59696
rect 30460 59687 30518 59693
rect 30460 59653 30472 59687
rect 30506 59684 30518 59687
rect 33980 59684 34008 59715
rect 38746 59712 38752 59764
rect 38804 59752 38810 59764
rect 38933 59755 38991 59761
rect 38933 59752 38945 59755
rect 38804 59724 38945 59752
rect 38804 59712 38810 59724
rect 38933 59721 38945 59724
rect 38979 59721 38991 59755
rect 46934 59752 46940 59764
rect 46895 59724 46940 59752
rect 38933 59715 38991 59721
rect 46934 59712 46940 59724
rect 46992 59712 46998 59764
rect 54938 59752 54944 59764
rect 54899 59724 54944 59752
rect 54938 59712 54944 59724
rect 54996 59712 55002 59764
rect 30506 59656 34008 59684
rect 30506 59653 30518 59656
rect 30460 59647 30518 59653
rect 34054 59644 34060 59696
rect 34112 59684 34118 59696
rect 55398 59684 55404 59696
rect 34112 59656 55404 59684
rect 34112 59644 34118 59656
rect 55398 59644 55404 59656
rect 55456 59644 55462 59696
rect 26973 59619 27031 59625
rect 26973 59585 26985 59619
rect 27019 59585 27031 59619
rect 26973 59579 27031 59585
rect 27240 59619 27298 59625
rect 27240 59585 27252 59619
rect 27286 59616 27298 59619
rect 28534 59616 28540 59628
rect 27286 59588 28540 59616
rect 27286 59585 27298 59588
rect 27240 59579 27298 59585
rect 28534 59576 28540 59588
rect 28592 59576 28598 59628
rect 29914 59576 29920 59628
rect 29972 59616 29978 59628
rect 30193 59619 30251 59625
rect 30193 59616 30205 59619
rect 29972 59588 30205 59616
rect 29972 59576 29978 59588
rect 30193 59585 30205 59588
rect 30239 59616 30251 59619
rect 30282 59616 30288 59628
rect 30239 59588 30288 59616
rect 30239 59585 30251 59588
rect 30193 59579 30251 59585
rect 30282 59576 30288 59588
rect 30340 59576 30346 59628
rect 31754 59576 31760 59628
rect 31812 59616 31818 59628
rect 32841 59619 32899 59625
rect 32841 59616 32853 59619
rect 31812 59588 32853 59616
rect 31812 59576 31818 59588
rect 32841 59585 32853 59588
rect 32887 59585 32899 59619
rect 32841 59579 32899 59585
rect 34692 59619 34750 59625
rect 34692 59585 34704 59619
rect 34738 59616 34750 59619
rect 35434 59616 35440 59628
rect 34738 59588 35440 59616
rect 34738 59585 34750 59588
rect 34692 59579 34750 59585
rect 35434 59576 35440 59588
rect 35492 59576 35498 59628
rect 37550 59616 37556 59628
rect 37511 59588 37556 59616
rect 37550 59576 37556 59588
rect 37608 59576 37614 59628
rect 37820 59619 37878 59625
rect 37820 59585 37832 59619
rect 37866 59616 37878 59619
rect 39022 59616 39028 59628
rect 37866 59588 39028 59616
rect 37866 59585 37878 59588
rect 37820 59579 37878 59585
rect 39022 59576 39028 59588
rect 39080 59576 39086 59628
rect 40672 59619 40730 59625
rect 40672 59585 40684 59619
rect 40718 59616 40730 59619
rect 41874 59616 41880 59628
rect 40718 59588 41880 59616
rect 40718 59585 40730 59588
rect 40672 59579 40730 59585
rect 41874 59576 41880 59588
rect 41932 59576 41938 59628
rect 43892 59619 43950 59625
rect 43892 59585 43904 59619
rect 43938 59616 43950 59619
rect 44450 59616 44456 59628
rect 43938 59588 44456 59616
rect 43938 59585 43950 59588
rect 43892 59579 43950 59585
rect 44450 59576 44456 59588
rect 44508 59576 44514 59628
rect 45554 59576 45560 59628
rect 45612 59616 45618 59628
rect 45824 59619 45882 59625
rect 45612 59588 45657 59616
rect 45612 59576 45618 59588
rect 45824 59585 45836 59619
rect 45870 59616 45882 59619
rect 47026 59616 47032 59628
rect 45870 59588 47032 59616
rect 45870 59585 45882 59588
rect 45824 59579 45882 59585
rect 47026 59576 47032 59588
rect 47084 59576 47090 59628
rect 48869 59619 48927 59625
rect 48869 59585 48881 59619
rect 48915 59616 48927 59619
rect 48958 59616 48964 59628
rect 48915 59588 48964 59616
rect 48915 59585 48927 59588
rect 48869 59579 48927 59585
rect 48958 59576 48964 59588
rect 49016 59576 49022 59628
rect 49136 59619 49194 59625
rect 49136 59585 49148 59619
rect 49182 59616 49194 59619
rect 49510 59616 49516 59628
rect 49182 59588 49516 59616
rect 49182 59585 49194 59588
rect 49136 59579 49194 59585
rect 49510 59576 49516 59588
rect 49568 59576 49574 59628
rect 51068 59619 51126 59625
rect 51068 59585 51080 59619
rect 51114 59616 51126 59619
rect 51902 59616 51908 59628
rect 51114 59588 51908 59616
rect 51114 59585 51126 59588
rect 51068 59579 51126 59585
rect 51902 59576 51908 59588
rect 51960 59576 51966 59628
rect 53828 59619 53886 59625
rect 53828 59585 53840 59619
rect 53874 59616 53886 59619
rect 54754 59616 54760 59628
rect 53874 59588 54760 59616
rect 53874 59585 53886 59588
rect 53828 59579 53886 59585
rect 54754 59576 54760 59588
rect 54812 59576 54818 59628
rect 54846 59576 54852 59628
rect 54904 59616 54910 59628
rect 56209 59619 56267 59625
rect 56209 59616 56221 59619
rect 54904 59588 56221 59616
rect 54904 59576 54910 59588
rect 56209 59585 56221 59588
rect 56255 59585 56267 59619
rect 56209 59579 56267 59585
rect 11514 59548 11520 59560
rect 11475 59520 11520 59548
rect 11514 59508 11520 59520
rect 11572 59508 11578 59560
rect 22462 59548 22468 59560
rect 22423 59520 22468 59548
rect 22462 59508 22468 59520
rect 22520 59508 22526 59560
rect 32122 59508 32128 59560
rect 32180 59548 32186 59560
rect 32585 59551 32643 59557
rect 32585 59548 32597 59551
rect 32180 59520 32597 59548
rect 32180 59508 32186 59520
rect 32585 59517 32597 59520
rect 32631 59517 32643 59551
rect 34422 59548 34428 59560
rect 34383 59520 34428 59548
rect 32585 59511 32643 59517
rect 9582 59412 9588 59424
rect 9543 59384 9588 59412
rect 9582 59372 9588 59384
rect 9640 59372 9646 59424
rect 14734 59412 14740 59424
rect 14695 59384 14740 59412
rect 14734 59372 14740 59384
rect 14792 59372 14798 59424
rect 20162 59372 20168 59424
rect 20220 59412 20226 59424
rect 21269 59415 21327 59421
rect 21269 59412 21281 59415
rect 20220 59384 21281 59412
rect 20220 59372 20226 59384
rect 21269 59381 21281 59384
rect 21315 59381 21327 59415
rect 21269 59375 21327 59381
rect 23474 59372 23480 59424
rect 23532 59412 23538 59424
rect 23845 59415 23903 59421
rect 23845 59412 23857 59415
rect 23532 59384 23857 59412
rect 23532 59372 23538 59384
rect 23845 59381 23857 59384
rect 23891 59381 23903 59415
rect 23845 59375 23903 59381
rect 23934 59372 23940 59424
rect 23992 59412 23998 59424
rect 25685 59415 25743 59421
rect 25685 59412 25697 59415
rect 23992 59384 25697 59412
rect 23992 59372 23998 59384
rect 25685 59381 25697 59384
rect 25731 59381 25743 59415
rect 25685 59375 25743 59381
rect 27246 59372 27252 59424
rect 27304 59412 27310 59424
rect 28353 59415 28411 59421
rect 28353 59412 28365 59415
rect 27304 59384 28365 59412
rect 27304 59372 27310 59384
rect 28353 59381 28365 59384
rect 28399 59381 28411 59415
rect 32600 59412 32628 59511
rect 34422 59508 34428 59520
rect 34480 59508 34486 59560
rect 40402 59548 40408 59560
rect 40363 59520 40408 59548
rect 40402 59508 40408 59520
rect 40460 59508 40466 59560
rect 43622 59548 43628 59560
rect 43583 59520 43628 59548
rect 43622 59508 43628 59520
rect 43680 59508 43686 59560
rect 50798 59548 50804 59560
rect 50759 59520 50804 59548
rect 50798 59508 50804 59520
rect 50856 59508 50862 59560
rect 53374 59508 53380 59560
rect 53432 59548 53438 59560
rect 53561 59551 53619 59557
rect 53561 59548 53573 59551
rect 53432 59520 53573 59548
rect 53432 59508 53438 59520
rect 53561 59517 53573 59520
rect 53607 59517 53619 59551
rect 53561 59511 53619 59517
rect 55858 59508 55864 59560
rect 55916 59548 55922 59560
rect 55953 59551 56011 59557
rect 55953 59548 55965 59551
rect 55916 59520 55965 59548
rect 55916 59508 55922 59520
rect 55953 59517 55965 59520
rect 55999 59517 56011 59551
rect 55953 59511 56011 59517
rect 32858 59412 32864 59424
rect 32600 59384 32864 59412
rect 28353 59375 28411 59381
rect 32858 59372 32864 59384
rect 32916 59372 32922 59424
rect 34606 59372 34612 59424
rect 34664 59412 34670 59424
rect 35805 59415 35863 59421
rect 35805 59412 35817 59415
rect 34664 59384 35817 59412
rect 34664 59372 34670 59384
rect 35805 59381 35817 59384
rect 35851 59381 35863 59415
rect 35805 59375 35863 59381
rect 40678 59372 40684 59424
rect 40736 59412 40742 59424
rect 41785 59415 41843 59421
rect 41785 59412 41797 59415
rect 40736 59384 41797 59412
rect 40736 59372 40742 59384
rect 41785 59381 41797 59384
rect 41831 59381 41843 59415
rect 41785 59375 41843 59381
rect 43346 59372 43352 59424
rect 43404 59412 43410 59424
rect 45005 59415 45063 59421
rect 45005 59412 45017 59415
rect 43404 59384 45017 59412
rect 43404 59372 43410 59384
rect 45005 59381 45017 59384
rect 45051 59381 45063 59415
rect 45005 59375 45063 59381
rect 48498 59372 48504 59424
rect 48556 59412 48562 59424
rect 50249 59415 50307 59421
rect 50249 59412 50261 59415
rect 48556 59384 50261 59412
rect 48556 59372 48562 59384
rect 50249 59381 50261 59384
rect 50295 59381 50307 59415
rect 50249 59375 50307 59381
rect 51074 59372 51080 59424
rect 51132 59412 51138 59424
rect 52181 59415 52239 59421
rect 52181 59412 52193 59415
rect 51132 59384 52193 59412
rect 51132 59372 51138 59384
rect 52181 59381 52193 59384
rect 52227 59381 52239 59415
rect 52181 59375 52239 59381
rect 55950 59372 55956 59424
rect 56008 59412 56014 59424
rect 57333 59415 57391 59421
rect 57333 59412 57345 59415
rect 56008 59384 57345 59412
rect 56008 59372 56014 59384
rect 57333 59381 57345 59384
rect 57379 59381 57391 59415
rect 57333 59375 57391 59381
rect 1104 59322 59340 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 34934 59322
rect 34986 59270 34998 59322
rect 35050 59270 35062 59322
rect 35114 59270 35126 59322
rect 35178 59270 35190 59322
rect 35242 59270 59340 59322
rect 1104 59248 59340 59270
rect 8110 59208 8116 59220
rect 8071 59180 8116 59208
rect 8110 59168 8116 59180
rect 8168 59168 8174 59220
rect 23842 59208 23848 59220
rect 23803 59180 23848 59208
rect 23842 59168 23848 59180
rect 23900 59168 23906 59220
rect 27522 59208 27528 59220
rect 25792 59180 27528 59208
rect 25792 59081 25820 59180
rect 27522 59168 27528 59180
rect 27580 59168 27586 59220
rect 39022 59208 39028 59220
rect 38983 59180 39028 59208
rect 39022 59168 39028 59180
rect 39080 59168 39086 59220
rect 44450 59208 44456 59220
rect 44411 59180 44456 59208
rect 44450 59168 44456 59180
rect 44508 59168 44514 59220
rect 54754 59208 54760 59220
rect 54715 59180 54760 59208
rect 54754 59168 54760 59180
rect 54812 59168 54818 59220
rect 56689 59211 56747 59217
rect 56689 59177 56701 59211
rect 56735 59208 56747 59211
rect 57514 59208 57520 59220
rect 56735 59180 57520 59208
rect 56735 59177 56747 59180
rect 56689 59171 56747 59177
rect 57514 59168 57520 59180
rect 57572 59208 57578 59220
rect 58434 59208 58440 59220
rect 57572 59180 58440 59208
rect 57572 59168 57578 59180
rect 58434 59168 58440 59180
rect 58492 59168 58498 59220
rect 25777 59075 25835 59081
rect 25777 59041 25789 59075
rect 25823 59041 25835 59075
rect 25777 59035 25835 59041
rect 37550 59032 37556 59084
rect 37608 59072 37614 59084
rect 37645 59075 37703 59081
rect 37645 59072 37657 59075
rect 37608 59044 37657 59072
rect 37608 59032 37614 59044
rect 37645 59041 37657 59044
rect 37691 59041 37703 59075
rect 37645 59035 37703 59041
rect 4893 59007 4951 59013
rect 4893 58973 4905 59007
rect 4939 59004 4951 59007
rect 6178 59004 6184 59016
rect 4939 58976 6184 59004
rect 4939 58973 4951 58976
rect 4893 58967 4951 58973
rect 6178 58964 6184 58976
rect 6236 58964 6242 59016
rect 6733 59007 6791 59013
rect 6733 58973 6745 59007
rect 6779 59004 6791 59007
rect 6822 59004 6828 59016
rect 6779 58976 6828 59004
rect 6779 58973 6791 58976
rect 6733 58967 6791 58973
rect 6822 58964 6828 58976
rect 6880 58964 6886 59016
rect 8202 58964 8208 59016
rect 8260 59004 8266 59016
rect 8941 59007 8999 59013
rect 8941 59004 8953 59007
rect 8260 58976 8953 59004
rect 8260 58964 8266 58976
rect 8941 58973 8953 58976
rect 8987 58973 8999 59007
rect 8941 58967 8999 58973
rect 9208 59007 9266 59013
rect 9208 58973 9220 59007
rect 9254 59004 9266 59007
rect 9582 59004 9588 59016
rect 9254 58976 9588 59004
rect 9254 58973 9266 58976
rect 9208 58967 9266 58973
rect 9582 58964 9588 58976
rect 9640 58964 9646 59016
rect 10781 59007 10839 59013
rect 10781 58973 10793 59007
rect 10827 59004 10839 59007
rect 11514 59004 11520 59016
rect 10827 58976 11520 59004
rect 10827 58973 10839 58976
rect 10781 58967 10839 58973
rect 11514 58964 11520 58976
rect 11572 58964 11578 59016
rect 14090 59004 14096 59016
rect 14051 58976 14096 59004
rect 14090 58964 14096 58976
rect 14148 58964 14154 59016
rect 14360 59007 14418 59013
rect 14360 58973 14372 59007
rect 14406 59004 14418 59007
rect 14734 59004 14740 59016
rect 14406 58976 14740 59004
rect 14406 58973 14418 58976
rect 14360 58967 14418 58973
rect 14734 58964 14740 58976
rect 14792 58964 14798 59016
rect 15930 59004 15936 59016
rect 15891 58976 15936 59004
rect 15930 58964 15936 58976
rect 15988 58964 15994 59016
rect 19978 58964 19984 59016
rect 20036 59004 20042 59016
rect 20533 59007 20591 59013
rect 20533 59004 20545 59007
rect 20036 58976 20545 59004
rect 20036 58964 20042 58976
rect 20533 58973 20545 58976
rect 20579 59004 20591 59007
rect 22465 59007 22523 59013
rect 22465 59004 22477 59007
rect 20579 58976 22477 59004
rect 20579 58973 20591 58976
rect 20533 58967 20591 58973
rect 22465 58973 22477 58976
rect 22511 58973 22523 59007
rect 22465 58967 22523 58973
rect 26044 59007 26102 59013
rect 26044 58973 26056 59007
rect 26090 59004 26102 59007
rect 27246 59004 27252 59016
rect 26090 58976 27252 59004
rect 26090 58973 26102 58976
rect 26044 58967 26102 58973
rect 27246 58964 27252 58976
rect 27304 58964 27310 59016
rect 27522 58964 27528 59016
rect 27580 59004 27586 59016
rect 27617 59007 27675 59013
rect 27617 59004 27629 59007
rect 27580 58976 27629 59004
rect 27580 58964 27586 58976
rect 27617 58973 27629 58976
rect 27663 58973 27675 59007
rect 27617 58967 27675 58973
rect 27884 59007 27942 59013
rect 27884 58973 27896 59007
rect 27930 59004 27942 59007
rect 29362 59004 29368 59016
rect 27930 58976 29368 59004
rect 27930 58973 27942 58976
rect 27884 58967 27942 58973
rect 29362 58964 29368 58976
rect 29420 58964 29426 59016
rect 30282 59004 30288 59016
rect 30243 58976 30288 59004
rect 30282 58964 30288 58976
rect 30340 58964 30346 59016
rect 32125 59007 32183 59013
rect 32125 58973 32137 59007
rect 32171 59004 32183 59007
rect 32858 59004 32864 59016
rect 32171 58976 32864 59004
rect 32171 58973 32183 58976
rect 32125 58967 32183 58973
rect 32858 58964 32864 58976
rect 32916 58964 32922 59016
rect 34514 58964 34520 59016
rect 34572 59004 34578 59016
rect 35342 59004 35348 59016
rect 34572 58976 35348 59004
rect 34572 58964 34578 58976
rect 35342 58964 35348 58976
rect 35400 59004 35406 59016
rect 35621 59007 35679 59013
rect 35621 59004 35633 59007
rect 35400 58976 35633 59004
rect 35400 58964 35406 58976
rect 35621 58973 35633 58976
rect 35667 58973 35679 59007
rect 35621 58967 35679 58973
rect 35888 59007 35946 59013
rect 35888 58973 35900 59007
rect 35934 59004 35946 59007
rect 36722 59004 36728 59016
rect 35934 58976 36728 59004
rect 35934 58973 35946 58976
rect 35888 58967 35946 58973
rect 36722 58964 36728 58976
rect 36780 58964 36786 59016
rect 41233 59007 41291 59013
rect 41233 58973 41245 59007
rect 41279 59004 41291 59007
rect 42794 59004 42800 59016
rect 41279 58976 42800 59004
rect 41279 58973 41291 58976
rect 41233 58967 41291 58973
rect 42794 58964 42800 58976
rect 42852 59004 42858 59016
rect 43073 59007 43131 59013
rect 43073 59004 43085 59007
rect 42852 58976 43085 59004
rect 42852 58964 42858 58976
rect 43073 58973 43085 58976
rect 43119 58973 43131 59007
rect 43073 58967 43131 58973
rect 46385 59007 46443 59013
rect 46385 58973 46397 59007
rect 46431 59004 46443 59007
rect 48225 59007 48283 59013
rect 48225 59004 48237 59007
rect 46431 58976 48237 59004
rect 46431 58973 46443 58976
rect 46385 58967 46443 58973
rect 48225 58973 48237 58976
rect 48271 59004 48283 59007
rect 48958 59004 48964 59016
rect 48271 58976 48964 59004
rect 48271 58973 48283 58976
rect 48225 58967 48283 58973
rect 48958 58964 48964 58976
rect 49016 58964 49022 59016
rect 50798 58964 50804 59016
rect 50856 59004 50862 59016
rect 51537 59007 51595 59013
rect 51537 59004 51549 59007
rect 50856 58976 51549 59004
rect 50856 58964 50862 58976
rect 51537 58973 51549 58976
rect 51583 58973 51595 59007
rect 51537 58967 51595 58973
rect 51804 59007 51862 59013
rect 51804 58973 51816 59007
rect 51850 59004 51862 59007
rect 53190 59004 53196 59016
rect 51850 58976 53196 59004
rect 51850 58973 51862 58976
rect 51804 58967 51862 58973
rect 53190 58964 53196 58976
rect 53248 58964 53254 59016
rect 53374 59004 53380 59016
rect 53335 58976 53380 59004
rect 53374 58964 53380 58976
rect 53432 59004 53438 59016
rect 55309 59007 55367 59013
rect 55309 59004 55321 59007
rect 53432 58976 55321 59004
rect 53432 58964 53438 58976
rect 55309 58973 55321 58976
rect 55355 58973 55367 59007
rect 55309 58967 55367 58973
rect 55398 58964 55404 59016
rect 55456 59004 55462 59016
rect 55565 59007 55623 59013
rect 55565 59004 55577 59007
rect 55456 58976 55577 59004
rect 55456 58964 55462 58976
rect 55565 58973 55577 58976
rect 55611 58973 55623 59007
rect 55565 58967 55623 58973
rect 57054 58964 57060 59016
rect 57112 59004 57118 59016
rect 57241 59007 57299 59013
rect 57241 59004 57253 59007
rect 57112 58976 57253 59004
rect 57112 58964 57118 58976
rect 57241 58973 57253 58976
rect 57287 58973 57299 59007
rect 57241 58967 57299 58973
rect 5160 58939 5218 58945
rect 5160 58905 5172 58939
rect 5206 58936 5218 58939
rect 5994 58936 6000 58948
rect 5206 58908 6000 58936
rect 5206 58905 5218 58908
rect 5160 58899 5218 58905
rect 5994 58896 6000 58908
rect 6052 58896 6058 58948
rect 7000 58939 7058 58945
rect 7000 58905 7012 58939
rect 7046 58936 7058 58939
rect 7742 58936 7748 58948
rect 7046 58908 7748 58936
rect 7046 58905 7058 58908
rect 7000 58899 7058 58905
rect 7742 58896 7748 58908
rect 7800 58896 7806 58948
rect 11048 58939 11106 58945
rect 11048 58905 11060 58939
rect 11094 58936 11106 58939
rect 12802 58936 12808 58948
rect 11094 58908 12808 58936
rect 11094 58905 11106 58908
rect 11048 58899 11106 58905
rect 12802 58896 12808 58908
rect 12860 58896 12866 58948
rect 15838 58896 15844 58948
rect 15896 58936 15902 58948
rect 16178 58939 16236 58945
rect 16178 58936 16190 58939
rect 15896 58908 16190 58936
rect 15896 58896 15902 58908
rect 16178 58905 16190 58908
rect 16224 58905 16236 58939
rect 16178 58899 16236 58905
rect 20800 58939 20858 58945
rect 20800 58905 20812 58939
rect 20846 58936 20858 58939
rect 21266 58936 21272 58948
rect 20846 58908 21272 58936
rect 20846 58905 20858 58908
rect 20800 58899 20858 58905
rect 21266 58896 21272 58908
rect 21324 58896 21330 58948
rect 22732 58939 22790 58945
rect 22732 58905 22744 58939
rect 22778 58936 22790 58939
rect 23842 58936 23848 58948
rect 22778 58908 23848 58936
rect 22778 58905 22790 58908
rect 22732 58899 22790 58905
rect 23842 58896 23848 58908
rect 23900 58896 23906 58948
rect 30552 58939 30610 58945
rect 30552 58905 30564 58939
rect 30598 58936 30610 58939
rect 30598 58908 31800 58936
rect 30598 58905 30610 58908
rect 30552 58899 30610 58905
rect 6270 58868 6276 58880
rect 6231 58840 6276 58868
rect 6270 58828 6276 58840
rect 6328 58828 6334 58880
rect 10318 58868 10324 58880
rect 10279 58840 10324 58868
rect 10318 58828 10324 58840
rect 10376 58828 10382 58880
rect 12158 58868 12164 58880
rect 12119 58840 12164 58868
rect 12158 58828 12164 58840
rect 12216 58828 12222 58880
rect 15470 58868 15476 58880
rect 15431 58840 15476 58868
rect 15470 58828 15476 58840
rect 15528 58828 15534 58880
rect 17310 58868 17316 58880
rect 17271 58840 17316 58868
rect 17310 58828 17316 58840
rect 17368 58828 17374 58880
rect 21910 58868 21916 58880
rect 21871 58840 21916 58868
rect 21910 58828 21916 58840
rect 21968 58828 21974 58880
rect 27154 58868 27160 58880
rect 27115 58840 27160 58868
rect 27154 58828 27160 58840
rect 27212 58828 27218 58880
rect 28994 58868 29000 58880
rect 28955 58840 29000 58868
rect 28994 58828 29000 58840
rect 29052 58828 29058 58880
rect 31662 58868 31668 58880
rect 31623 58840 31668 58868
rect 31662 58828 31668 58840
rect 31720 58828 31726 58880
rect 31772 58868 31800 58908
rect 31846 58896 31852 58948
rect 31904 58936 31910 58948
rect 32370 58939 32428 58945
rect 32370 58936 32382 58939
rect 31904 58908 32382 58936
rect 31904 58896 31910 58908
rect 32370 58905 32382 58908
rect 32416 58905 32428 58939
rect 32370 58899 32428 58905
rect 37912 58939 37970 58945
rect 37912 58905 37924 58939
rect 37958 58936 37970 58939
rect 38838 58936 38844 58948
rect 37958 58908 38844 58936
rect 37958 58905 37970 58908
rect 37912 58899 37970 58905
rect 38838 58896 38844 58908
rect 38896 58896 38902 58948
rect 41500 58939 41558 58945
rect 41500 58905 41512 58939
rect 41546 58936 41558 58939
rect 43162 58936 43168 58948
rect 41546 58908 43168 58936
rect 41546 58905 41558 58908
rect 41500 58899 41558 58905
rect 43162 58896 43168 58908
rect 43220 58896 43226 58948
rect 43340 58939 43398 58945
rect 43340 58905 43352 58939
rect 43386 58936 43398 58939
rect 45186 58936 45192 58948
rect 43386 58908 45192 58936
rect 43386 58905 43398 58908
rect 43340 58899 43398 58905
rect 45186 58896 45192 58908
rect 45244 58896 45250 58948
rect 46652 58939 46710 58945
rect 46652 58905 46664 58939
rect 46698 58936 46710 58939
rect 47302 58936 47308 58948
rect 46698 58908 47308 58936
rect 46698 58905 46710 58908
rect 46652 58899 46710 58905
rect 47302 58896 47308 58908
rect 47360 58896 47366 58948
rect 48492 58939 48550 58945
rect 48492 58905 48504 58939
rect 48538 58936 48550 58939
rect 49418 58936 49424 58948
rect 48538 58908 49424 58936
rect 48538 58905 48550 58908
rect 48492 58899 48550 58905
rect 49418 58896 49424 58908
rect 49476 58896 49482 58948
rect 53644 58939 53702 58945
rect 53644 58905 53656 58939
rect 53690 58936 53702 58939
rect 54754 58936 54760 58948
rect 53690 58908 54760 58936
rect 53690 58905 53702 58908
rect 53644 58899 53702 58905
rect 54754 58896 54760 58908
rect 54812 58896 54818 58948
rect 56778 58896 56784 58948
rect 56836 58936 56842 58948
rect 57486 58939 57544 58945
rect 57486 58936 57498 58939
rect 56836 58908 57498 58936
rect 56836 58896 56842 58908
rect 57486 58905 57498 58908
rect 57532 58905 57544 58939
rect 57486 58899 57544 58905
rect 33505 58871 33563 58877
rect 33505 58868 33517 58871
rect 31772 58840 33517 58868
rect 33505 58837 33517 58840
rect 33551 58837 33563 58871
rect 36998 58868 37004 58880
rect 36959 58840 37004 58868
rect 33505 58831 33563 58837
rect 36998 58828 37004 58840
rect 37056 58828 37062 58880
rect 42610 58868 42616 58880
rect 42571 58840 42616 58868
rect 42610 58828 42616 58840
rect 42668 58828 42674 58880
rect 47762 58868 47768 58880
rect 47723 58840 47768 58868
rect 47762 58828 47768 58840
rect 47820 58828 47826 58880
rect 48314 58828 48320 58880
rect 48372 58868 48378 58880
rect 49605 58871 49663 58877
rect 49605 58868 49617 58871
rect 48372 58840 49617 58868
rect 48372 58828 48378 58840
rect 49605 58837 49617 58840
rect 49651 58837 49663 58871
rect 49605 58831 49663 58837
rect 52546 58828 52552 58880
rect 52604 58868 52610 58880
rect 52917 58871 52975 58877
rect 52917 58868 52929 58871
rect 52604 58840 52929 58868
rect 52604 58828 52610 58840
rect 52917 58837 52929 58840
rect 52963 58837 52975 58871
rect 58618 58868 58624 58880
rect 58579 58840 58624 58868
rect 52917 58831 52975 58837
rect 58618 58828 58624 58840
rect 58676 58828 58682 58880
rect 1104 58778 59340 58800
rect 1104 58726 19574 58778
rect 19626 58726 19638 58778
rect 19690 58726 19702 58778
rect 19754 58726 19766 58778
rect 19818 58726 19830 58778
rect 19882 58726 50294 58778
rect 50346 58726 50358 58778
rect 50410 58726 50422 58778
rect 50474 58726 50486 58778
rect 50538 58726 50550 58778
rect 50602 58726 59340 58778
rect 1104 58704 59340 58726
rect 7742 58664 7748 58676
rect 7703 58636 7748 58664
rect 7742 58624 7748 58636
rect 7800 58624 7806 58676
rect 9490 58624 9496 58676
rect 9548 58664 9554 58676
rect 9585 58667 9643 58673
rect 9585 58664 9597 58667
rect 9548 58636 9597 58664
rect 9548 58624 9554 58636
rect 9585 58633 9597 58636
rect 9631 58633 9643 58667
rect 9585 58627 9643 58633
rect 14642 58624 14648 58676
rect 14700 58664 14706 58676
rect 14737 58667 14795 58673
rect 14737 58664 14749 58667
rect 14700 58636 14749 58664
rect 14700 58624 14706 58636
rect 14737 58633 14749 58636
rect 14783 58633 14795 58667
rect 14737 58627 14795 58633
rect 21174 58624 21180 58676
rect 21232 58664 21238 58676
rect 21269 58667 21327 58673
rect 21269 58664 21281 58667
rect 21232 58636 21281 58664
rect 21232 58624 21238 58636
rect 21269 58633 21281 58636
rect 21315 58633 21327 58667
rect 25958 58664 25964 58676
rect 25919 58636 25964 58664
rect 21269 58627 21327 58633
rect 25958 58624 25964 58636
rect 26016 58624 26022 58676
rect 31573 58667 31631 58673
rect 31573 58633 31585 58667
rect 31619 58664 31631 58667
rect 31754 58664 31760 58676
rect 31619 58636 31760 58664
rect 31619 58633 31631 58636
rect 31573 58627 31631 58633
rect 31754 58624 31760 58636
rect 31812 58624 31818 58676
rect 38838 58664 38844 58676
rect 38799 58636 38844 58664
rect 38838 58624 38844 58636
rect 38896 58624 38902 58676
rect 41874 58664 41880 58676
rect 41835 58636 41880 58664
rect 41874 58624 41880 58636
rect 41932 58624 41938 58676
rect 45186 58664 45192 58676
rect 45147 58636 45192 58664
rect 45186 58624 45192 58636
rect 45244 58624 45250 58676
rect 47026 58664 47032 58676
rect 46987 58636 47032 58664
rect 47026 58624 47032 58636
rect 47084 58624 47090 58676
rect 6178 58596 6184 58608
rect 4172 58568 6184 58596
rect 4172 58537 4200 58568
rect 6178 58556 6184 58568
rect 6236 58556 6242 58608
rect 6270 58556 6276 58608
rect 6328 58596 6334 58608
rect 8478 58605 8484 58608
rect 6610 58599 6668 58605
rect 6610 58596 6622 58599
rect 6328 58568 6622 58596
rect 6328 58556 6334 58568
rect 6610 58565 6622 58568
rect 6656 58565 6668 58599
rect 8472 58596 8484 58605
rect 8439 58568 8484 58596
rect 6610 58559 6668 58565
rect 8472 58559 8484 58568
rect 8478 58556 8484 58559
rect 8536 58556 8542 58608
rect 11784 58599 11842 58605
rect 11784 58565 11796 58599
rect 11830 58596 11842 58599
rect 12158 58596 12164 58608
rect 11830 58568 12164 58596
rect 11830 58565 11842 58568
rect 11784 58559 11842 58565
rect 12158 58556 12164 58568
rect 12216 58556 12222 58608
rect 13078 58556 13084 58608
rect 13136 58596 13142 58608
rect 13602 58599 13660 58605
rect 13602 58596 13614 58599
rect 13136 58568 13614 58596
rect 13136 58556 13142 58568
rect 13602 58565 13614 58568
rect 13648 58565 13660 58599
rect 13602 58559 13660 58565
rect 20156 58599 20214 58605
rect 20156 58565 20168 58599
rect 20202 58596 20214 58599
rect 21910 58596 21916 58608
rect 20202 58568 21916 58596
rect 20202 58565 20214 58568
rect 20156 58559 20214 58565
rect 21910 58556 21916 58568
rect 21968 58556 21974 58608
rect 23008 58599 23066 58605
rect 23008 58565 23020 58599
rect 23054 58596 23066 58599
rect 23934 58596 23940 58608
rect 23054 58568 23940 58596
rect 23054 58565 23066 58568
rect 23008 58559 23066 58565
rect 23934 58556 23940 58568
rect 23992 58556 23998 58608
rect 28160 58599 28218 58605
rect 28160 58565 28172 58599
rect 28206 58596 28218 58599
rect 28994 58596 29000 58608
rect 28206 58568 29000 58596
rect 28206 58565 28218 58568
rect 28160 58559 28218 58565
rect 28994 58556 29000 58568
rect 29052 58556 29058 58608
rect 30460 58599 30518 58605
rect 30460 58565 30472 58599
rect 30506 58596 30518 58599
rect 31662 58596 31668 58608
rect 30506 58568 31668 58596
rect 30506 58565 30518 58568
rect 30460 58559 30518 58565
rect 31662 58556 31668 58568
rect 31720 58556 31726 58608
rect 33873 58599 33931 58605
rect 33873 58565 33885 58599
rect 33919 58596 33931 58599
rect 39022 58596 39028 58608
rect 33919 58568 39028 58596
rect 33919 58565 33931 58568
rect 33873 58559 33931 58565
rect 39022 58556 39028 58568
rect 39080 58556 39086 58608
rect 40764 58599 40822 58605
rect 40764 58565 40776 58599
rect 40810 58596 40822 58599
rect 42610 58596 42616 58608
rect 40810 58568 42616 58596
rect 40810 58565 40822 58568
rect 40764 58559 40822 58565
rect 42610 58556 42616 58568
rect 42668 58556 42674 58608
rect 44076 58599 44134 58605
rect 44076 58565 44088 58599
rect 44122 58596 44134 58599
rect 44174 58596 44180 58608
rect 44122 58568 44180 58596
rect 44122 58565 44134 58568
rect 44076 58559 44134 58565
rect 44174 58556 44180 58568
rect 44232 58556 44238 58608
rect 45916 58599 45974 58605
rect 45916 58565 45928 58599
rect 45962 58596 45974 58599
rect 47762 58596 47768 58608
rect 45962 58568 47768 58596
rect 45962 58565 45974 58568
rect 45916 58559 45974 58565
rect 47762 58556 47768 58568
rect 47820 58556 47826 58608
rect 53098 58596 53104 58608
rect 47964 58568 53104 58596
rect 4157 58531 4215 58537
rect 4157 58497 4169 58531
rect 4203 58497 4215 58531
rect 4157 58491 4215 58497
rect 4424 58531 4482 58537
rect 4424 58497 4436 58531
rect 4470 58528 4482 58531
rect 5166 58528 5172 58540
rect 4470 58500 5172 58528
rect 4470 58497 4482 58500
rect 4424 58491 4482 58497
rect 5166 58488 5172 58500
rect 5224 58488 5230 58540
rect 6914 58488 6920 58540
rect 6972 58528 6978 58540
rect 8202 58528 8208 58540
rect 6972 58500 8208 58528
rect 6972 58488 6978 58500
rect 8202 58488 8208 58500
rect 8260 58488 8266 58540
rect 13357 58531 13415 58537
rect 13357 58528 13369 58531
rect 11532 58500 13369 58528
rect 11532 58472 11560 58500
rect 13357 58497 13369 58500
rect 13403 58528 13415 58531
rect 14090 58528 14096 58540
rect 13403 58500 14096 58528
rect 13403 58497 13415 58500
rect 13357 58491 13415 58497
rect 14090 58488 14096 58500
rect 14148 58488 14154 58540
rect 18316 58531 18374 58537
rect 18316 58497 18328 58531
rect 18362 58528 18374 58531
rect 19150 58528 19156 58540
rect 18362 58500 19156 58528
rect 18362 58497 18374 58500
rect 18316 58491 18374 58497
rect 19150 58488 19156 58500
rect 19208 58488 19214 58540
rect 19889 58531 19947 58537
rect 19889 58497 19901 58531
rect 19935 58528 19947 58531
rect 19978 58528 19984 58540
rect 19935 58500 19984 58528
rect 19935 58497 19947 58500
rect 19889 58491 19947 58497
rect 19978 58488 19984 58500
rect 20036 58488 20042 58540
rect 22462 58488 22468 58540
rect 22520 58528 22526 58540
rect 22741 58531 22799 58537
rect 22741 58528 22753 58531
rect 22520 58500 22753 58528
rect 22520 58488 22526 58500
rect 22741 58497 22753 58500
rect 22787 58528 22799 58531
rect 24581 58531 24639 58537
rect 24581 58528 24593 58531
rect 22787 58500 24593 58528
rect 22787 58497 22799 58500
rect 22741 58491 22799 58497
rect 24581 58497 24593 58500
rect 24627 58497 24639 58531
rect 24581 58491 24639 58497
rect 24848 58531 24906 58537
rect 24848 58497 24860 58531
rect 24894 58528 24906 58531
rect 26418 58528 26424 58540
rect 24894 58500 26424 58528
rect 24894 58497 24906 58500
rect 24848 58491 24906 58497
rect 26418 58488 26424 58500
rect 26476 58488 26482 58540
rect 30193 58531 30251 58537
rect 30193 58497 30205 58531
rect 30239 58528 30251 58531
rect 30282 58528 30288 58540
rect 30239 58500 30288 58528
rect 30239 58497 30251 58500
rect 30193 58491 30251 58497
rect 30282 58488 30288 58500
rect 30340 58488 30346 58540
rect 37274 58488 37280 58540
rect 37332 58528 37338 58540
rect 37461 58531 37519 58537
rect 37461 58528 37473 58531
rect 37332 58500 37473 58528
rect 37332 58488 37338 58500
rect 37461 58497 37473 58500
rect 37507 58528 37519 58531
rect 37550 58528 37556 58540
rect 37507 58500 37556 58528
rect 37507 58497 37519 58500
rect 37461 58491 37519 58497
rect 37550 58488 37556 58500
rect 37608 58488 37614 58540
rect 37728 58531 37786 58537
rect 37728 58497 37740 58531
rect 37774 58528 37786 58531
rect 38562 58528 38568 58540
rect 37774 58500 38568 58528
rect 37774 58497 37786 58500
rect 37728 58491 37786 58497
rect 38562 58488 38568 58500
rect 38620 58488 38626 58540
rect 43622 58488 43628 58540
rect 43680 58528 43686 58540
rect 43809 58531 43867 58537
rect 43809 58528 43821 58531
rect 43680 58500 43821 58528
rect 43680 58488 43686 58500
rect 43809 58497 43821 58500
rect 43855 58497 43867 58531
rect 43809 58491 43867 58497
rect 45554 58488 45560 58540
rect 45612 58528 45618 58540
rect 45649 58531 45707 58537
rect 45649 58528 45661 58531
rect 45612 58500 45661 58528
rect 45612 58488 45618 58500
rect 45649 58497 45661 58500
rect 45695 58497 45707 58531
rect 45649 58491 45707 58497
rect 47118 58488 47124 58540
rect 47176 58528 47182 58540
rect 47964 58537 47992 58568
rect 53098 58556 53104 58568
rect 53156 58556 53162 58608
rect 54380 58599 54438 58605
rect 54380 58565 54392 58599
rect 54426 58596 54438 58599
rect 55950 58596 55956 58608
rect 54426 58568 55956 58596
rect 54426 58565 54438 58568
rect 54380 58559 54438 58565
rect 55950 58556 55956 58568
rect 56008 58556 56014 58608
rect 56220 58599 56278 58605
rect 56220 58565 56232 58599
rect 56266 58596 56278 58599
rect 58618 58596 58624 58608
rect 56266 58568 58624 58596
rect 56266 58565 56278 58568
rect 56220 58559 56278 58565
rect 58618 58556 58624 58568
rect 58676 58556 58682 58608
rect 47949 58531 48007 58537
rect 47949 58528 47961 58531
rect 47176 58500 47961 58528
rect 47176 58488 47182 58500
rect 47949 58497 47961 58500
rect 47995 58497 48007 58531
rect 47949 58491 48007 58497
rect 51068 58531 51126 58537
rect 51068 58497 51080 58531
rect 51114 58528 51126 58531
rect 52914 58528 52920 58540
rect 51114 58500 52920 58528
rect 51114 58497 51126 58500
rect 51068 58491 51126 58497
rect 52914 58488 52920 58500
rect 52972 58488 52978 58540
rect 54110 58528 54116 58540
rect 54071 58500 54116 58528
rect 54110 58488 54116 58500
rect 54168 58528 54174 58540
rect 55214 58528 55220 58540
rect 54168 58500 55220 58528
rect 54168 58488 54174 58500
rect 55214 58488 55220 58500
rect 55272 58528 55278 58540
rect 55858 58528 55864 58540
rect 55272 58500 55864 58528
rect 55272 58488 55278 58500
rect 55858 58488 55864 58500
rect 55916 58528 55922 58540
rect 57054 58528 57060 58540
rect 55916 58500 57060 58528
rect 55916 58488 55922 58500
rect 6270 58420 6276 58472
rect 6328 58460 6334 58472
rect 6365 58463 6423 58469
rect 6365 58460 6377 58463
rect 6328 58432 6377 58460
rect 6328 58420 6334 58432
rect 6365 58429 6377 58432
rect 6411 58429 6423 58463
rect 11514 58460 11520 58472
rect 11475 58432 11520 58460
rect 6365 58423 6423 58429
rect 11514 58420 11520 58432
rect 11572 58420 11578 58472
rect 18046 58460 18052 58472
rect 18007 58432 18052 58460
rect 18046 58420 18052 58432
rect 18104 58420 18110 58472
rect 27522 58420 27528 58472
rect 27580 58460 27586 58472
rect 27893 58463 27951 58469
rect 27893 58460 27905 58463
rect 27580 58432 27905 58460
rect 27580 58420 27586 58432
rect 27893 58429 27905 58432
rect 27939 58429 27951 58463
rect 27893 58423 27951 58429
rect 40402 58420 40408 58472
rect 40460 58460 40466 58472
rect 40497 58463 40555 58469
rect 40497 58460 40509 58463
rect 40460 58432 40509 58460
rect 40460 58420 40466 58432
rect 40497 58429 40509 58432
rect 40543 58429 40555 58463
rect 50798 58460 50804 58472
rect 50759 58432 50804 58460
rect 40497 58423 40555 58429
rect 50798 58420 50804 58432
rect 50856 58420 50862 58472
rect 55968 58469 55996 58500
rect 57054 58488 57060 58500
rect 57112 58488 57118 58540
rect 55953 58463 56011 58469
rect 55953 58429 55965 58463
rect 55999 58429 56011 58463
rect 55953 58423 56011 58429
rect 5534 58324 5540 58336
rect 5495 58296 5540 58324
rect 5534 58284 5540 58296
rect 5592 58284 5598 58336
rect 12894 58324 12900 58336
rect 12855 58296 12900 58324
rect 12894 58284 12900 58296
rect 12952 58284 12958 58336
rect 19334 58284 19340 58336
rect 19392 58324 19398 58336
rect 19429 58327 19487 58333
rect 19429 58324 19441 58327
rect 19392 58296 19441 58324
rect 19392 58284 19398 58296
rect 19429 58293 19441 58296
rect 19475 58293 19487 58327
rect 24118 58324 24124 58336
rect 24079 58296 24124 58324
rect 19429 58287 19487 58293
rect 24118 58284 24124 58296
rect 24176 58284 24182 58336
rect 29270 58324 29276 58336
rect 29231 58296 29276 58324
rect 29270 58284 29276 58296
rect 29328 58284 29334 58336
rect 35342 58324 35348 58336
rect 35303 58296 35348 58324
rect 35342 58284 35348 58296
rect 35400 58284 35406 58336
rect 48958 58284 48964 58336
rect 49016 58324 49022 58336
rect 49237 58327 49295 58333
rect 49237 58324 49249 58327
rect 49016 58296 49249 58324
rect 49016 58284 49022 58296
rect 49237 58293 49249 58296
rect 49283 58293 49295 58327
rect 52178 58324 52184 58336
rect 52139 58296 52184 58324
rect 49237 58287 49295 58293
rect 52178 58284 52184 58296
rect 52236 58284 52242 58336
rect 54386 58284 54392 58336
rect 54444 58324 54450 58336
rect 55493 58327 55551 58333
rect 55493 58324 55505 58327
rect 54444 58296 55505 58324
rect 54444 58284 54450 58296
rect 55493 58293 55505 58296
rect 55539 58293 55551 58327
rect 55493 58287 55551 58293
rect 56870 58284 56876 58336
rect 56928 58324 56934 58336
rect 57333 58327 57391 58333
rect 57333 58324 57345 58327
rect 56928 58296 57345 58324
rect 56928 58284 56934 58296
rect 57333 58293 57345 58296
rect 57379 58293 57391 58327
rect 57333 58287 57391 58293
rect 1104 58234 59340 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 34934 58234
rect 34986 58182 34998 58234
rect 35050 58182 35062 58234
rect 35114 58182 35126 58234
rect 35178 58182 35190 58234
rect 35242 58182 59340 58234
rect 1104 58160 59340 58182
rect 5166 58120 5172 58132
rect 5127 58092 5172 58120
rect 5166 58080 5172 58092
rect 5224 58080 5230 58132
rect 38562 58120 38568 58132
rect 38523 58092 38568 58120
rect 38562 58080 38568 58092
rect 38620 58080 38626 58132
rect 47302 58080 47308 58132
rect 47360 58120 47366 58132
rect 47765 58123 47823 58129
rect 47765 58120 47777 58123
rect 47360 58092 47777 58120
rect 47360 58080 47366 58092
rect 47765 58089 47777 58092
rect 47811 58089 47823 58123
rect 48958 58120 48964 58132
rect 47765 58083 47823 58089
rect 48240 58092 48964 58120
rect 10321 58055 10379 58061
rect 10321 58021 10333 58055
rect 10367 58021 10379 58055
rect 10321 58015 10379 58021
rect 10336 57984 10364 58015
rect 19978 58012 19984 58064
rect 20036 58052 20042 58064
rect 21729 58055 21787 58061
rect 21729 58052 21741 58055
rect 20036 58024 21741 58052
rect 20036 58012 20042 58024
rect 21729 58021 21741 58024
rect 21775 58021 21787 58055
rect 21729 58015 21787 58021
rect 10336 57956 10456 57984
rect 3789 57919 3847 57925
rect 3789 57885 3801 57919
rect 3835 57916 3847 57919
rect 3878 57916 3884 57928
rect 3835 57888 3884 57916
rect 3835 57885 3847 57888
rect 3789 57879 3847 57885
rect 3878 57876 3884 57888
rect 3936 57876 3942 57928
rect 5629 57919 5687 57925
rect 5629 57885 5641 57919
rect 5675 57916 5687 57919
rect 6914 57916 6920 57928
rect 5675 57888 6920 57916
rect 5675 57885 5687 57888
rect 5629 57879 5687 57885
rect 6914 57876 6920 57888
rect 6972 57876 6978 57928
rect 8941 57919 8999 57925
rect 8941 57885 8953 57919
rect 8987 57885 8999 57919
rect 8941 57879 8999 57885
rect 9208 57919 9266 57925
rect 9208 57885 9220 57919
rect 9254 57916 9266 57919
rect 10318 57916 10324 57928
rect 9254 57888 10324 57916
rect 9254 57885 9266 57888
rect 9208 57879 9266 57885
rect 4056 57851 4114 57857
rect 4056 57817 4068 57851
rect 4102 57848 4114 57851
rect 4982 57848 4988 57860
rect 4102 57820 4988 57848
rect 4102 57817 4114 57820
rect 4056 57811 4114 57817
rect 4982 57808 4988 57820
rect 5040 57808 5046 57860
rect 5534 57808 5540 57860
rect 5592 57848 5598 57860
rect 5874 57851 5932 57857
rect 5874 57848 5886 57851
rect 5592 57820 5886 57848
rect 5592 57808 5598 57820
rect 5874 57817 5886 57820
rect 5920 57817 5932 57851
rect 5874 57811 5932 57817
rect 8956 57792 8984 57879
rect 10318 57876 10324 57888
rect 10376 57876 10382 57928
rect 10428 57848 10456 57956
rect 15930 57944 15936 57996
rect 15988 57984 15994 57996
rect 40402 57984 40408 57996
rect 15988 57956 17356 57984
rect 40363 57956 40408 57984
rect 15988 57944 15994 57956
rect 10778 57916 10784 57928
rect 10739 57888 10784 57916
rect 10778 57876 10784 57888
rect 10836 57876 10842 57928
rect 17328 57925 17356 57956
rect 40402 57944 40408 57956
rect 40460 57944 40466 57996
rect 48240 57993 48268 58092
rect 48958 58080 48964 58092
rect 49016 58080 49022 58132
rect 52914 58120 52920 58132
rect 52875 58092 52920 58120
rect 52914 58080 52920 58092
rect 52972 58080 52978 58132
rect 54754 58120 54760 58132
rect 54715 58092 54760 58120
rect 54754 58080 54760 58092
rect 54812 58080 54818 58132
rect 48225 57987 48283 57993
rect 48225 57953 48237 57987
rect 48271 57953 48283 57987
rect 48225 57947 48283 57953
rect 17313 57919 17371 57925
rect 17313 57885 17325 57919
rect 17359 57916 17371 57919
rect 18046 57916 18052 57928
rect 17359 57888 18052 57916
rect 17359 57885 17371 57888
rect 17313 57879 17371 57885
rect 18046 57876 18052 57888
rect 18104 57876 18110 57928
rect 25038 57876 25044 57928
rect 25096 57916 25102 57928
rect 25777 57919 25835 57925
rect 25777 57916 25789 57919
rect 25096 57888 25789 57916
rect 25096 57876 25102 57888
rect 25777 57885 25789 57888
rect 25823 57885 25835 57919
rect 25777 57879 25835 57885
rect 27522 57876 27528 57928
rect 27580 57916 27586 57928
rect 27617 57919 27675 57925
rect 27617 57916 27629 57919
rect 27580 57888 27629 57916
rect 27580 57876 27586 57888
rect 27617 57885 27629 57888
rect 27663 57885 27675 57919
rect 27617 57879 27675 57885
rect 27884 57919 27942 57925
rect 27884 57885 27896 57919
rect 27930 57916 27942 57919
rect 29270 57916 29276 57928
rect 27930 57888 29276 57916
rect 27930 57885 27942 57888
rect 27884 57879 27942 57885
rect 29270 57876 29276 57888
rect 29328 57876 29334 57928
rect 30282 57876 30288 57928
rect 30340 57916 30346 57928
rect 30929 57919 30987 57925
rect 30929 57916 30941 57919
rect 30340 57888 30941 57916
rect 30340 57876 30346 57888
rect 30929 57885 30941 57888
rect 30975 57916 30987 57919
rect 32769 57919 32827 57925
rect 32769 57916 32781 57919
rect 30975 57888 32781 57916
rect 30975 57885 30987 57888
rect 30929 57879 30987 57885
rect 32769 57885 32781 57888
rect 32815 57916 32827 57919
rect 32858 57916 32864 57928
rect 32815 57888 32864 57916
rect 32815 57885 32827 57888
rect 32769 57879 32827 57885
rect 32858 57876 32864 57888
rect 32916 57876 32922 57928
rect 33036 57919 33094 57925
rect 33036 57885 33048 57919
rect 33082 57916 33094 57919
rect 34606 57916 34612 57928
rect 33082 57888 34612 57916
rect 33082 57885 33094 57888
rect 33036 57879 33094 57885
rect 34606 57876 34612 57888
rect 34664 57876 34670 57928
rect 34698 57876 34704 57928
rect 34756 57916 34762 57928
rect 35342 57916 35348 57928
rect 34756 57888 35348 57916
rect 34756 57876 34762 57888
rect 35342 57876 35348 57888
rect 35400 57876 35406 57928
rect 35612 57919 35670 57925
rect 35612 57885 35624 57919
rect 35658 57916 35670 57919
rect 36998 57916 37004 57928
rect 35658 57888 37004 57916
rect 35658 57885 35670 57888
rect 35612 57879 35670 57885
rect 36998 57876 37004 57888
rect 37056 57876 37062 57928
rect 37185 57919 37243 57925
rect 37185 57885 37197 57919
rect 37231 57916 37243 57919
rect 37274 57916 37280 57928
rect 37231 57888 37280 57916
rect 37231 57885 37243 57888
rect 37185 57879 37243 57885
rect 37274 57876 37280 57888
rect 37332 57876 37338 57928
rect 40678 57925 40684 57928
rect 40672 57916 40684 57925
rect 40639 57888 40684 57916
rect 40672 57879 40684 57888
rect 40678 57876 40684 57879
rect 40736 57876 40742 57928
rect 43346 57925 43352 57928
rect 43073 57919 43131 57925
rect 43073 57885 43085 57919
rect 43119 57885 43131 57919
rect 43340 57916 43352 57925
rect 43307 57888 43352 57916
rect 43073 57879 43131 57885
rect 43340 57879 43352 57888
rect 11026 57851 11084 57857
rect 11026 57848 11038 57851
rect 10428 57820 11038 57848
rect 11026 57817 11038 57820
rect 11072 57817 11084 57851
rect 11026 57811 11084 57817
rect 13814 57808 13820 57860
rect 13872 57848 13878 57860
rect 14461 57851 14519 57857
rect 14461 57848 14473 57851
rect 13872 57820 14473 57848
rect 13872 57808 13878 57820
rect 14461 57817 14473 57820
rect 14507 57817 14519 57851
rect 14461 57811 14519 57817
rect 17580 57851 17638 57857
rect 17580 57817 17592 57851
rect 17626 57848 17638 57851
rect 18598 57848 18604 57860
rect 17626 57820 18604 57848
rect 17626 57817 17638 57820
rect 17580 57811 17638 57817
rect 18598 57808 18604 57820
rect 18656 57808 18662 57860
rect 20438 57848 20444 57860
rect 20399 57820 20444 57848
rect 20438 57808 20444 57820
rect 20496 57808 20502 57860
rect 26044 57851 26102 57857
rect 26044 57817 26056 57851
rect 26090 57848 26102 57851
rect 28902 57848 28908 57860
rect 26090 57820 28908 57848
rect 26090 57817 26102 57820
rect 26044 57811 26102 57817
rect 28902 57808 28908 57820
rect 28960 57808 28966 57860
rect 31196 57851 31254 57857
rect 31196 57817 31208 57851
rect 31242 57848 31254 57851
rect 32214 57848 32220 57860
rect 31242 57820 32220 57848
rect 31242 57817 31254 57820
rect 31196 57811 31254 57817
rect 32214 57808 32220 57820
rect 32272 57808 32278 57860
rect 37452 57851 37510 57857
rect 37452 57817 37464 57851
rect 37498 57848 37510 57851
rect 38654 57848 38660 57860
rect 37498 57820 38660 57848
rect 37498 57817 37510 57820
rect 37452 57811 37510 57817
rect 38654 57808 38660 57820
rect 38712 57808 38718 57860
rect 43088 57848 43116 57879
rect 43346 57876 43352 57879
rect 43404 57876 43410 57928
rect 46385 57919 46443 57925
rect 46385 57885 46397 57919
rect 46431 57916 46443 57919
rect 48240 57916 48268 57947
rect 48774 57916 48780 57928
rect 46431 57888 48268 57916
rect 48332 57888 48780 57916
rect 46431 57885 46443 57888
rect 46385 57879 46443 57885
rect 44266 57848 44272 57860
rect 43088 57820 44272 57848
rect 44266 57808 44272 57820
rect 44324 57848 44330 57860
rect 46400 57848 46428 57879
rect 44324 57820 46428 57848
rect 46652 57851 46710 57857
rect 44324 57808 44330 57820
rect 46652 57817 46664 57851
rect 46698 57848 46710 57851
rect 48332 57848 48360 57888
rect 48774 57876 48780 57888
rect 48832 57876 48838 57928
rect 50798 57876 50804 57928
rect 50856 57916 50862 57928
rect 51537 57919 51595 57925
rect 51537 57916 51549 57919
rect 50856 57888 51549 57916
rect 50856 57876 50862 57888
rect 51537 57885 51549 57888
rect 51583 57885 51595 57919
rect 53374 57916 53380 57928
rect 53335 57888 53380 57916
rect 51537 57879 51595 57885
rect 53374 57876 53380 57888
rect 53432 57876 53438 57928
rect 53644 57919 53702 57925
rect 53644 57885 53656 57919
rect 53690 57916 53702 57919
rect 54386 57916 54392 57928
rect 53690 57888 54392 57916
rect 53690 57885 53702 57888
rect 53644 57879 53702 57885
rect 54386 57876 54392 57888
rect 54444 57876 54450 57928
rect 55214 57876 55220 57928
rect 55272 57916 55278 57928
rect 55309 57919 55367 57925
rect 55309 57916 55321 57919
rect 55272 57888 55321 57916
rect 55272 57876 55278 57888
rect 55309 57885 55321 57888
rect 55355 57885 55367 57919
rect 55309 57879 55367 57885
rect 57054 57876 57060 57928
rect 57112 57916 57118 57928
rect 57149 57919 57207 57925
rect 57149 57916 57161 57919
rect 57112 57888 57161 57916
rect 57112 57876 57118 57888
rect 57149 57885 57161 57888
rect 57195 57885 57207 57919
rect 57149 57879 57207 57885
rect 46698 57820 48360 57848
rect 48492 57851 48550 57857
rect 46698 57817 46710 57820
rect 46652 57811 46710 57817
rect 48492 57817 48504 57851
rect 48538 57848 48550 57851
rect 51074 57848 51080 57860
rect 48538 57820 51080 57848
rect 48538 57817 48550 57820
rect 48492 57811 48550 57817
rect 51074 57808 51080 57820
rect 51132 57808 51138 57860
rect 51804 57851 51862 57857
rect 51804 57817 51816 57851
rect 51850 57848 51862 57851
rect 52822 57848 52828 57860
rect 51850 57820 52828 57848
rect 51850 57817 51862 57820
rect 51804 57811 51862 57817
rect 52822 57808 52828 57820
rect 52880 57808 52886 57860
rect 55576 57851 55634 57857
rect 55576 57817 55588 57851
rect 55622 57848 55634 57851
rect 57416 57851 57474 57857
rect 55622 57820 57100 57848
rect 55622 57817 55634 57820
rect 55576 57811 55634 57817
rect 5994 57740 6000 57792
rect 6052 57780 6058 57792
rect 7009 57783 7067 57789
rect 7009 57780 7021 57783
rect 6052 57752 7021 57780
rect 6052 57740 6058 57752
rect 7009 57749 7021 57752
rect 7055 57749 7067 57783
rect 8938 57780 8944 57792
rect 8851 57752 8944 57780
rect 7009 57743 7067 57749
rect 8938 57740 8944 57752
rect 8996 57780 9002 57792
rect 10778 57780 10784 57792
rect 8996 57752 10784 57780
rect 8996 57740 9002 57752
rect 10778 57740 10784 57752
rect 10836 57740 10842 57792
rect 12158 57780 12164 57792
rect 12119 57752 12164 57780
rect 12158 57740 12164 57752
rect 12216 57740 12222 57792
rect 14090 57740 14096 57792
rect 14148 57780 14154 57792
rect 15749 57783 15807 57789
rect 15749 57780 15761 57783
rect 14148 57752 15761 57780
rect 14148 57740 14154 57752
rect 15749 57749 15761 57752
rect 15795 57749 15807 57783
rect 18690 57780 18696 57792
rect 18651 57752 18696 57780
rect 15749 57743 15807 57749
rect 18690 57740 18696 57752
rect 18748 57740 18754 57792
rect 27157 57783 27215 57789
rect 27157 57749 27169 57783
rect 27203 57780 27215 57783
rect 27246 57780 27252 57792
rect 27203 57752 27252 57780
rect 27203 57749 27215 57752
rect 27157 57743 27215 57749
rect 27246 57740 27252 57752
rect 27304 57740 27310 57792
rect 28994 57780 29000 57792
rect 28955 57752 29000 57780
rect 28994 57740 29000 57752
rect 29052 57740 29058 57792
rect 32306 57780 32312 57792
rect 32267 57752 32312 57780
rect 32306 57740 32312 57752
rect 32364 57740 32370 57792
rect 34146 57780 34152 57792
rect 34107 57752 34152 57780
rect 34146 57740 34152 57752
rect 34204 57740 34210 57792
rect 35434 57740 35440 57792
rect 35492 57780 35498 57792
rect 36725 57783 36783 57789
rect 36725 57780 36737 57783
rect 35492 57752 36737 57780
rect 35492 57740 35498 57752
rect 36725 57749 36737 57752
rect 36771 57749 36783 57783
rect 36725 57743 36783 57749
rect 41138 57740 41144 57792
rect 41196 57780 41202 57792
rect 41785 57783 41843 57789
rect 41785 57780 41797 57783
rect 41196 57752 41797 57780
rect 41196 57740 41202 57752
rect 41785 57749 41797 57752
rect 41831 57749 41843 57783
rect 41785 57743 41843 57749
rect 43162 57740 43168 57792
rect 43220 57780 43226 57792
rect 44453 57783 44511 57789
rect 44453 57780 44465 57783
rect 43220 57752 44465 57780
rect 43220 57740 43226 57752
rect 44453 57749 44465 57752
rect 44499 57749 44511 57783
rect 49602 57780 49608 57792
rect 49563 57752 49608 57780
rect 44453 57743 44511 57749
rect 49602 57740 49608 57752
rect 49660 57740 49666 57792
rect 56594 57740 56600 57792
rect 56652 57780 56658 57792
rect 56689 57783 56747 57789
rect 56689 57780 56701 57783
rect 56652 57752 56701 57780
rect 56652 57740 56658 57752
rect 56689 57749 56701 57752
rect 56735 57749 56747 57783
rect 57072 57780 57100 57820
rect 57416 57817 57428 57851
rect 57462 57848 57474 57851
rect 58434 57848 58440 57860
rect 57462 57820 58440 57848
rect 57462 57817 57474 57820
rect 57416 57811 57474 57817
rect 58434 57808 58440 57820
rect 58492 57808 58498 57860
rect 58529 57783 58587 57789
rect 58529 57780 58541 57783
rect 57072 57752 58541 57780
rect 56689 57743 56747 57749
rect 58529 57749 58541 57752
rect 58575 57749 58587 57783
rect 58529 57743 58587 57749
rect 1104 57690 59340 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 59340 57690
rect 1104 57616 59340 57638
rect 4982 57576 4988 57588
rect 4943 57548 4988 57576
rect 4982 57536 4988 57548
rect 5040 57536 5046 57588
rect 12802 57536 12808 57588
rect 12860 57576 12866 57588
rect 12897 57579 12955 57585
rect 12897 57576 12909 57579
rect 12860 57548 12909 57576
rect 12860 57536 12866 57548
rect 12897 57545 12909 57548
rect 12943 57545 12955 57579
rect 21266 57576 21272 57588
rect 21227 57548 21272 57576
rect 12897 57539 12955 57545
rect 21266 57536 21272 57548
rect 21324 57536 21330 57588
rect 26418 57576 26424 57588
rect 26379 57548 26424 57576
rect 26418 57536 26424 57548
rect 26476 57536 26482 57588
rect 31573 57579 31631 57585
rect 31573 57545 31585 57579
rect 31619 57576 31631 57579
rect 31846 57576 31852 57588
rect 31619 57548 31852 57576
rect 31619 57545 31631 57548
rect 31573 57539 31631 57545
rect 31846 57536 31852 57548
rect 31904 57536 31910 57588
rect 40313 57579 40371 57585
rect 40313 57545 40325 57579
rect 40359 57576 40371 57579
rect 40402 57576 40408 57588
rect 40359 57548 40408 57576
rect 40359 57545 40371 57548
rect 40313 57539 40371 57545
rect 40402 57536 40408 57548
rect 40460 57536 40466 57588
rect 49510 57536 49516 57588
rect 49568 57576 49574 57588
rect 50341 57579 50399 57585
rect 50341 57576 50353 57579
rect 49568 57548 50353 57576
rect 49568 57536 49574 57548
rect 50341 57545 50353 57548
rect 50387 57545 50399 57579
rect 50341 57539 50399 57545
rect 53374 57536 53380 57588
rect 53432 57576 53438 57588
rect 54389 57579 54447 57585
rect 54389 57576 54401 57579
rect 53432 57548 54401 57576
rect 53432 57536 53438 57548
rect 54389 57545 54401 57548
rect 54435 57545 54447 57579
rect 54389 57539 54447 57545
rect 11784 57511 11842 57517
rect 11784 57477 11796 57511
rect 11830 57508 11842 57511
rect 12158 57508 12164 57520
rect 11830 57480 12164 57508
rect 11830 57477 11842 57480
rect 11784 57471 11842 57477
rect 12158 57468 12164 57480
rect 12216 57468 12222 57520
rect 14360 57511 14418 57517
rect 14360 57477 14372 57511
rect 14406 57508 14418 57511
rect 15470 57508 15476 57520
rect 14406 57480 15476 57508
rect 14406 57477 14418 57480
rect 14360 57471 14418 57477
rect 15470 57468 15476 57480
rect 15528 57468 15534 57520
rect 18316 57511 18374 57517
rect 18316 57477 18328 57511
rect 18362 57508 18374 57511
rect 20622 57508 20628 57520
rect 18362 57480 20628 57508
rect 18362 57477 18374 57480
rect 18316 57471 18374 57477
rect 20622 57468 20628 57480
rect 20680 57468 20686 57520
rect 23468 57511 23526 57517
rect 23468 57477 23480 57511
rect 23514 57508 23526 57511
rect 24118 57508 24124 57520
rect 23514 57480 24124 57508
rect 23514 57477 23526 57480
rect 23468 57471 23526 57477
rect 24118 57468 24124 57480
rect 24176 57468 24182 57520
rect 25308 57511 25366 57517
rect 25308 57477 25320 57511
rect 25354 57508 25366 57511
rect 27154 57508 27160 57520
rect 25354 57480 27160 57508
rect 25354 57477 25366 57480
rect 25308 57471 25366 57477
rect 27154 57468 27160 57480
rect 27212 57468 27218 57520
rect 27884 57511 27942 57517
rect 27884 57477 27896 57511
rect 27930 57508 27942 57511
rect 28994 57508 29000 57520
rect 27930 57480 29000 57508
rect 27930 57477 27942 57480
rect 27884 57471 27942 57477
rect 28994 57468 29000 57480
rect 29052 57468 29058 57520
rect 30460 57511 30518 57517
rect 30460 57477 30472 57511
rect 30506 57508 30518 57511
rect 32306 57508 32312 57520
rect 30506 57480 32312 57508
rect 30506 57477 30518 57480
rect 30460 57471 30518 57477
rect 32306 57468 32312 57480
rect 32364 57468 32370 57520
rect 34146 57468 34152 57520
rect 34204 57508 34210 57520
rect 34946 57511 35004 57517
rect 34946 57508 34958 57511
rect 34204 57480 34958 57508
rect 34204 57468 34210 57480
rect 34946 57477 34958 57480
rect 34992 57477 35004 57511
rect 39022 57508 39028 57520
rect 38983 57480 39028 57508
rect 34946 57471 35004 57477
rect 39022 57468 39028 57480
rect 39080 57508 39086 57520
rect 41782 57508 41788 57520
rect 39080 57480 41788 57508
rect 39080 57468 39086 57480
rect 41782 57468 41788 57480
rect 41840 57468 41846 57520
rect 42794 57508 42800 57520
rect 42444 57480 42800 57508
rect 3872 57443 3930 57449
rect 3872 57409 3884 57443
rect 3918 57440 3930 57443
rect 5166 57440 5172 57452
rect 3918 57412 5172 57440
rect 3918 57409 3930 57412
rect 3872 57403 3930 57409
rect 5166 57400 5172 57412
rect 5224 57400 5230 57452
rect 7184 57443 7242 57449
rect 7184 57409 7196 57443
rect 7230 57440 7242 57443
rect 8294 57440 8300 57452
rect 7230 57412 8300 57440
rect 7230 57409 7242 57412
rect 7184 57403 7242 57409
rect 8294 57400 8300 57412
rect 8352 57400 8358 57452
rect 8754 57440 8760 57452
rect 8667 57412 8760 57440
rect 8754 57400 8760 57412
rect 8812 57440 8818 57452
rect 13814 57440 13820 57452
rect 8812 57412 13820 57440
rect 8812 57400 8818 57412
rect 13814 57400 13820 57412
rect 13872 57400 13878 57452
rect 14090 57440 14096 57452
rect 14051 57412 14096 57440
rect 14090 57400 14096 57412
rect 14148 57400 14154 57452
rect 18046 57440 18052 57452
rect 18007 57412 18052 57440
rect 18046 57400 18052 57412
rect 18104 57440 18110 57452
rect 19886 57440 19892 57452
rect 18104 57412 19892 57440
rect 18104 57400 18110 57412
rect 19886 57400 19892 57412
rect 19944 57400 19950 57452
rect 20156 57443 20214 57449
rect 20156 57409 20168 57443
rect 20202 57440 20214 57443
rect 23750 57440 23756 57452
rect 20202 57412 23756 57440
rect 20202 57409 20214 57412
rect 20156 57403 20214 57409
rect 23750 57400 23756 57412
rect 23808 57400 23814 57452
rect 30193 57443 30251 57449
rect 30193 57409 30205 57443
rect 30239 57440 30251 57443
rect 30282 57440 30288 57452
rect 30239 57412 30288 57440
rect 30239 57409 30251 57412
rect 30193 57403 30251 57409
rect 30282 57400 30288 57412
rect 30340 57400 30346 57452
rect 33128 57443 33186 57449
rect 33128 57409 33140 57443
rect 33174 57440 33186 57443
rect 34054 57440 34060 57452
rect 33174 57412 34060 57440
rect 33174 57409 33186 57412
rect 33128 57403 33186 57409
rect 34054 57400 34060 57412
rect 34112 57400 34118 57452
rect 42444 57449 42472 57480
rect 42794 57468 42800 57480
rect 42852 57468 42858 57520
rect 51068 57511 51126 57517
rect 51068 57477 51080 57511
rect 51114 57508 51126 57511
rect 52178 57508 52184 57520
rect 51114 57480 52184 57508
rect 51114 57477 51126 57480
rect 51068 57471 51126 57477
rect 52178 57468 52184 57480
rect 52236 57468 52242 57520
rect 53098 57508 53104 57520
rect 53059 57480 53104 57508
rect 53098 57468 53104 57480
rect 53156 57508 53162 57520
rect 56134 57508 56140 57520
rect 53156 57480 56140 57508
rect 53156 57468 53162 57480
rect 56134 57468 56140 57480
rect 56192 57468 56198 57520
rect 42429 57443 42487 57449
rect 42429 57409 42441 57443
rect 42475 57409 42487 57443
rect 42429 57403 42487 57409
rect 42696 57443 42754 57449
rect 42696 57409 42708 57443
rect 42742 57440 42754 57443
rect 43806 57440 43812 57452
rect 42742 57412 43812 57440
rect 42742 57409 42754 57412
rect 42696 57403 42754 57409
rect 43806 57400 43812 57412
rect 43864 57400 43870 57452
rect 44266 57440 44272 57452
rect 44227 57412 44272 57440
rect 44266 57400 44272 57412
rect 44324 57400 44330 57452
rect 44536 57443 44594 57449
rect 44536 57409 44548 57443
rect 44582 57440 44594 57443
rect 45646 57440 45652 57452
rect 44582 57412 45652 57440
rect 44582 57409 44594 57412
rect 44536 57403 44594 57409
rect 45646 57400 45652 57412
rect 45704 57400 45710 57452
rect 49228 57443 49286 57449
rect 49228 57409 49240 57443
rect 49274 57440 49286 57443
rect 51534 57440 51540 57452
rect 49274 57412 51540 57440
rect 49274 57409 49286 57412
rect 49228 57403 49286 57409
rect 51534 57400 51540 57412
rect 51592 57400 51598 57452
rect 55214 57400 55220 57452
rect 55272 57440 55278 57452
rect 55309 57443 55367 57449
rect 55309 57440 55321 57443
rect 55272 57412 55321 57440
rect 55272 57400 55278 57412
rect 55309 57409 55321 57412
rect 55355 57409 55367 57443
rect 55309 57403 55367 57409
rect 55576 57443 55634 57449
rect 55576 57409 55588 57443
rect 55622 57440 55634 57443
rect 56686 57440 56692 57452
rect 55622 57412 56692 57440
rect 55622 57409 55634 57412
rect 55576 57403 55634 57409
rect 56686 57400 56692 57412
rect 56744 57400 56750 57452
rect 3605 57375 3663 57381
rect 3605 57341 3617 57375
rect 3651 57341 3663 57375
rect 3605 57335 3663 57341
rect 3620 57236 3648 57335
rect 6914 57332 6920 57384
rect 6972 57372 6978 57384
rect 10505 57375 10563 57381
rect 6972 57344 7017 57372
rect 6972 57332 6978 57344
rect 10505 57341 10517 57375
rect 10551 57372 10563 57375
rect 10778 57372 10784 57384
rect 10551 57344 10784 57372
rect 10551 57341 10563 57344
rect 10505 57335 10563 57341
rect 10778 57332 10784 57344
rect 10836 57372 10842 57384
rect 11517 57375 11575 57381
rect 11517 57372 11529 57375
rect 10836 57344 11529 57372
rect 10836 57332 10842 57344
rect 11517 57341 11529 57344
rect 11563 57341 11575 57375
rect 11517 57335 11575 57341
rect 22462 57332 22468 57384
rect 22520 57372 22526 57384
rect 23201 57375 23259 57381
rect 23201 57372 23213 57375
rect 22520 57344 23213 57372
rect 22520 57332 22526 57344
rect 23201 57341 23213 57344
rect 23247 57341 23259 57375
rect 25038 57372 25044 57384
rect 23201 57335 23259 57341
rect 24228 57344 25044 57372
rect 3878 57236 3884 57248
rect 3620 57208 3884 57236
rect 3878 57196 3884 57208
rect 3936 57196 3942 57248
rect 8297 57239 8355 57245
rect 8297 57205 8309 57239
rect 8343 57236 8355 57239
rect 8386 57236 8392 57248
rect 8343 57208 8392 57236
rect 8343 57205 8355 57208
rect 8297 57199 8355 57205
rect 8386 57196 8392 57208
rect 8444 57196 8450 57248
rect 15470 57236 15476 57248
rect 15431 57208 15476 57236
rect 15470 57196 15476 57208
rect 15528 57196 15534 57248
rect 19426 57236 19432 57248
rect 19387 57208 19432 57236
rect 19426 57196 19432 57208
rect 19484 57196 19490 57248
rect 23216 57236 23244 57335
rect 24228 57236 24256 57344
rect 25038 57332 25044 57344
rect 25096 57332 25102 57384
rect 27522 57332 27528 57384
rect 27580 57372 27586 57384
rect 27617 57375 27675 57381
rect 27617 57372 27629 57375
rect 27580 57344 27629 57372
rect 27580 57332 27586 57344
rect 27617 57341 27629 57344
rect 27663 57341 27675 57375
rect 27617 57335 27675 57341
rect 32766 57332 32772 57384
rect 32824 57372 32830 57384
rect 32861 57375 32919 57381
rect 32861 57372 32873 57375
rect 32824 57344 32873 57372
rect 32824 57332 32830 57344
rect 32861 57341 32873 57344
rect 32907 57341 32919 57375
rect 34698 57372 34704 57384
rect 34659 57344 34704 57372
rect 32861 57335 32919 57341
rect 34698 57332 34704 57344
rect 34756 57332 34762 57384
rect 48958 57372 48964 57384
rect 48919 57344 48964 57372
rect 48958 57332 48964 57344
rect 49016 57332 49022 57384
rect 50154 57332 50160 57384
rect 50212 57372 50218 57384
rect 50798 57372 50804 57384
rect 50212 57344 50804 57372
rect 50212 57332 50218 57344
rect 50798 57332 50804 57344
rect 50856 57332 50862 57384
rect 24578 57236 24584 57248
rect 23216 57208 24256 57236
rect 24539 57208 24584 57236
rect 24578 57196 24584 57208
rect 24636 57196 24642 57248
rect 28994 57236 29000 57248
rect 28955 57208 29000 57236
rect 28994 57196 29000 57208
rect 29052 57196 29058 57248
rect 31202 57196 31208 57248
rect 31260 57236 31266 57248
rect 34241 57239 34299 57245
rect 34241 57236 34253 57239
rect 31260 57208 34253 57236
rect 31260 57196 31266 57208
rect 34241 57205 34253 57208
rect 34287 57205 34299 57239
rect 36078 57236 36084 57248
rect 36039 57208 36084 57236
rect 34241 57199 34299 57205
rect 36078 57196 36084 57208
rect 36136 57196 36142 57248
rect 43809 57239 43867 57245
rect 43809 57205 43821 57239
rect 43855 57236 43867 57239
rect 44542 57236 44548 57248
rect 43855 57208 44548 57236
rect 43855 57205 43867 57208
rect 43809 57199 43867 57205
rect 44542 57196 44548 57208
rect 44600 57196 44606 57248
rect 45554 57196 45560 57248
rect 45612 57236 45618 57248
rect 45649 57239 45707 57245
rect 45649 57236 45661 57239
rect 45612 57208 45661 57236
rect 45612 57196 45618 57208
rect 45649 57205 45661 57208
rect 45695 57205 45707 57239
rect 52178 57236 52184 57248
rect 52139 57208 52184 57236
rect 45649 57199 45707 57205
rect 52178 57196 52184 57208
rect 52236 57196 52242 57248
rect 56689 57239 56747 57245
rect 56689 57205 56701 57239
rect 56735 57236 56747 57239
rect 57238 57236 57244 57248
rect 56735 57208 57244 57236
rect 56735 57205 56747 57208
rect 56689 57199 56747 57205
rect 57238 57196 57244 57208
rect 57296 57196 57302 57248
rect 1104 57146 59340 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 59340 57146
rect 1104 57072 59340 57094
rect 5166 57032 5172 57044
rect 5127 57004 5172 57032
rect 5166 56992 5172 57004
rect 5224 56992 5230 57044
rect 8294 57032 8300 57044
rect 8255 57004 8300 57032
rect 8294 56992 8300 57004
rect 8352 56992 8358 57044
rect 12250 56992 12256 57044
rect 12308 57032 12314 57044
rect 12897 57035 12955 57041
rect 12897 57032 12909 57035
rect 12308 57004 12909 57032
rect 12308 56992 12314 57004
rect 12897 57001 12909 57004
rect 12943 57001 12955 57035
rect 15838 57032 15844 57044
rect 15799 57004 15844 57032
rect 12897 56995 12955 57001
rect 15838 56992 15844 57004
rect 15896 56992 15902 57044
rect 18598 56992 18604 57044
rect 18656 57032 18662 57044
rect 18693 57035 18751 57041
rect 18693 57032 18705 57035
rect 18656 57004 18705 57032
rect 18656 56992 18662 57004
rect 18693 57001 18705 57004
rect 18739 57001 18751 57035
rect 23842 57032 23848 57044
rect 23803 57004 23848 57032
rect 18693 56995 18751 57001
rect 23842 56992 23848 57004
rect 23900 56992 23906 57044
rect 25038 56992 25044 57044
rect 25096 57032 25102 57044
rect 26053 57035 26111 57041
rect 26053 57032 26065 57035
rect 25096 57004 26065 57032
rect 25096 56992 25102 57004
rect 26053 57001 26065 57004
rect 26099 57001 26111 57035
rect 28902 57032 28908 57044
rect 28863 57004 28908 57032
rect 26053 56995 26111 57001
rect 28902 56992 28908 57004
rect 28960 56992 28966 57044
rect 32214 56992 32220 57044
rect 32272 57032 32278 57044
rect 32309 57035 32367 57041
rect 32309 57032 32321 57035
rect 32272 57004 32321 57032
rect 32272 56992 32278 57004
rect 32309 57001 32321 57004
rect 32355 57001 32367 57035
rect 32309 56995 32367 57001
rect 34054 56992 34060 57044
rect 34112 57032 34118 57044
rect 34149 57035 34207 57041
rect 34149 57032 34161 57035
rect 34112 57004 34161 57032
rect 34112 56992 34118 57004
rect 34149 57001 34161 57004
rect 34195 57001 34207 57035
rect 38654 57032 38660 57044
rect 38615 57004 38660 57032
rect 34149 56995 34207 57001
rect 38654 56992 38660 57004
rect 38712 56992 38718 57044
rect 49418 56992 49424 57044
rect 49476 57032 49482 57044
rect 49605 57035 49663 57041
rect 49605 57032 49617 57035
rect 49476 57004 49617 57032
rect 49476 56992 49482 57004
rect 49605 57001 49617 57004
rect 49651 57001 49663 57035
rect 49605 56995 49663 57001
rect 52822 56992 52828 57044
rect 52880 57032 52886 57044
rect 52917 57035 52975 57041
rect 52917 57032 52929 57035
rect 52880 57004 52929 57032
rect 52880 56992 52886 57004
rect 52917 57001 52929 57004
rect 52963 57001 52975 57035
rect 52917 56995 52975 57001
rect 54757 57035 54815 57041
rect 54757 57001 54769 57035
rect 54803 57032 54815 57035
rect 54846 57032 54852 57044
rect 54803 57004 54852 57032
rect 54803 57001 54815 57004
rect 54757 56995 54815 57001
rect 54846 56992 54852 57004
rect 54904 56992 54910 57044
rect 56686 57032 56692 57044
rect 56647 57004 56692 57032
rect 56686 56992 56692 57004
rect 56744 56992 56750 57044
rect 58434 56992 58440 57044
rect 58492 57032 58498 57044
rect 58529 57035 58587 57041
rect 58529 57032 58541 57035
rect 58492 57004 58541 57032
rect 58492 56992 58498 57004
rect 58529 57001 58541 57004
rect 58575 57001 58587 57035
rect 58529 56995 58587 57001
rect 8938 56896 8944 56908
rect 8899 56868 8944 56896
rect 8938 56856 8944 56868
rect 8996 56856 9002 56908
rect 14090 56856 14096 56908
rect 14148 56896 14154 56908
rect 14461 56899 14519 56905
rect 14461 56896 14473 56899
rect 14148 56868 14473 56896
rect 14148 56856 14154 56868
rect 14461 56865 14473 56868
rect 14507 56865 14519 56899
rect 19886 56896 19892 56908
rect 19847 56868 19892 56896
rect 14461 56859 14519 56865
rect 19886 56856 19892 56868
rect 19944 56856 19950 56908
rect 22462 56896 22468 56908
rect 22423 56868 22468 56896
rect 22462 56856 22468 56868
rect 22520 56856 22526 56908
rect 32766 56896 32772 56908
rect 32727 56868 32772 56896
rect 32766 56856 32772 56868
rect 32824 56856 32830 56908
rect 37274 56896 37280 56908
rect 37235 56868 37280 56896
rect 37274 56856 37280 56868
rect 37332 56856 37338 56908
rect 40402 56856 40408 56908
rect 40460 56896 40466 56908
rect 40865 56899 40923 56905
rect 40865 56896 40877 56899
rect 40460 56868 40877 56896
rect 40460 56856 40466 56868
rect 40865 56865 40877 56868
rect 40911 56865 40923 56899
rect 42702 56896 42708 56908
rect 42663 56868 42708 56896
rect 40865 56859 40923 56865
rect 42702 56856 42708 56868
rect 42760 56856 42766 56908
rect 44266 56856 44272 56908
rect 44324 56896 44330 56908
rect 45002 56896 45008 56908
rect 44324 56868 45008 56896
rect 44324 56856 44330 56868
rect 45002 56856 45008 56868
rect 45060 56856 45066 56908
rect 50154 56856 50160 56908
rect 50212 56896 50218 56908
rect 51537 56899 51595 56905
rect 51537 56896 51549 56899
rect 50212 56868 51549 56896
rect 50212 56856 50218 56868
rect 51537 56865 51549 56868
rect 51583 56865 51595 56899
rect 51537 56859 51595 56865
rect 3789 56831 3847 56837
rect 3789 56797 3801 56831
rect 3835 56828 3847 56831
rect 3878 56828 3884 56840
rect 3835 56800 3884 56828
rect 3835 56797 3847 56800
rect 3789 56791 3847 56797
rect 3878 56788 3884 56800
rect 3936 56788 3942 56840
rect 6914 56788 6920 56840
rect 6972 56828 6978 56840
rect 7184 56831 7242 56837
rect 6972 56800 7017 56828
rect 6972 56788 6978 56800
rect 7184 56797 7196 56831
rect 7230 56828 7242 56831
rect 8294 56828 8300 56840
rect 7230 56800 8300 56828
rect 7230 56797 7242 56800
rect 7184 56791 7242 56797
rect 8294 56788 8300 56800
rect 8352 56788 8358 56840
rect 11514 56828 11520 56840
rect 11475 56800 11520 56828
rect 11514 56788 11520 56800
rect 11572 56788 11578 56840
rect 11784 56831 11842 56837
rect 11784 56797 11796 56831
rect 11830 56828 11842 56831
rect 12894 56828 12900 56840
rect 11830 56800 12900 56828
rect 11830 56797 11842 56800
rect 11784 56791 11842 56797
rect 12894 56788 12900 56800
rect 12952 56788 12958 56840
rect 14728 56831 14786 56837
rect 14728 56797 14740 56831
rect 14774 56828 14786 56831
rect 15470 56828 15476 56840
rect 14774 56800 15476 56828
rect 14774 56797 14786 56800
rect 14728 56791 14786 56797
rect 15470 56788 15476 56800
rect 15528 56788 15534 56840
rect 17313 56831 17371 56837
rect 17313 56797 17325 56831
rect 17359 56828 17371 56831
rect 17862 56828 17868 56840
rect 17359 56800 17868 56828
rect 17359 56797 17371 56800
rect 17313 56791 17371 56797
rect 17862 56788 17868 56800
rect 17920 56788 17926 56840
rect 20162 56837 20168 56840
rect 20156 56828 20168 56837
rect 20123 56800 20168 56828
rect 20156 56791 20168 56800
rect 20162 56788 20168 56791
rect 20220 56788 20226 56840
rect 22732 56831 22790 56837
rect 22732 56797 22744 56831
rect 22778 56828 22790 56831
rect 24578 56828 24584 56840
rect 22778 56800 24584 56828
rect 22778 56797 22790 56800
rect 22732 56791 22790 56797
rect 24578 56788 24584 56800
rect 24636 56788 24642 56840
rect 26970 56788 26976 56840
rect 27028 56828 27034 56840
rect 27522 56828 27528 56840
rect 27028 56800 27528 56828
rect 27028 56788 27034 56800
rect 27522 56788 27528 56800
rect 27580 56788 27586 56840
rect 27792 56831 27850 56837
rect 27792 56797 27804 56831
rect 27838 56828 27850 56831
rect 28994 56828 29000 56840
rect 27838 56800 29000 56828
rect 27838 56797 27850 56800
rect 27792 56791 27850 56797
rect 28994 56788 29000 56800
rect 29052 56788 29058 56840
rect 31202 56837 31208 56840
rect 30929 56831 30987 56837
rect 30929 56797 30941 56831
rect 30975 56797 30987 56831
rect 31196 56828 31208 56837
rect 31163 56800 31208 56828
rect 30929 56791 30987 56797
rect 31196 56791 31208 56800
rect 4056 56763 4114 56769
rect 4056 56729 4068 56763
rect 4102 56760 4114 56763
rect 4982 56760 4988 56772
rect 4102 56732 4988 56760
rect 4102 56729 4114 56732
rect 4056 56723 4114 56729
rect 4982 56720 4988 56732
rect 5040 56720 5046 56772
rect 9208 56763 9266 56769
rect 9208 56729 9220 56763
rect 9254 56760 9266 56763
rect 17580 56763 17638 56769
rect 9254 56732 12434 56760
rect 9254 56729 9266 56732
rect 9208 56723 9266 56729
rect 10318 56692 10324 56704
rect 10279 56664 10324 56692
rect 10318 56652 10324 56664
rect 10376 56652 10382 56704
rect 12406 56692 12434 56732
rect 17580 56729 17592 56763
rect 17626 56760 17638 56763
rect 19242 56760 19248 56772
rect 17626 56732 19248 56760
rect 17626 56729 17638 56732
rect 17580 56723 17638 56729
rect 19242 56720 19248 56732
rect 19300 56720 19306 56772
rect 24765 56763 24823 56769
rect 24765 56729 24777 56763
rect 24811 56760 24823 56763
rect 27614 56760 27620 56772
rect 24811 56732 27620 56760
rect 24811 56729 24823 56732
rect 24765 56723 24823 56729
rect 27614 56720 27620 56732
rect 27672 56720 27678 56772
rect 30944 56760 30972 56791
rect 31202 56788 31208 56791
rect 31260 56788 31266 56840
rect 32858 56788 32864 56840
rect 32916 56828 32922 56840
rect 34698 56828 34704 56840
rect 32916 56800 34704 56828
rect 32916 56788 32922 56800
rect 34698 56788 34704 56800
rect 34756 56788 34762 56840
rect 34968 56831 35026 56837
rect 34968 56797 34980 56831
rect 35014 56828 35026 56831
rect 36078 56828 36084 56840
rect 35014 56800 36084 56828
rect 35014 56797 35026 56800
rect 34968 56791 35026 56797
rect 36078 56788 36084 56800
rect 36136 56788 36142 56840
rect 41138 56837 41144 56840
rect 41132 56828 41144 56837
rect 41099 56800 41144 56828
rect 41132 56791 41144 56800
rect 41138 56788 41144 56791
rect 41196 56788 41202 56840
rect 48498 56837 48504 56840
rect 48225 56831 48283 56837
rect 48225 56797 48237 56831
rect 48271 56797 48283 56831
rect 48492 56828 48504 56837
rect 48459 56800 48504 56828
rect 48225 56791 48283 56797
rect 48492 56791 48504 56800
rect 32766 56760 32772 56772
rect 30944 56732 32772 56760
rect 32766 56720 32772 56732
rect 32824 56720 32830 56772
rect 33036 56763 33094 56769
rect 33036 56729 33048 56763
rect 33082 56760 33094 56763
rect 34238 56760 34244 56772
rect 33082 56732 34244 56760
rect 33082 56729 33094 56732
rect 33036 56723 33094 56729
rect 34238 56720 34244 56732
rect 34296 56720 34302 56772
rect 37544 56763 37602 56769
rect 37544 56729 37556 56763
rect 37590 56760 37602 56763
rect 39022 56760 39028 56772
rect 37590 56732 39028 56760
rect 37590 56729 37602 56732
rect 37544 56723 37602 56729
rect 39022 56720 39028 56732
rect 39080 56720 39086 56772
rect 42794 56720 42800 56772
rect 42852 56760 42858 56772
rect 42950 56763 43008 56769
rect 42950 56760 42962 56763
rect 42852 56732 42962 56760
rect 42852 56720 42858 56732
rect 42950 56729 42962 56732
rect 42996 56729 43008 56763
rect 42950 56723 43008 56729
rect 45272 56763 45330 56769
rect 45272 56729 45284 56763
rect 45318 56760 45330 56763
rect 46290 56760 46296 56772
rect 45318 56732 46296 56760
rect 45318 56729 45330 56732
rect 45272 56723 45330 56729
rect 46290 56720 46296 56732
rect 46348 56720 46354 56772
rect 48240 56760 48268 56791
rect 48498 56788 48504 56791
rect 48556 56788 48562 56840
rect 48958 56760 48964 56772
rect 48240 56732 48964 56760
rect 48958 56720 48964 56732
rect 49016 56720 49022 56772
rect 51552 56760 51580 56859
rect 55214 56856 55220 56908
rect 55272 56896 55278 56908
rect 55309 56899 55367 56905
rect 55309 56896 55321 56899
rect 55272 56868 55321 56896
rect 55272 56856 55278 56868
rect 55309 56865 55321 56868
rect 55355 56865 55367 56899
rect 55309 56859 55367 56865
rect 51804 56831 51862 56837
rect 51804 56797 51816 56831
rect 51850 56828 51862 56831
rect 52546 56828 52552 56840
rect 51850 56800 52552 56828
rect 51850 56797 51862 56800
rect 51804 56791 51862 56797
rect 52546 56788 52552 56800
rect 52604 56788 52610 56840
rect 53374 56828 53380 56840
rect 52656 56800 53380 56828
rect 52656 56772 52684 56800
rect 53374 56788 53380 56800
rect 53432 56788 53438 56840
rect 56870 56828 56876 56840
rect 55508 56800 56876 56828
rect 52638 56760 52644 56772
rect 51552 56732 52644 56760
rect 52638 56720 52644 56732
rect 52696 56720 52702 56772
rect 53644 56763 53702 56769
rect 53644 56729 53656 56763
rect 53690 56760 53702 56763
rect 55508 56760 55536 56800
rect 56870 56788 56876 56800
rect 56928 56788 56934 56840
rect 57054 56788 57060 56840
rect 57112 56828 57118 56840
rect 57149 56831 57207 56837
rect 57149 56828 57161 56831
rect 57112 56800 57161 56828
rect 57112 56788 57118 56800
rect 57149 56797 57161 56800
rect 57195 56797 57207 56831
rect 57149 56791 57207 56797
rect 57238 56788 57244 56840
rect 57296 56828 57302 56840
rect 57405 56831 57463 56837
rect 57405 56828 57417 56831
rect 57296 56800 57417 56828
rect 57296 56788 57302 56800
rect 57405 56797 57417 56800
rect 57451 56797 57463 56831
rect 57405 56791 57463 56797
rect 53690 56732 55536 56760
rect 55576 56763 55634 56769
rect 53690 56729 53702 56732
rect 53644 56723 53702 56729
rect 55576 56729 55588 56763
rect 55622 56760 55634 56763
rect 55674 56760 55680 56772
rect 55622 56732 55680 56760
rect 55622 56729 55634 56732
rect 55576 56723 55634 56729
rect 55674 56720 55680 56732
rect 55732 56720 55738 56772
rect 20990 56692 20996 56704
rect 12406 56664 20996 56692
rect 20990 56652 20996 56664
rect 21048 56652 21054 56704
rect 21266 56692 21272 56704
rect 21227 56664 21272 56692
rect 21266 56652 21272 56664
rect 21324 56652 21330 56704
rect 36078 56692 36084 56704
rect 36039 56664 36084 56692
rect 36078 56652 36084 56664
rect 36136 56652 36142 56704
rect 42242 56692 42248 56704
rect 42203 56664 42248 56692
rect 42242 56652 42248 56664
rect 42300 56652 42306 56704
rect 42334 56652 42340 56704
rect 42392 56692 42398 56704
rect 44085 56695 44143 56701
rect 44085 56692 44097 56695
rect 42392 56664 44097 56692
rect 42392 56652 42398 56664
rect 44085 56661 44097 56664
rect 44131 56661 44143 56695
rect 46382 56692 46388 56704
rect 46343 56664 46388 56692
rect 44085 56655 44143 56661
rect 46382 56652 46388 56664
rect 46440 56652 46446 56704
rect 1104 56602 59340 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 59340 56602
rect 1104 56528 59340 56550
rect 4982 56488 4988 56500
rect 4943 56460 4988 56488
rect 4982 56448 4988 56460
rect 5040 56448 5046 56500
rect 8294 56488 8300 56500
rect 8255 56460 8300 56488
rect 8294 56448 8300 56460
rect 8352 56448 8358 56500
rect 8938 56448 8944 56500
rect 8996 56448 9002 56500
rect 14645 56491 14703 56497
rect 14645 56457 14657 56491
rect 14691 56488 14703 56491
rect 15930 56488 15936 56500
rect 14691 56460 15936 56488
rect 14691 56457 14703 56460
rect 14645 56451 14703 56457
rect 15930 56448 15936 56460
rect 15988 56448 15994 56500
rect 23750 56488 23756 56500
rect 23711 56460 23756 56488
rect 23750 56448 23756 56460
rect 23808 56448 23814 56500
rect 34238 56488 34244 56500
rect 34199 56460 34244 56488
rect 34238 56448 34244 56460
rect 34296 56448 34302 56500
rect 39022 56488 39028 56500
rect 38983 56460 39028 56488
rect 39022 56448 39028 56460
rect 39080 56448 39086 56500
rect 41785 56491 41843 56497
rect 41785 56457 41797 56491
rect 41831 56488 41843 56491
rect 42794 56488 42800 56500
rect 41831 56460 42800 56488
rect 41831 56457 41843 56460
rect 41785 56451 41843 56457
rect 42794 56448 42800 56460
rect 42852 56448 42858 56500
rect 43806 56488 43812 56500
rect 43767 56460 43812 56488
rect 43806 56448 43812 56460
rect 43864 56448 43870 56500
rect 45646 56488 45652 56500
rect 45607 56460 45652 56488
rect 45646 56448 45652 56460
rect 45704 56448 45710 56500
rect 50341 56491 50399 56497
rect 50341 56457 50353 56491
rect 50387 56488 50399 56491
rect 50614 56488 50620 56500
rect 50387 56460 50620 56488
rect 50387 56457 50399 56460
rect 50341 56451 50399 56457
rect 50614 56448 50620 56460
rect 50672 56448 50678 56500
rect 55674 56488 55680 56500
rect 55635 56460 55680 56488
rect 55674 56448 55680 56460
rect 55732 56448 55738 56500
rect 3872 56355 3930 56361
rect 3872 56321 3884 56355
rect 3918 56352 3930 56355
rect 5166 56352 5172 56364
rect 3918 56324 5172 56352
rect 3918 56321 3930 56324
rect 3872 56315 3930 56321
rect 5166 56312 5172 56324
rect 5224 56312 5230 56364
rect 7184 56355 7242 56361
rect 7184 56321 7196 56355
rect 7230 56352 7242 56355
rect 8202 56352 8208 56364
rect 7230 56324 8208 56352
rect 7230 56321 7242 56324
rect 7184 56315 7242 56321
rect 8202 56312 8208 56324
rect 8260 56312 8266 56364
rect 8757 56355 8815 56361
rect 8757 56321 8769 56355
rect 8803 56352 8815 56355
rect 8956 56352 8984 56448
rect 9024 56423 9082 56429
rect 9024 56389 9036 56423
rect 9070 56420 9082 56423
rect 10318 56420 10324 56432
rect 9070 56392 10324 56420
rect 9070 56389 9082 56392
rect 9024 56383 9082 56389
rect 10318 56380 10324 56392
rect 10376 56380 10382 56432
rect 11514 56380 11520 56432
rect 11572 56420 11578 56432
rect 14090 56420 14096 56432
rect 11572 56392 14096 56420
rect 11572 56380 11578 56392
rect 12820 56361 12848 56392
rect 14090 56380 14096 56392
rect 14148 56380 14154 56432
rect 15004 56423 15062 56429
rect 15004 56389 15016 56423
rect 15050 56420 15062 56423
rect 17310 56420 17316 56432
rect 15050 56392 17316 56420
rect 15050 56389 15062 56392
rect 15004 56383 15062 56389
rect 17310 56380 17316 56392
rect 17368 56380 17374 56432
rect 18316 56423 18374 56429
rect 18316 56389 18328 56423
rect 18362 56420 18374 56423
rect 19426 56420 19432 56432
rect 18362 56392 19432 56420
rect 18362 56389 18374 56392
rect 18316 56383 18374 56389
rect 19426 56380 19432 56392
rect 19484 56380 19490 56432
rect 20156 56423 20214 56429
rect 20156 56389 20168 56423
rect 20202 56420 20214 56423
rect 21266 56420 21272 56432
rect 20202 56392 21272 56420
rect 20202 56389 20214 56392
rect 20156 56383 20214 56389
rect 21266 56380 21272 56392
rect 21324 56380 21330 56432
rect 22640 56423 22698 56429
rect 22640 56389 22652 56423
rect 22686 56420 22698 56423
rect 23474 56420 23480 56432
rect 22686 56392 23480 56420
rect 22686 56389 22698 56392
rect 22640 56383 22698 56389
rect 23474 56380 23480 56392
rect 23532 56380 23538 56432
rect 27614 56380 27620 56432
rect 27672 56420 27678 56432
rect 27985 56423 28043 56429
rect 27985 56420 27997 56423
rect 27672 56392 27997 56420
rect 27672 56380 27678 56392
rect 27985 56389 27997 56392
rect 28031 56389 28043 56423
rect 27985 56383 28043 56389
rect 34968 56423 35026 56429
rect 34968 56389 34980 56423
rect 35014 56420 35026 56423
rect 36078 56420 36084 56432
rect 35014 56392 36084 56420
rect 35014 56389 35026 56392
rect 34968 56383 35026 56389
rect 36078 56380 36084 56392
rect 36136 56380 36142 56432
rect 40672 56423 40730 56429
rect 40672 56389 40684 56423
rect 40718 56420 40730 56423
rect 42242 56420 42248 56432
rect 40718 56392 42248 56420
rect 40718 56389 40730 56392
rect 40672 56383 40730 56389
rect 42242 56380 42248 56392
rect 42300 56380 42306 56432
rect 44542 56429 44548 56432
rect 44536 56420 44548 56429
rect 44503 56392 44548 56420
rect 44536 56383 44548 56392
rect 44542 56380 44548 56383
rect 44600 56380 44606 56432
rect 49228 56423 49286 56429
rect 49228 56389 49240 56423
rect 49274 56420 49286 56423
rect 49602 56420 49608 56432
rect 49274 56392 49608 56420
rect 49274 56389 49286 56392
rect 49228 56383 49286 56389
rect 49602 56380 49608 56392
rect 49660 56380 49666 56432
rect 51068 56423 51126 56429
rect 51068 56389 51080 56423
rect 51114 56420 51126 56423
rect 52178 56420 52184 56432
rect 51114 56392 52184 56420
rect 51114 56389 51126 56392
rect 51068 56383 51126 56389
rect 52178 56380 52184 56392
rect 52236 56380 52242 56432
rect 55122 56420 55128 56432
rect 54312 56392 55128 56420
rect 8803 56324 8984 56352
rect 12805 56355 12863 56361
rect 8803 56321 8815 56324
rect 8757 56315 8815 56321
rect 12805 56321 12817 56355
rect 12851 56321 12863 56355
rect 12805 56315 12863 56321
rect 13072 56355 13130 56361
rect 13072 56321 13084 56355
rect 13118 56352 13130 56355
rect 15562 56352 15568 56364
rect 13118 56324 15568 56352
rect 13118 56321 13130 56324
rect 13072 56315 13130 56321
rect 15562 56312 15568 56324
rect 15620 56312 15626 56364
rect 19889 56355 19947 56361
rect 19889 56321 19901 56355
rect 19935 56352 19947 56355
rect 19978 56352 19984 56364
rect 19935 56324 19984 56352
rect 19935 56321 19947 56324
rect 19889 56315 19947 56321
rect 19978 56312 19984 56324
rect 20036 56312 20042 56364
rect 22373 56355 22431 56361
rect 22373 56321 22385 56355
rect 22419 56352 22431 56355
rect 22462 56352 22468 56364
rect 22419 56324 22468 56352
rect 22419 56321 22431 56324
rect 22373 56315 22431 56321
rect 22462 56312 22468 56324
rect 22520 56312 22526 56364
rect 24480 56355 24538 56361
rect 24480 56321 24492 56355
rect 24526 56352 24538 56355
rect 25038 56352 25044 56364
rect 24526 56324 25044 56352
rect 24526 56321 24538 56324
rect 24480 56315 24538 56321
rect 25038 56312 25044 56324
rect 25096 56312 25102 56364
rect 28350 56312 28356 56364
rect 28408 56352 28414 56364
rect 30449 56355 30507 56361
rect 30449 56352 30461 56355
rect 28408 56324 30461 56352
rect 28408 56312 28414 56324
rect 30449 56321 30461 56324
rect 30495 56321 30507 56355
rect 32858 56352 32864 56364
rect 32819 56324 32864 56352
rect 30449 56315 30507 56321
rect 32858 56312 32864 56324
rect 32916 56312 32922 56364
rect 33128 56355 33186 56361
rect 33128 56321 33140 56355
rect 33174 56352 33186 56355
rect 33174 56324 35894 56352
rect 33174 56321 33186 56324
rect 33128 56315 33186 56321
rect 3605 56287 3663 56293
rect 3605 56253 3617 56287
rect 3651 56253 3663 56287
rect 3605 56247 3663 56253
rect 3620 56148 3648 56247
rect 6914 56244 6920 56296
rect 6972 56284 6978 56296
rect 14645 56287 14703 56293
rect 6972 56256 7017 56284
rect 6972 56244 6978 56256
rect 14645 56253 14657 56287
rect 14691 56284 14703 56287
rect 14737 56287 14795 56293
rect 14737 56284 14749 56287
rect 14691 56256 14749 56284
rect 14691 56253 14703 56256
rect 14645 56247 14703 56253
rect 14737 56253 14749 56256
rect 14783 56253 14795 56287
rect 14737 56247 14795 56253
rect 17862 56244 17868 56296
rect 17920 56284 17926 56296
rect 18049 56287 18107 56293
rect 18049 56284 18061 56287
rect 17920 56256 18061 56284
rect 17920 56244 17926 56256
rect 18049 56253 18061 56256
rect 18095 56253 18107 56287
rect 18049 56247 18107 56253
rect 24213 56287 24271 56293
rect 24213 56253 24225 56287
rect 24259 56253 24271 56287
rect 24213 56247 24271 56253
rect 19242 56176 19248 56228
rect 19300 56216 19306 56228
rect 19429 56219 19487 56225
rect 19429 56216 19441 56219
rect 19300 56188 19441 56216
rect 19300 56176 19306 56188
rect 19429 56185 19441 56188
rect 19475 56185 19487 56219
rect 19429 56179 19487 56185
rect 3878 56148 3884 56160
rect 3620 56120 3884 56148
rect 3878 56108 3884 56120
rect 3936 56108 3942 56160
rect 10134 56148 10140 56160
rect 10095 56120 10140 56148
rect 10134 56108 10140 56120
rect 10192 56108 10198 56160
rect 14182 56148 14188 56160
rect 14143 56120 14188 56148
rect 14182 56108 14188 56120
rect 14240 56108 14246 56160
rect 16114 56148 16120 56160
rect 16075 56120 16120 56148
rect 16114 56108 16120 56120
rect 16172 56108 16178 56160
rect 21266 56148 21272 56160
rect 21227 56120 21272 56148
rect 21266 56108 21272 56120
rect 21324 56108 21330 56160
rect 21726 56108 21732 56160
rect 21784 56148 21790 56160
rect 24228 56148 24256 56247
rect 28258 56244 28264 56296
rect 28316 56284 28322 56296
rect 30193 56287 30251 56293
rect 30193 56284 30205 56287
rect 28316 56256 30205 56284
rect 28316 56244 28322 56256
rect 30193 56253 30205 56256
rect 30239 56253 30251 56287
rect 34698 56284 34704 56296
rect 34611 56256 34704 56284
rect 30193 56247 30251 56253
rect 34698 56244 34704 56256
rect 34756 56244 34762 56296
rect 25590 56148 25596 56160
rect 21784 56120 24256 56148
rect 25551 56120 25596 56148
rect 21784 56108 21790 56120
rect 25590 56108 25596 56120
rect 25648 56108 25654 56160
rect 29178 56108 29184 56160
rect 29236 56148 29242 56160
rect 29273 56151 29331 56157
rect 29273 56148 29285 56151
rect 29236 56120 29285 56148
rect 29236 56108 29242 56120
rect 29273 56117 29285 56120
rect 29319 56117 29331 56151
rect 29273 56111 29331 56117
rect 30374 56108 30380 56160
rect 30432 56148 30438 56160
rect 31573 56151 31631 56157
rect 31573 56148 31585 56151
rect 30432 56120 31585 56148
rect 30432 56108 30438 56120
rect 31573 56117 31585 56120
rect 31619 56117 31631 56151
rect 34716 56148 34744 56244
rect 35866 56216 35894 56324
rect 37274 56312 37280 56364
rect 37332 56352 37338 56364
rect 37642 56352 37648 56364
rect 37332 56324 37648 56352
rect 37332 56312 37338 56324
rect 37642 56312 37648 56324
rect 37700 56312 37706 56364
rect 37912 56355 37970 56361
rect 37912 56321 37924 56355
rect 37958 56352 37970 56355
rect 39022 56352 39028 56364
rect 37958 56324 39028 56352
rect 37958 56321 37970 56324
rect 37912 56315 37970 56321
rect 39022 56312 39028 56324
rect 39080 56312 39086 56364
rect 40402 56352 40408 56364
rect 40363 56324 40408 56352
rect 40402 56312 40408 56324
rect 40460 56312 40466 56364
rect 41874 56312 41880 56364
rect 41932 56352 41938 56364
rect 42685 56355 42743 56361
rect 42685 56352 42697 56355
rect 41932 56324 42697 56352
rect 41932 56312 41938 56324
rect 42685 56321 42697 56324
rect 42731 56321 42743 56355
rect 48958 56352 48964 56364
rect 48871 56324 48964 56352
rect 42685 56315 42743 56321
rect 48958 56312 48964 56324
rect 49016 56352 49022 56364
rect 50801 56355 50859 56361
rect 50801 56352 50813 56355
rect 49016 56324 50813 56352
rect 49016 56312 49022 56324
rect 50801 56321 50813 56324
rect 50847 56321 50859 56355
rect 50801 56315 50859 56321
rect 42429 56287 42487 56293
rect 42429 56253 42441 56287
rect 42475 56253 42487 56287
rect 42429 56247 42487 56253
rect 44269 56287 44327 56293
rect 44269 56253 44281 56287
rect 44315 56253 44327 56287
rect 44269 56247 44327 56253
rect 36081 56219 36139 56225
rect 36081 56216 36093 56219
rect 35866 56188 36093 56216
rect 36081 56185 36093 56188
rect 36127 56185 36139 56219
rect 36081 56179 36139 56185
rect 35342 56148 35348 56160
rect 34716 56120 35348 56148
rect 31573 56111 31631 56117
rect 35342 56108 35348 56120
rect 35400 56108 35406 56160
rect 42444 56148 42472 56247
rect 42794 56148 42800 56160
rect 42444 56120 42800 56148
rect 42794 56108 42800 56120
rect 42852 56148 42858 56160
rect 44284 56148 44312 56247
rect 53374 56244 53380 56296
rect 53432 56284 53438 56296
rect 54312 56293 54340 56392
rect 55122 56380 55128 56392
rect 55180 56380 55186 56432
rect 54564 56355 54622 56361
rect 54564 56321 54576 56355
rect 54610 56352 54622 56355
rect 55950 56352 55956 56364
rect 54610 56324 55956 56352
rect 54610 56321 54622 56324
rect 54564 56315 54622 56321
rect 55950 56312 55956 56324
rect 56008 56312 56014 56364
rect 54297 56287 54355 56293
rect 54297 56284 54309 56287
rect 53432 56256 54309 56284
rect 53432 56244 53438 56256
rect 54297 56253 54309 56256
rect 54343 56253 54355 56287
rect 54297 56247 54355 56253
rect 51902 56176 51908 56228
rect 51960 56216 51966 56228
rect 52181 56219 52239 56225
rect 52181 56216 52193 56219
rect 51960 56188 52193 56216
rect 51960 56176 51966 56188
rect 52181 56185 52193 56188
rect 52227 56185 52239 56219
rect 52181 56179 52239 56185
rect 42852 56120 44312 56148
rect 42852 56108 42858 56120
rect 1104 56058 59340 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 59340 56058
rect 1104 55984 59340 56006
rect 20622 55904 20628 55956
rect 20680 55944 20686 55956
rect 21269 55947 21327 55953
rect 21269 55944 21281 55947
rect 20680 55916 21281 55944
rect 20680 55904 20686 55916
rect 21269 55913 21281 55916
rect 21315 55913 21327 55947
rect 28534 55944 28540 55956
rect 28495 55916 28540 55944
rect 21269 55907 21327 55913
rect 28534 55904 28540 55916
rect 28592 55904 28598 55956
rect 39022 55944 39028 55956
rect 38983 55916 39028 55944
rect 39022 55904 39028 55916
rect 39080 55904 39086 55956
rect 42794 55904 42800 55956
rect 42852 55944 42858 55956
rect 43070 55944 43076 55956
rect 42852 55916 43076 55944
rect 42852 55904 42858 55916
rect 43070 55904 43076 55916
rect 43128 55944 43134 55956
rect 43165 55947 43223 55953
rect 43165 55944 43177 55947
rect 43128 55916 43177 55944
rect 43128 55904 43134 55916
rect 43165 55913 43177 55916
rect 43211 55913 43223 55947
rect 43165 55907 43223 55913
rect 46290 55904 46296 55956
rect 46348 55944 46354 55956
rect 46385 55947 46443 55953
rect 46385 55944 46397 55947
rect 46348 55916 46397 55944
rect 46348 55904 46354 55916
rect 46385 55913 46397 55916
rect 46431 55913 46443 55947
rect 46385 55907 46443 55913
rect 49326 55904 49332 55956
rect 49384 55944 49390 55956
rect 49421 55947 49479 55953
rect 49421 55944 49433 55947
rect 49384 55916 49433 55944
rect 49384 55904 49390 55916
rect 49421 55913 49433 55916
rect 49467 55913 49479 55947
rect 49421 55907 49479 55913
rect 54757 55947 54815 55953
rect 54757 55913 54769 55947
rect 54803 55944 54815 55947
rect 56778 55944 56784 55956
rect 54803 55916 56784 55944
rect 54803 55913 54815 55916
rect 54757 55907 54815 55913
rect 56778 55904 56784 55916
rect 56836 55904 56842 55956
rect 8938 55808 8944 55820
rect 8899 55780 8944 55808
rect 8938 55768 8944 55780
rect 8996 55768 9002 55820
rect 14090 55768 14096 55820
rect 14148 55808 14154 55820
rect 14645 55811 14703 55817
rect 14645 55808 14657 55811
rect 14148 55780 14657 55808
rect 14148 55768 14154 55780
rect 14645 55777 14657 55780
rect 14691 55777 14703 55811
rect 37642 55808 37648 55820
rect 37603 55780 37648 55808
rect 14645 55771 14703 55777
rect 37642 55768 37648 55780
rect 37700 55768 37706 55820
rect 45002 55808 45008 55820
rect 44963 55780 45008 55808
rect 45002 55768 45008 55780
rect 45060 55768 45066 55820
rect 4985 55675 5043 55681
rect 4985 55641 4997 55675
rect 5031 55672 5043 55675
rect 5534 55672 5540 55684
rect 5031 55644 5540 55672
rect 5031 55641 5043 55644
rect 4985 55635 5043 55641
rect 5534 55632 5540 55644
rect 5592 55672 5598 55684
rect 8754 55672 8760 55684
rect 5592 55644 8760 55672
rect 5592 55632 5598 55644
rect 8754 55632 8760 55644
rect 8812 55632 8818 55684
rect 8956 55672 8984 55768
rect 9208 55743 9266 55749
rect 9208 55709 9220 55743
rect 9254 55740 9266 55743
rect 10134 55740 10140 55752
rect 9254 55712 10140 55740
rect 9254 55709 9266 55712
rect 9208 55703 9266 55709
rect 10134 55700 10140 55712
rect 10192 55700 10198 55752
rect 11698 55700 11704 55752
rect 11756 55740 11762 55752
rect 12161 55743 12219 55749
rect 12161 55740 12173 55743
rect 11756 55712 12173 55740
rect 11756 55700 11762 55712
rect 12161 55709 12173 55712
rect 12207 55709 12219 55743
rect 12161 55703 12219 55709
rect 14912 55743 14970 55749
rect 14912 55709 14924 55743
rect 14958 55740 14970 55743
rect 16114 55740 16120 55752
rect 14958 55712 16120 55740
rect 14958 55709 14970 55712
rect 14912 55703 14970 55709
rect 16114 55700 16120 55712
rect 16172 55700 16178 55752
rect 17313 55743 17371 55749
rect 17313 55709 17325 55743
rect 17359 55709 17371 55743
rect 17313 55703 17371 55709
rect 17580 55743 17638 55749
rect 17580 55709 17592 55743
rect 17626 55740 17638 55743
rect 18690 55740 18696 55752
rect 17626 55712 18696 55740
rect 17626 55709 17638 55712
rect 17580 55703 17638 55709
rect 9306 55672 9312 55684
rect 8956 55644 9312 55672
rect 9306 55632 9312 55644
rect 9364 55632 9370 55684
rect 12428 55675 12486 55681
rect 12428 55641 12440 55675
rect 12474 55672 12486 55675
rect 13722 55672 13728 55684
rect 12474 55644 13728 55672
rect 12474 55641 12486 55644
rect 12428 55635 12486 55641
rect 13722 55632 13728 55644
rect 13780 55632 13786 55684
rect 17328 55672 17356 55703
rect 18690 55700 18696 55712
rect 18748 55700 18754 55752
rect 19889 55743 19947 55749
rect 19889 55709 19901 55743
rect 19935 55740 19947 55743
rect 19978 55740 19984 55752
rect 19935 55712 19984 55740
rect 19935 55709 19947 55712
rect 19889 55703 19947 55709
rect 19978 55700 19984 55712
rect 20036 55700 20042 55752
rect 20156 55743 20214 55749
rect 20156 55709 20168 55743
rect 20202 55740 20214 55743
rect 21266 55740 21272 55752
rect 20202 55712 21272 55740
rect 20202 55709 20214 55712
rect 20156 55703 20214 55709
rect 21266 55700 21272 55712
rect 21324 55700 21330 55752
rect 21726 55740 21732 55752
rect 21639 55712 21732 55740
rect 21726 55700 21732 55712
rect 21784 55700 21790 55752
rect 21818 55700 21824 55752
rect 21876 55740 21882 55752
rect 22462 55740 22468 55752
rect 21876 55712 22468 55740
rect 21876 55700 21882 55712
rect 22462 55700 22468 55712
rect 22520 55740 22526 55752
rect 23658 55740 23664 55752
rect 22520 55712 23664 55740
rect 22520 55700 22526 55712
rect 23658 55700 23664 55712
rect 23716 55740 23722 55752
rect 24394 55740 24400 55752
rect 23716 55712 24400 55740
rect 23716 55700 23722 55712
rect 24394 55700 24400 55712
rect 24452 55700 24458 55752
rect 26970 55700 26976 55752
rect 27028 55740 27034 55752
rect 27157 55743 27215 55749
rect 27157 55740 27169 55743
rect 27028 55712 27169 55740
rect 27028 55700 27034 55712
rect 27157 55709 27169 55712
rect 27203 55709 27215 55743
rect 27157 55703 27215 55709
rect 27246 55700 27252 55752
rect 27304 55740 27310 55752
rect 27413 55743 27471 55749
rect 27413 55740 27425 55743
rect 27304 55712 27425 55740
rect 27304 55700 27310 55712
rect 27413 55709 27425 55712
rect 27459 55709 27471 55743
rect 32122 55740 32128 55752
rect 32035 55712 32128 55740
rect 27413 55703 27471 55709
rect 32122 55700 32128 55712
rect 32180 55740 32186 55752
rect 32766 55740 32772 55752
rect 32180 55712 32772 55740
rect 32180 55700 32186 55712
rect 32766 55700 32772 55712
rect 32824 55700 32830 55752
rect 35342 55700 35348 55752
rect 35400 55740 35406 55752
rect 35805 55743 35863 55749
rect 35805 55740 35817 55743
rect 35400 55712 35817 55740
rect 35400 55700 35406 55712
rect 35805 55709 35817 55712
rect 35851 55709 35863 55743
rect 35805 55703 35863 55709
rect 40037 55743 40095 55749
rect 40037 55709 40049 55743
rect 40083 55740 40095 55743
rect 40126 55740 40132 55752
rect 40083 55712 40132 55740
rect 40083 55709 40095 55712
rect 40037 55703 40095 55709
rect 40126 55700 40132 55712
rect 40184 55700 40190 55752
rect 40304 55743 40362 55749
rect 40304 55709 40316 55743
rect 40350 55740 40362 55743
rect 42334 55740 42340 55752
rect 40350 55712 42340 55740
rect 40350 55709 40362 55712
rect 40304 55703 40362 55709
rect 42334 55700 42340 55712
rect 42392 55700 42398 55752
rect 17862 55672 17868 55684
rect 17328 55644 17868 55672
rect 17862 55632 17868 55644
rect 17920 55632 17926 55684
rect 19996 55672 20024 55700
rect 21744 55672 21772 55700
rect 19996 55644 21772 55672
rect 21996 55675 22054 55681
rect 21996 55641 22008 55675
rect 22042 55672 22054 55675
rect 23198 55672 23204 55684
rect 22042 55644 23204 55672
rect 22042 55641 22054 55644
rect 21996 55635 22054 55641
rect 23198 55632 23204 55644
rect 23256 55632 23262 55684
rect 24664 55675 24722 55681
rect 24664 55641 24676 55675
rect 24710 55672 24722 55675
rect 25406 55672 25412 55684
rect 24710 55644 25412 55672
rect 24710 55641 24722 55644
rect 24664 55635 24722 55641
rect 25406 55632 25412 55644
rect 25464 55632 25470 55684
rect 32392 55675 32450 55681
rect 32392 55641 32404 55675
rect 32438 55672 32450 55675
rect 33134 55672 33140 55684
rect 32438 55644 33140 55672
rect 32438 55641 32450 55644
rect 32392 55635 32450 55641
rect 33134 55632 33140 55644
rect 33192 55632 33198 55684
rect 36072 55675 36130 55681
rect 36072 55641 36084 55675
rect 36118 55672 36130 55675
rect 36722 55672 36728 55684
rect 36118 55644 36728 55672
rect 36118 55641 36130 55644
rect 36072 55635 36130 55641
rect 36722 55632 36728 55644
rect 36780 55632 36786 55684
rect 37890 55675 37948 55681
rect 37890 55672 37902 55675
rect 37200 55644 37902 55672
rect 6270 55604 6276 55616
rect 6231 55576 6276 55604
rect 6270 55564 6276 55576
rect 6328 55564 6334 55616
rect 10318 55604 10324 55616
rect 10279 55576 10324 55604
rect 10318 55564 10324 55576
rect 10376 55564 10382 55616
rect 13541 55607 13599 55613
rect 13541 55573 13553 55607
rect 13587 55604 13599 55607
rect 14366 55604 14372 55616
rect 13587 55576 14372 55604
rect 13587 55573 13599 55576
rect 13541 55567 13599 55573
rect 14366 55564 14372 55576
rect 14424 55564 14430 55616
rect 16022 55604 16028 55616
rect 15983 55576 16028 55604
rect 16022 55564 16028 55576
rect 16080 55564 16086 55616
rect 18690 55604 18696 55616
rect 18651 55576 18696 55604
rect 18690 55564 18696 55576
rect 18748 55564 18754 55616
rect 23109 55607 23167 55613
rect 23109 55573 23121 55607
rect 23155 55604 23167 55607
rect 23842 55604 23848 55616
rect 23155 55576 23848 55604
rect 23155 55573 23167 55576
rect 23109 55567 23167 55573
rect 23842 55564 23848 55576
rect 23900 55564 23906 55616
rect 25777 55607 25835 55613
rect 25777 55573 25789 55607
rect 25823 55604 25835 55607
rect 28350 55604 28356 55616
rect 25823 55576 28356 55604
rect 25823 55573 25835 55576
rect 25777 55567 25835 55573
rect 28350 55564 28356 55576
rect 28408 55564 28414 55616
rect 33502 55604 33508 55616
rect 33463 55576 33508 55604
rect 33502 55564 33508 55576
rect 33560 55564 33566 55616
rect 37200 55613 37228 55644
rect 37890 55641 37902 55644
rect 37936 55641 37948 55675
rect 37890 55635 37948 55641
rect 41782 55632 41788 55684
rect 41840 55672 41846 55684
rect 41877 55675 41935 55681
rect 41877 55672 41889 55675
rect 41840 55644 41889 55672
rect 41840 55632 41846 55644
rect 41877 55641 41889 55644
rect 41923 55641 41935 55675
rect 45020 55672 45048 55768
rect 45272 55743 45330 55749
rect 45272 55709 45284 55743
rect 45318 55740 45330 55743
rect 45554 55740 45560 55752
rect 45318 55712 45560 55740
rect 45318 55709 45330 55712
rect 45272 55703 45330 55709
rect 45554 55700 45560 55712
rect 45612 55700 45618 55752
rect 48314 55749 48320 55752
rect 48041 55743 48099 55749
rect 48041 55709 48053 55743
rect 48087 55709 48099 55743
rect 48308 55740 48320 55749
rect 48275 55712 48320 55740
rect 48041 55703 48099 55709
rect 48308 55703 48320 55712
rect 48056 55672 48084 55703
rect 48314 55700 48320 55703
rect 48372 55700 48378 55752
rect 50154 55740 50160 55752
rect 50115 55712 50160 55740
rect 50154 55700 50160 55712
rect 50212 55700 50218 55752
rect 52730 55700 52736 55752
rect 52788 55740 52794 55752
rect 53374 55740 53380 55752
rect 52788 55712 53380 55740
rect 52788 55700 52794 55712
rect 53374 55700 53380 55712
rect 53432 55700 53438 55752
rect 53644 55743 53702 55749
rect 53644 55709 53656 55743
rect 53690 55740 53702 55743
rect 56594 55740 56600 55752
rect 53690 55712 56600 55740
rect 53690 55709 53702 55712
rect 53644 55703 53702 55709
rect 56594 55700 56600 55712
rect 56652 55700 56658 55752
rect 45020 55644 48084 55672
rect 50424 55675 50482 55681
rect 41877 55635 41935 55641
rect 50424 55641 50436 55675
rect 50470 55672 50482 55675
rect 51166 55672 51172 55684
rect 50470 55644 51172 55672
rect 50470 55641 50482 55644
rect 50424 55635 50482 55641
rect 51166 55632 51172 55644
rect 51224 55632 51230 55684
rect 56134 55672 56140 55684
rect 56095 55644 56140 55672
rect 56134 55632 56140 55644
rect 56192 55632 56198 55684
rect 37185 55607 37243 55613
rect 37185 55573 37197 55607
rect 37231 55573 37243 55607
rect 41414 55604 41420 55616
rect 41375 55576 41420 55604
rect 37185 55567 37243 55573
rect 41414 55564 41420 55576
rect 41472 55564 41478 55616
rect 51534 55604 51540 55616
rect 51495 55576 51540 55604
rect 51534 55564 51540 55576
rect 51592 55564 51598 55616
rect 57054 55564 57060 55616
rect 57112 55604 57118 55616
rect 57425 55607 57483 55613
rect 57425 55604 57437 55607
rect 57112 55576 57437 55604
rect 57112 55564 57118 55576
rect 57425 55573 57437 55576
rect 57471 55573 57483 55607
rect 57425 55567 57483 55573
rect 1104 55514 59340 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 59340 55514
rect 1104 55440 59340 55462
rect 5166 55400 5172 55412
rect 5127 55372 5172 55400
rect 5166 55360 5172 55372
rect 5224 55360 5230 55412
rect 8202 55400 8208 55412
rect 8163 55372 8208 55400
rect 8202 55360 8208 55372
rect 8260 55360 8266 55412
rect 13722 55400 13728 55412
rect 13683 55372 13728 55400
rect 13722 55360 13728 55372
rect 13780 55360 13786 55412
rect 15562 55400 15568 55412
rect 15523 55372 15568 55400
rect 15562 55360 15568 55372
rect 15620 55360 15626 55412
rect 19150 55400 19156 55412
rect 19111 55372 19156 55400
rect 19150 55360 19156 55372
rect 19208 55360 19214 55412
rect 20990 55400 20996 55412
rect 20951 55372 20996 55400
rect 20990 55360 20996 55372
rect 21048 55360 21054 55412
rect 23198 55400 23204 55412
rect 23159 55372 23204 55400
rect 23198 55360 23204 55372
rect 23256 55360 23262 55412
rect 25038 55400 25044 55412
rect 24999 55372 25044 55400
rect 25038 55360 25044 55372
rect 25096 55360 25102 55412
rect 29822 55360 29828 55412
rect 29880 55400 29886 55412
rect 30561 55403 30619 55409
rect 30561 55400 30573 55403
rect 29880 55372 30573 55400
rect 29880 55360 29886 55372
rect 30561 55369 30573 55372
rect 30607 55369 30619 55403
rect 30561 55363 30619 55369
rect 32398 55360 32404 55412
rect 32456 55400 32462 55412
rect 33505 55403 33563 55409
rect 33505 55400 33517 55403
rect 32456 55372 33517 55400
rect 32456 55360 32462 55372
rect 33505 55369 33517 55372
rect 33551 55369 33563 55403
rect 36722 55400 36728 55412
rect 36683 55372 36728 55400
rect 33505 55363 33563 55369
rect 36722 55360 36728 55372
rect 36780 55360 36786 55412
rect 38930 55360 38936 55412
rect 38988 55400 38994 55412
rect 40037 55403 40095 55409
rect 40037 55400 40049 55403
rect 38988 55372 40049 55400
rect 38988 55360 38994 55372
rect 40037 55369 40049 55372
rect 40083 55369 40095 55403
rect 41874 55400 41880 55412
rect 41835 55372 41880 55400
rect 40037 55363 40095 55369
rect 41874 55360 41880 55372
rect 41932 55360 41938 55412
rect 49421 55403 49479 55409
rect 49421 55369 49433 55403
rect 49467 55400 49479 55403
rect 49694 55400 49700 55412
rect 49467 55372 49700 55400
rect 49467 55369 49479 55372
rect 49421 55363 49479 55369
rect 49694 55360 49700 55372
rect 49752 55360 49758 55412
rect 52546 55360 52552 55412
rect 52604 55400 52610 55412
rect 54113 55403 54171 55409
rect 54113 55400 54125 55403
rect 52604 55372 54125 55400
rect 52604 55360 52610 55372
rect 54113 55369 54125 55372
rect 54159 55369 54171 55403
rect 55950 55400 55956 55412
rect 55911 55372 55956 55400
rect 54113 55363 54171 55369
rect 55950 55360 55956 55372
rect 56008 55360 56014 55412
rect 4056 55335 4114 55341
rect 4056 55301 4068 55335
rect 4102 55332 4114 55335
rect 8386 55332 8392 55344
rect 4102 55304 8392 55332
rect 4102 55301 4114 55304
rect 4056 55295 4114 55301
rect 8386 55292 8392 55304
rect 8444 55292 8450 55344
rect 9576 55335 9634 55341
rect 9576 55301 9588 55335
rect 9622 55332 9634 55335
rect 10318 55332 10324 55344
rect 9622 55304 10324 55332
rect 9622 55301 9634 55304
rect 9576 55295 9634 55301
rect 10318 55292 10324 55304
rect 10376 55292 10382 55344
rect 12612 55335 12670 55341
rect 12612 55301 12624 55335
rect 12658 55332 12670 55335
rect 14182 55332 14188 55344
rect 12658 55304 14188 55332
rect 12658 55301 12670 55304
rect 12612 55295 12670 55301
rect 14182 55292 14188 55304
rect 14240 55292 14246 55344
rect 14452 55335 14510 55341
rect 14452 55301 14464 55335
rect 14498 55332 14510 55335
rect 16022 55332 16028 55344
rect 14498 55304 16028 55332
rect 14498 55301 14510 55304
rect 14452 55295 14510 55301
rect 16022 55292 16028 55304
rect 16080 55292 16086 55344
rect 18040 55335 18098 55341
rect 18040 55301 18052 55335
rect 18086 55332 18098 55335
rect 18690 55332 18696 55344
rect 18086 55304 18696 55332
rect 18086 55301 18098 55304
rect 18040 55295 18098 55301
rect 18690 55292 18696 55304
rect 18748 55292 18754 55344
rect 19334 55292 19340 55344
rect 19392 55332 19398 55344
rect 19858 55335 19916 55341
rect 19858 55332 19870 55335
rect 19392 55304 19870 55332
rect 19392 55292 19398 55304
rect 19858 55301 19870 55304
rect 19904 55301 19916 55335
rect 19858 55295 19916 55301
rect 19978 55292 19984 55344
rect 20036 55292 20042 55344
rect 24394 55292 24400 55344
rect 24452 55332 24458 55344
rect 28258 55332 28264 55344
rect 24452 55304 28264 55332
rect 24452 55292 24458 55304
rect 28258 55292 28264 55304
rect 28316 55292 28322 55344
rect 40126 55332 40132 55344
rect 38672 55304 40132 55332
rect 3789 55267 3847 55273
rect 3789 55233 3801 55267
rect 3835 55264 3847 55267
rect 3878 55264 3884 55276
rect 3835 55236 3884 55264
rect 3835 55233 3847 55236
rect 3789 55227 3847 55233
rect 3878 55224 3884 55236
rect 3936 55224 3942 55276
rect 6825 55267 6883 55273
rect 6825 55233 6837 55267
rect 6871 55264 6883 55267
rect 6914 55264 6920 55276
rect 6871 55236 6920 55264
rect 6871 55233 6883 55236
rect 6825 55227 6883 55233
rect 6914 55224 6920 55236
rect 6972 55224 6978 55276
rect 7092 55267 7150 55273
rect 7092 55233 7104 55267
rect 7138 55264 7150 55267
rect 7926 55264 7932 55276
rect 7138 55236 7932 55264
rect 7138 55233 7150 55236
rect 7092 55227 7150 55233
rect 7926 55224 7932 55236
rect 7984 55224 7990 55276
rect 12345 55267 12403 55273
rect 12345 55233 12357 55267
rect 12391 55264 12403 55267
rect 17773 55267 17831 55273
rect 12391 55236 14136 55264
rect 12391 55233 12403 55236
rect 12345 55227 12403 55233
rect 14108 55208 14136 55236
rect 17773 55233 17785 55267
rect 17819 55264 17831 55267
rect 17862 55264 17868 55276
rect 17819 55236 17868 55264
rect 17819 55233 17831 55236
rect 17773 55227 17831 55233
rect 17862 55224 17868 55236
rect 17920 55224 17926 55276
rect 19613 55267 19671 55273
rect 19613 55233 19625 55267
rect 19659 55264 19671 55267
rect 19996 55264 20024 55292
rect 19659 55236 20024 55264
rect 22088 55267 22146 55273
rect 19659 55233 19671 55236
rect 19613 55227 19671 55233
rect 22088 55233 22100 55267
rect 22134 55264 22146 55267
rect 23106 55264 23112 55276
rect 22134 55236 23112 55264
rect 22134 55233 22146 55236
rect 22088 55227 22146 55233
rect 23106 55224 23112 55236
rect 23164 55224 23170 55276
rect 23658 55264 23664 55276
rect 23619 55236 23664 55264
rect 23658 55224 23664 55236
rect 23716 55224 23722 55276
rect 23928 55267 23986 55273
rect 23928 55233 23940 55267
rect 23974 55264 23986 55267
rect 25038 55264 25044 55276
rect 23974 55236 25044 55264
rect 23974 55233 23986 55236
rect 23928 55227 23986 55233
rect 25038 55224 25044 55236
rect 25096 55224 25102 55276
rect 27608 55267 27666 55273
rect 27608 55233 27620 55267
rect 27654 55264 27666 55267
rect 28166 55264 28172 55276
rect 27654 55236 28172 55264
rect 27654 55233 27666 55236
rect 27608 55227 27666 55233
rect 28166 55224 28172 55236
rect 28224 55224 28230 55276
rect 29270 55264 29276 55276
rect 28736 55236 29276 55264
rect 9306 55196 9312 55208
rect 9219 55168 9312 55196
rect 9306 55156 9312 55168
rect 9364 55156 9370 55208
rect 14090 55156 14096 55208
rect 14148 55196 14154 55208
rect 14185 55199 14243 55205
rect 14185 55196 14197 55199
rect 14148 55168 14197 55196
rect 14148 55156 14154 55168
rect 14185 55165 14197 55168
rect 14231 55165 14243 55199
rect 21818 55196 21824 55208
rect 21779 55168 21824 55196
rect 14185 55159 14243 55165
rect 21818 55156 21824 55168
rect 21876 55156 21882 55208
rect 27341 55199 27399 55205
rect 27341 55165 27353 55199
rect 27387 55165 27399 55199
rect 27341 55159 27399 55165
rect 7006 55020 7012 55072
rect 7064 55060 7070 55072
rect 9315 55060 9343 55156
rect 10686 55060 10692 55072
rect 7064 55032 9343 55060
rect 10647 55032 10692 55060
rect 7064 55020 7070 55032
rect 10686 55020 10692 55032
rect 10744 55020 10750 55072
rect 26970 55020 26976 55072
rect 27028 55060 27034 55072
rect 27356 55060 27384 55159
rect 28736 55137 28764 55236
rect 29270 55224 29276 55236
rect 29328 55224 29334 55276
rect 29448 55267 29506 55273
rect 29448 55233 29460 55267
rect 29494 55264 29506 55267
rect 30190 55264 30196 55276
rect 29494 55236 30196 55264
rect 29494 55233 29506 55236
rect 29448 55227 29506 55233
rect 30190 55224 30196 55236
rect 30248 55224 30254 55276
rect 32392 55267 32450 55273
rect 32392 55233 32404 55267
rect 32438 55264 32450 55267
rect 33410 55264 33416 55276
rect 32438 55236 33416 55264
rect 32438 55233 32450 55236
rect 32392 55227 32450 55233
rect 33410 55224 33416 55236
rect 33468 55224 33474 55276
rect 35342 55264 35348 55276
rect 35303 55236 35348 55264
rect 35342 55224 35348 55236
rect 35400 55224 35406 55276
rect 35612 55267 35670 55273
rect 35612 55233 35624 55267
rect 35658 55264 35670 55267
rect 36630 55264 36636 55276
rect 35658 55236 36636 55264
rect 35658 55233 35670 55236
rect 35612 55227 35670 55233
rect 36630 55224 36636 55236
rect 36688 55224 36694 55276
rect 38672 55273 38700 55304
rect 40126 55292 40132 55304
rect 40184 55332 40190 55344
rect 40494 55332 40500 55344
rect 40184 55304 40500 55332
rect 40184 55292 40190 55304
rect 40494 55292 40500 55304
rect 40552 55292 40558 55344
rect 40764 55335 40822 55341
rect 40764 55301 40776 55335
rect 40810 55332 40822 55335
rect 41414 55332 41420 55344
rect 40810 55304 41420 55332
rect 40810 55301 40822 55304
rect 40764 55295 40822 55301
rect 41414 55292 41420 55304
rect 41472 55292 41478 55344
rect 45364 55335 45422 55341
rect 45364 55301 45376 55335
rect 45410 55332 45422 55335
rect 46382 55332 46388 55344
rect 45410 55304 46388 55332
rect 45410 55301 45422 55304
rect 45364 55295 45422 55301
rect 46382 55292 46388 55304
rect 46440 55292 46446 55344
rect 48056 55304 49924 55332
rect 38657 55267 38715 55273
rect 38657 55233 38669 55267
rect 38703 55233 38715 55267
rect 38657 55227 38715 55233
rect 38924 55267 38982 55273
rect 38924 55233 38936 55267
rect 38970 55264 38982 55267
rect 41322 55264 41328 55276
rect 38970 55236 41328 55264
rect 38970 55233 38982 55236
rect 38924 55227 38982 55233
rect 41322 55224 41328 55236
rect 41380 55224 41386 55276
rect 45097 55267 45155 55273
rect 45097 55233 45109 55267
rect 45143 55264 45155 55267
rect 45186 55264 45192 55276
rect 45143 55236 45192 55264
rect 45143 55233 45155 55236
rect 45097 55227 45155 55233
rect 45186 55224 45192 55236
rect 45244 55224 45250 55276
rect 29178 55196 29184 55208
rect 29091 55168 29184 55196
rect 29178 55156 29184 55168
rect 29236 55156 29242 55208
rect 32122 55196 32128 55208
rect 32083 55168 32128 55196
rect 32122 55156 32128 55168
rect 32180 55156 32186 55208
rect 40494 55196 40500 55208
rect 40455 55168 40500 55196
rect 40494 55156 40500 55168
rect 40552 55156 40558 55208
rect 47578 55156 47584 55208
rect 47636 55196 47642 55208
rect 48056 55205 48084 55304
rect 48308 55267 48366 55273
rect 48308 55233 48320 55267
rect 48354 55264 48366 55267
rect 49050 55264 49056 55276
rect 48354 55236 49056 55264
rect 48354 55233 48366 55236
rect 48308 55227 48366 55233
rect 49050 55224 49056 55236
rect 49108 55224 49114 55276
rect 49896 55273 49924 55304
rect 51534 55292 51540 55344
rect 51592 55332 51598 55344
rect 52978 55335 53036 55341
rect 52978 55332 52990 55335
rect 51592 55304 52990 55332
rect 51592 55292 51598 55304
rect 52978 55301 52990 55304
rect 53024 55301 53036 55335
rect 52978 55295 53036 55301
rect 49881 55267 49939 55273
rect 49881 55233 49893 55267
rect 49927 55233 49939 55267
rect 49881 55227 49939 55233
rect 50148 55267 50206 55273
rect 50148 55233 50160 55267
rect 50194 55264 50206 55267
rect 50890 55264 50896 55276
rect 50194 55236 50896 55264
rect 50194 55233 50206 55236
rect 50148 55227 50206 55233
rect 50890 55224 50896 55236
rect 50948 55224 50954 55276
rect 52638 55224 52644 55276
rect 52696 55264 52702 55276
rect 52733 55267 52791 55273
rect 52733 55264 52745 55267
rect 52696 55236 52745 55264
rect 52696 55224 52702 55236
rect 52733 55233 52745 55236
rect 52779 55233 52791 55267
rect 52733 55227 52791 55233
rect 54573 55267 54631 55273
rect 54573 55233 54585 55267
rect 54619 55233 54631 55267
rect 54573 55227 54631 55233
rect 54840 55267 54898 55273
rect 54840 55233 54852 55267
rect 54886 55264 54898 55267
rect 56134 55264 56140 55276
rect 54886 55236 56140 55264
rect 54886 55233 54898 55236
rect 54840 55227 54898 55233
rect 48041 55199 48099 55205
rect 48041 55196 48053 55199
rect 47636 55168 48053 55196
rect 47636 55156 47642 55168
rect 48041 55165 48053 55168
rect 48087 55165 48099 55199
rect 48041 55159 48099 55165
rect 28721 55131 28779 55137
rect 28721 55097 28733 55131
rect 28767 55097 28779 55131
rect 28721 55091 28779 55097
rect 29196 55060 29224 55156
rect 29454 55060 29460 55072
rect 27028 55032 29460 55060
rect 27028 55020 27034 55032
rect 29454 55020 29460 55032
rect 29512 55020 29518 55072
rect 46474 55060 46480 55072
rect 46435 55032 46480 55060
rect 46474 55020 46480 55032
rect 46532 55020 46538 55072
rect 51258 55060 51264 55072
rect 51219 55032 51264 55060
rect 51258 55020 51264 55032
rect 51316 55020 51322 55072
rect 54588 55060 54616 55227
rect 56134 55224 56140 55236
rect 56192 55224 56198 55276
rect 55490 55060 55496 55072
rect 54588 55032 55496 55060
rect 55490 55020 55496 55032
rect 55548 55060 55554 55072
rect 57054 55060 57060 55072
rect 55548 55032 57060 55060
rect 55548 55020 55554 55032
rect 57054 55020 57060 55032
rect 57112 55020 57118 55072
rect 1104 54970 59340 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 59340 54970
rect 1104 54896 59340 54918
rect 23106 54856 23112 54868
rect 23067 54828 23112 54856
rect 23106 54816 23112 54828
rect 23164 54816 23170 54868
rect 25406 54816 25412 54868
rect 25464 54856 25470 54868
rect 25777 54859 25835 54865
rect 25777 54856 25789 54859
rect 25464 54828 25789 54856
rect 25464 54816 25470 54828
rect 25777 54825 25789 54828
rect 25823 54825 25835 54859
rect 25777 54819 25835 54825
rect 28166 54816 28172 54868
rect 28224 54856 28230 54868
rect 28261 54859 28319 54865
rect 28261 54856 28273 54859
rect 28224 54828 28273 54856
rect 28224 54816 28230 54828
rect 28261 54825 28273 54828
rect 28307 54825 28319 54859
rect 36630 54856 36636 54868
rect 36591 54828 36636 54856
rect 28261 54819 28319 54825
rect 36630 54816 36636 54828
rect 36688 54816 36694 54868
rect 41322 54816 41328 54868
rect 41380 54856 41386 54868
rect 41417 54859 41475 54865
rect 41417 54856 41429 54859
rect 41380 54828 41429 54856
rect 41380 54816 41386 54828
rect 41417 54825 41429 54828
rect 41463 54825 41475 54859
rect 49050 54856 49056 54868
rect 49011 54828 49056 54856
rect 41417 54819 41475 54825
rect 49050 54816 49056 54828
rect 49108 54816 49114 54868
rect 51166 54816 51172 54868
rect 51224 54856 51230 54868
rect 51537 54859 51595 54865
rect 51537 54856 51549 54859
rect 51224 54828 51549 54856
rect 51224 54816 51230 54828
rect 51537 54825 51549 54828
rect 51583 54825 51595 54859
rect 51537 54819 51595 54825
rect 6914 54680 6920 54732
rect 6972 54720 6978 54732
rect 14090 54720 14096 54732
rect 6972 54692 7017 54720
rect 14051 54692 14096 54720
rect 6972 54680 6978 54692
rect 14090 54680 14096 54692
rect 14148 54680 14154 54732
rect 21726 54720 21732 54732
rect 21687 54692 21732 54720
rect 21726 54680 21732 54692
rect 21784 54680 21790 54732
rect 57054 54720 57060 54732
rect 57015 54692 57060 54720
rect 57054 54680 57060 54692
rect 57112 54680 57118 54732
rect 3878 54612 3884 54664
rect 3936 54652 3942 54664
rect 5077 54655 5135 54661
rect 5077 54652 5089 54655
rect 3936 54624 5089 54652
rect 3936 54612 3942 54624
rect 5077 54621 5089 54624
rect 5123 54652 5135 54655
rect 5626 54652 5632 54664
rect 5123 54624 5632 54652
rect 5123 54621 5135 54624
rect 5077 54615 5135 54621
rect 5626 54612 5632 54624
rect 5684 54652 5690 54664
rect 6270 54652 6276 54664
rect 5684 54624 6276 54652
rect 5684 54612 5690 54624
rect 6270 54612 6276 54624
rect 6328 54612 6334 54664
rect 9490 54652 9496 54664
rect 9451 54624 9496 54652
rect 9490 54612 9496 54624
rect 9548 54612 9554 54664
rect 9760 54655 9818 54661
rect 9760 54621 9772 54655
rect 9806 54652 9818 54655
rect 10686 54652 10692 54664
rect 9806 54624 10692 54652
rect 9806 54621 9818 54624
rect 9760 54615 9818 54621
rect 10686 54612 10692 54624
rect 10744 54612 10750 54664
rect 14366 54661 14372 54664
rect 14360 54652 14372 54661
rect 14327 54624 14372 54652
rect 14360 54615 14372 54624
rect 14366 54612 14372 54615
rect 14424 54612 14430 54664
rect 15933 54655 15991 54661
rect 15933 54621 15945 54655
rect 15979 54652 15991 54655
rect 16574 54652 16580 54664
rect 15979 54624 16580 54652
rect 15979 54621 15991 54624
rect 15933 54615 15991 54621
rect 16574 54612 16580 54624
rect 16632 54612 16638 54664
rect 19889 54655 19947 54661
rect 19889 54621 19901 54655
rect 19935 54652 19947 54655
rect 20714 54652 20720 54664
rect 19935 54624 20720 54652
rect 19935 54621 19947 54624
rect 19889 54615 19947 54621
rect 20714 54612 20720 54624
rect 20772 54612 20778 54664
rect 23658 54612 23664 54664
rect 23716 54652 23722 54664
rect 24394 54652 24400 54664
rect 23716 54624 24400 54652
rect 23716 54612 23722 54624
rect 24394 54612 24400 54624
rect 24452 54612 24458 54664
rect 24664 54655 24722 54661
rect 24664 54621 24676 54655
rect 24710 54652 24722 54655
rect 25590 54652 25596 54664
rect 24710 54624 25596 54652
rect 24710 54621 24722 54624
rect 24664 54615 24722 54621
rect 25590 54612 25596 54624
rect 25648 54612 25654 54664
rect 26881 54655 26939 54661
rect 26881 54621 26893 54655
rect 26927 54652 26939 54655
rect 26970 54652 26976 54664
rect 26927 54624 26976 54652
rect 26927 54621 26939 54624
rect 26881 54615 26939 54621
rect 26970 54612 26976 54624
rect 27028 54612 27034 54664
rect 29454 54612 29460 54664
rect 29512 54652 29518 54664
rect 29549 54655 29607 54661
rect 29549 54652 29561 54655
rect 29512 54624 29561 54652
rect 29512 54612 29518 54624
rect 29549 54621 29561 54624
rect 29595 54621 29607 54655
rect 29549 54615 29607 54621
rect 35253 54655 35311 54661
rect 35253 54621 35265 54655
rect 35299 54652 35311 54655
rect 37093 54655 37151 54661
rect 37093 54652 37105 54655
rect 35299 54624 37105 54652
rect 35299 54621 35311 54624
rect 35253 54615 35311 54621
rect 37093 54621 37105 54624
rect 37139 54652 37151 54655
rect 37642 54652 37648 54664
rect 37139 54624 37648 54652
rect 37139 54621 37151 54624
rect 37093 54615 37151 54621
rect 37642 54612 37648 54624
rect 37700 54612 37706 54664
rect 40037 54655 40095 54661
rect 40037 54621 40049 54655
rect 40083 54652 40095 54655
rect 40586 54652 40592 54664
rect 40083 54624 40592 54652
rect 40083 54621 40095 54624
rect 40037 54615 40095 54621
rect 40586 54612 40592 54624
rect 40644 54612 40650 54664
rect 42981 54655 43039 54661
rect 42981 54621 42993 54655
rect 43027 54652 43039 54655
rect 45278 54652 45284 54664
rect 43027 54624 45284 54652
rect 43027 54621 43039 54624
rect 42981 54615 43039 54621
rect 45278 54612 45284 54624
rect 45336 54652 45342 54664
rect 45833 54655 45891 54661
rect 45833 54652 45845 54655
rect 45336 54624 45845 54652
rect 45336 54612 45342 54624
rect 45833 54621 45845 54624
rect 45879 54621 45891 54655
rect 45833 54615 45891 54621
rect 46100 54655 46158 54661
rect 46100 54621 46112 54655
rect 46146 54652 46158 54655
rect 46474 54652 46480 54664
rect 46146 54624 46480 54652
rect 46146 54621 46158 54624
rect 46100 54615 46158 54621
rect 46474 54612 46480 54624
rect 46532 54612 46538 54664
rect 47578 54612 47584 54664
rect 47636 54652 47642 54664
rect 47673 54655 47731 54661
rect 47673 54652 47685 54655
rect 47636 54624 47685 54652
rect 47636 54612 47642 54624
rect 47673 54621 47685 54624
rect 47719 54621 47731 54655
rect 50154 54652 50160 54664
rect 50115 54624 50160 54652
rect 47673 54615 47731 54621
rect 50154 54612 50160 54624
rect 50212 54612 50218 54664
rect 50424 54655 50482 54661
rect 50424 54621 50436 54655
rect 50470 54652 50482 54655
rect 51258 54652 51264 54664
rect 50470 54624 51264 54652
rect 50470 54621 50482 54624
rect 50424 54615 50482 54621
rect 51258 54612 51264 54624
rect 51316 54612 51322 54664
rect 51997 54655 52055 54661
rect 51997 54621 52009 54655
rect 52043 54621 52055 54655
rect 51997 54615 52055 54621
rect 52264 54655 52322 54661
rect 52264 54621 52276 54655
rect 52310 54652 52322 54655
rect 52546 54652 52552 54664
rect 52310 54624 52552 54652
rect 52310 54621 52322 54624
rect 52264 54615 52322 54621
rect 5344 54587 5402 54593
rect 5344 54553 5356 54587
rect 5390 54584 5402 54587
rect 5810 54584 5816 54596
rect 5390 54556 5816 54584
rect 5390 54553 5402 54556
rect 5344 54547 5402 54553
rect 5810 54544 5816 54556
rect 5868 54544 5874 54596
rect 7184 54587 7242 54593
rect 7184 54553 7196 54587
rect 7230 54584 7242 54587
rect 7742 54584 7748 54596
rect 7230 54556 7748 54584
rect 7230 54553 7242 54556
rect 7184 54547 7242 54553
rect 7742 54544 7748 54556
rect 7800 54544 7806 54596
rect 16206 54593 16212 54596
rect 16200 54547 16212 54593
rect 16264 54584 16270 54596
rect 20156 54587 20214 54593
rect 16264 54556 16300 54584
rect 16206 54544 16212 54547
rect 16264 54544 16270 54556
rect 20156 54553 20168 54587
rect 20202 54584 20214 54587
rect 21082 54584 21088 54596
rect 20202 54556 21088 54584
rect 20202 54553 20214 54556
rect 20156 54547 20214 54553
rect 21082 54544 21088 54556
rect 21140 54544 21146 54596
rect 21996 54587 22054 54593
rect 21996 54553 22008 54587
rect 22042 54584 22054 54587
rect 23198 54584 23204 54596
rect 22042 54556 23204 54584
rect 22042 54553 22054 54556
rect 21996 54547 22054 54553
rect 23198 54544 23204 54556
rect 23256 54544 23262 54596
rect 27148 54587 27206 54593
rect 27148 54553 27160 54587
rect 27194 54584 27206 54587
rect 28350 54584 28356 54596
rect 27194 54556 28356 54584
rect 27194 54553 27206 54556
rect 27148 54547 27206 54553
rect 28350 54544 28356 54556
rect 28408 54544 28414 54596
rect 29270 54544 29276 54596
rect 29328 54584 29334 54596
rect 29794 54587 29852 54593
rect 29794 54584 29806 54587
rect 29328 54556 29806 54584
rect 29328 54544 29334 54556
rect 29794 54553 29806 54556
rect 29840 54553 29852 54587
rect 29794 54547 29852 54553
rect 32401 54587 32459 54593
rect 32401 54553 32413 54587
rect 32447 54584 32459 54587
rect 32490 54584 32496 54596
rect 32447 54556 32496 54584
rect 32447 54553 32459 54556
rect 32401 54547 32459 54553
rect 32490 54544 32496 54556
rect 32548 54544 32554 54596
rect 33962 54584 33968 54596
rect 33923 54556 33968 54584
rect 33962 54544 33968 54556
rect 34020 54544 34026 54596
rect 35520 54587 35578 54593
rect 35520 54553 35532 54587
rect 35566 54584 35578 54587
rect 37360 54587 37418 54593
rect 35566 54556 35894 54584
rect 35566 54553 35578 54556
rect 35520 54547 35578 54553
rect 6454 54516 6460 54528
rect 6415 54488 6460 54516
rect 6454 54476 6460 54488
rect 6512 54476 6518 54528
rect 7558 54476 7564 54528
rect 7616 54516 7622 54528
rect 8297 54519 8355 54525
rect 8297 54516 8309 54519
rect 7616 54488 8309 54516
rect 7616 54476 7622 54488
rect 8297 54485 8309 54488
rect 8343 54485 8355 54519
rect 10870 54516 10876 54528
rect 10831 54488 10876 54516
rect 8297 54479 8355 54485
rect 10870 54476 10876 54488
rect 10928 54476 10934 54528
rect 15470 54516 15476 54528
rect 15431 54488 15476 54516
rect 15470 54476 15476 54488
rect 15528 54476 15534 54528
rect 16666 54476 16672 54528
rect 16724 54516 16730 54528
rect 17313 54519 17371 54525
rect 17313 54516 17325 54519
rect 16724 54488 17325 54516
rect 16724 54476 16730 54488
rect 17313 54485 17325 54488
rect 17359 54485 17371 54519
rect 21266 54516 21272 54528
rect 21227 54488 21272 54516
rect 17313 54479 17371 54485
rect 21266 54476 21272 54488
rect 21324 54476 21330 54528
rect 30926 54516 30932 54528
rect 30887 54488 30932 54516
rect 30926 54476 30932 54488
rect 30984 54476 30990 54528
rect 35866 54516 35894 54556
rect 37360 54553 37372 54587
rect 37406 54584 37418 54587
rect 39298 54584 39304 54596
rect 37406 54556 39304 54584
rect 37406 54553 37418 54556
rect 37360 54547 37418 54553
rect 39298 54544 39304 54556
rect 39356 54544 39362 54596
rect 40304 54587 40362 54593
rect 40304 54553 40316 54587
rect 40350 54584 40362 54587
rect 41782 54584 41788 54596
rect 40350 54556 41788 54584
rect 40350 54553 40362 54556
rect 40304 54547 40362 54553
rect 41782 54544 41788 54556
rect 41840 54544 41846 54596
rect 43248 54587 43306 54593
rect 43248 54553 43260 54587
rect 43294 54584 43306 54587
rect 44542 54584 44548 54596
rect 43294 54556 44548 54584
rect 43294 54553 43306 54556
rect 43248 54547 43306 54553
rect 44542 54544 44548 54556
rect 44600 54544 44606 54596
rect 47940 54587 47998 54593
rect 47940 54553 47952 54587
rect 47986 54584 47998 54587
rect 48958 54584 48964 54596
rect 47986 54556 48964 54584
rect 47986 54553 47998 54556
rect 47940 54547 47998 54553
rect 48958 54544 48964 54556
rect 49016 54544 49022 54596
rect 52012 54584 52040 54615
rect 52546 54612 52552 54624
rect 52604 54612 52610 54664
rect 52730 54584 52736 54596
rect 52012 54556 52736 54584
rect 52730 54544 52736 54556
rect 52788 54544 52794 54596
rect 57330 54593 57336 54596
rect 57324 54547 57336 54593
rect 57388 54584 57394 54596
rect 57388 54556 57424 54584
rect 57330 54544 57336 54547
rect 57388 54544 57394 54556
rect 38473 54519 38531 54525
rect 38473 54516 38485 54519
rect 35866 54488 38485 54516
rect 38473 54485 38485 54488
rect 38519 54485 38531 54519
rect 38473 54479 38531 54485
rect 44174 54476 44180 54528
rect 44232 54516 44238 54528
rect 44361 54519 44419 54525
rect 44361 54516 44373 54519
rect 44232 54488 44373 54516
rect 44232 54476 44238 54488
rect 44361 54485 44373 54488
rect 44407 54485 44419 54519
rect 47210 54516 47216 54528
rect 47171 54488 47216 54516
rect 44361 54479 44419 54485
rect 47210 54476 47216 54488
rect 47268 54476 47274 54528
rect 52546 54476 52552 54528
rect 52604 54516 52610 54528
rect 53377 54519 53435 54525
rect 53377 54516 53389 54519
rect 52604 54488 53389 54516
rect 52604 54476 52610 54488
rect 53377 54485 53389 54488
rect 53423 54485 53435 54519
rect 53377 54479 53435 54485
rect 58437 54519 58495 54525
rect 58437 54485 58449 54519
rect 58483 54516 58495 54519
rect 59449 54519 59507 54525
rect 59449 54516 59461 54519
rect 58483 54488 59461 54516
rect 58483 54485 58495 54488
rect 58437 54479 58495 54485
rect 59449 54485 59461 54488
rect 59495 54485 59507 54519
rect 59449 54479 59507 54485
rect 1104 54426 59340 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 59340 54426
rect 1104 54352 59340 54374
rect 7742 54312 7748 54324
rect 7703 54284 7748 54312
rect 7742 54272 7748 54284
rect 7800 54272 7806 54324
rect 23198 54312 23204 54324
rect 23159 54284 23204 54312
rect 23198 54272 23204 54284
rect 23256 54272 23262 54324
rect 25038 54312 25044 54324
rect 24999 54284 25044 54312
rect 25038 54272 25044 54284
rect 25096 54272 25102 54324
rect 28350 54312 28356 54324
rect 28311 54284 28356 54312
rect 28350 54272 28356 54284
rect 28408 54272 28414 54324
rect 30190 54312 30196 54324
rect 30151 54284 30196 54312
rect 30190 54272 30196 54284
rect 30248 54272 30254 54324
rect 33410 54272 33416 54324
rect 33468 54312 33474 54324
rect 33505 54315 33563 54321
rect 33505 54312 33517 54315
rect 33468 54284 33517 54312
rect 33468 54272 33474 54284
rect 33505 54281 33517 54284
rect 33551 54281 33563 54315
rect 48958 54312 48964 54324
rect 48919 54284 48964 54312
rect 33505 54275 33563 54281
rect 48958 54272 48964 54284
rect 49016 54272 49022 54324
rect 49694 54272 49700 54324
rect 49752 54312 49758 54324
rect 50890 54312 50896 54324
rect 49752 54284 49832 54312
rect 50851 54284 50896 54312
rect 49752 54272 49758 54284
rect 6454 54204 6460 54256
rect 6512 54244 6518 54256
rect 6610 54247 6668 54253
rect 6610 54244 6622 54247
rect 6512 54216 6622 54244
rect 6512 54204 6518 54216
rect 6610 54213 6622 54216
rect 6656 54213 6668 54247
rect 6610 54207 6668 54213
rect 9852 54247 9910 54253
rect 9852 54213 9864 54247
rect 9898 54244 9910 54247
rect 10870 54244 10876 54256
rect 9898 54216 10876 54244
rect 9898 54213 9910 54216
rect 9852 54207 9910 54213
rect 10870 54204 10876 54216
rect 10928 54204 10934 54256
rect 14912 54247 14970 54253
rect 14912 54213 14924 54247
rect 14958 54244 14970 54247
rect 15470 54244 15476 54256
rect 14958 54216 15476 54244
rect 14958 54213 14970 54216
rect 14912 54207 14970 54213
rect 15470 54204 15476 54216
rect 15528 54204 15534 54256
rect 16574 54204 16580 54256
rect 16632 54244 16638 54256
rect 17862 54244 17868 54256
rect 16632 54216 17868 54244
rect 16632 54204 16638 54216
rect 3136 54179 3194 54185
rect 3136 54145 3148 54179
rect 3182 54176 3194 54179
rect 5350 54176 5356 54188
rect 3182 54148 5356 54176
rect 3182 54145 3194 54148
rect 3136 54139 3194 54145
rect 5350 54136 5356 54148
rect 5408 54136 5414 54188
rect 6270 54136 6276 54188
rect 6328 54176 6334 54188
rect 6365 54179 6423 54185
rect 6365 54176 6377 54179
rect 6328 54148 6377 54176
rect 6328 54136 6334 54148
rect 6365 54145 6377 54148
rect 6411 54145 6423 54179
rect 6365 54139 6423 54145
rect 9306 54136 9312 54188
rect 9364 54176 9370 54188
rect 9585 54179 9643 54185
rect 9585 54176 9597 54179
rect 9364 54148 9597 54176
rect 9364 54136 9370 54148
rect 9585 54145 9597 54148
rect 9631 54145 9643 54179
rect 9585 54139 9643 54145
rect 11238 54136 11244 54188
rect 11296 54176 11302 54188
rect 16684 54185 16712 54216
rect 17862 54204 17868 54216
rect 17920 54204 17926 54256
rect 18693 54247 18751 54253
rect 18693 54213 18705 54247
rect 18739 54244 18751 54247
rect 20070 54244 20076 54256
rect 18739 54216 20076 54244
rect 18739 54213 18751 54216
rect 18693 54207 18751 54213
rect 20070 54204 20076 54216
rect 20128 54244 20134 54256
rect 20438 54244 20444 54256
rect 20128 54216 20444 54244
rect 20128 54204 20134 54216
rect 20438 54204 20444 54216
rect 20496 54204 20502 54256
rect 21266 54204 21272 54256
rect 21324 54244 21330 54256
rect 23934 54253 23940 54256
rect 22066 54247 22124 54253
rect 22066 54244 22078 54247
rect 21324 54216 22078 54244
rect 21324 54204 21330 54216
rect 22066 54213 22078 54216
rect 22112 54213 22124 54247
rect 22066 54207 22124 54213
rect 23928 54207 23940 54253
rect 23992 54244 23998 54256
rect 29080 54247 29138 54253
rect 23992 54216 24028 54244
rect 23934 54204 23940 54207
rect 23992 54204 23998 54216
rect 29080 54213 29092 54247
rect 29126 54244 29138 54247
rect 30926 54244 30932 54256
rect 29126 54216 30932 54244
rect 29126 54213 29138 54216
rect 29080 54207 29138 54213
rect 30926 54204 30932 54216
rect 30984 54204 30990 54256
rect 33962 54244 33968 54256
rect 32324 54216 33968 54244
rect 11773 54179 11831 54185
rect 11773 54176 11785 54179
rect 11296 54148 11785 54176
rect 11296 54136 11302 54148
rect 11773 54145 11785 54148
rect 11819 54145 11831 54179
rect 11773 54139 11831 54145
rect 14645 54179 14703 54185
rect 14645 54145 14657 54179
rect 14691 54176 14703 54179
rect 16669 54179 16727 54185
rect 16669 54176 16681 54179
rect 14691 54148 16681 54176
rect 14691 54145 14703 54148
rect 14645 54139 14703 54145
rect 16669 54145 16681 54148
rect 16715 54145 16727 54179
rect 16669 54139 16727 54145
rect 16936 54179 16994 54185
rect 16936 54145 16948 54179
rect 16982 54176 16994 54179
rect 17770 54176 17776 54188
rect 16982 54148 17776 54176
rect 16982 54145 16994 54148
rect 16936 54139 16994 54145
rect 17770 54136 17776 54148
rect 17828 54136 17834 54188
rect 23658 54176 23664 54188
rect 23619 54148 23664 54176
rect 23658 54136 23664 54148
rect 23716 54136 23722 54188
rect 26970 54176 26976 54188
rect 26931 54148 26976 54176
rect 26970 54136 26976 54148
rect 27028 54136 27034 54188
rect 27246 54185 27252 54188
rect 27240 54139 27252 54185
rect 27304 54176 27310 54188
rect 28813 54179 28871 54185
rect 27304 54148 27340 54176
rect 27246 54136 27252 54139
rect 27304 54136 27310 54148
rect 28813 54145 28825 54179
rect 28859 54176 28871 54179
rect 29546 54176 29552 54188
rect 28859 54148 29552 54176
rect 28859 54145 28871 54148
rect 28813 54139 28871 54145
rect 29546 54136 29552 54148
rect 29604 54136 29610 54188
rect 32122 54176 32128 54188
rect 32035 54148 32128 54176
rect 32122 54136 32128 54148
rect 32180 54176 32186 54188
rect 32324 54176 32352 54216
rect 33962 54204 33968 54216
rect 34020 54204 34026 54256
rect 40494 54244 40500 54256
rect 38672 54216 40500 54244
rect 32180 54148 32352 54176
rect 32392 54179 32450 54185
rect 32180 54136 32186 54148
rect 32392 54145 32404 54179
rect 32438 54176 32450 54179
rect 32766 54176 32772 54188
rect 32438 54148 32772 54176
rect 32438 54145 32450 54148
rect 32392 54139 32450 54145
rect 32766 54136 32772 54148
rect 32824 54136 32830 54188
rect 33502 54136 33508 54188
rect 33560 54176 33566 54188
rect 38672 54185 38700 54216
rect 40494 54204 40500 54216
rect 40552 54204 40558 54256
rect 45278 54244 45284 54256
rect 43824 54216 45284 54244
rect 34221 54179 34279 54185
rect 34221 54176 34233 54179
rect 33560 54148 34233 54176
rect 33560 54136 33566 54148
rect 34221 54145 34233 54148
rect 34267 54145 34279 54179
rect 34221 54139 34279 54145
rect 38657 54179 38715 54185
rect 38657 54145 38669 54179
rect 38703 54145 38715 54179
rect 38657 54139 38715 54145
rect 38924 54179 38982 54185
rect 38924 54145 38936 54179
rect 38970 54176 38982 54179
rect 40034 54176 40040 54188
rect 38970 54148 40040 54176
rect 38970 54145 38982 54148
rect 38924 54139 38982 54145
rect 40034 54136 40040 54148
rect 40092 54136 40098 54188
rect 40764 54179 40822 54185
rect 40764 54145 40776 54179
rect 40810 54176 40822 54179
rect 42610 54176 42616 54188
rect 40810 54148 42616 54176
rect 40810 54145 40822 54148
rect 40764 54139 40822 54145
rect 42610 54136 42616 54148
rect 42668 54136 42674 54188
rect 43824 54185 43852 54216
rect 45278 54204 45284 54216
rect 45336 54204 45342 54256
rect 45916 54247 45974 54253
rect 45916 54213 45928 54247
rect 45962 54244 45974 54247
rect 47210 54244 47216 54256
rect 45962 54216 47216 54244
rect 45962 54213 45974 54216
rect 45916 54207 45974 54213
rect 47210 54204 47216 54216
rect 47268 54204 47274 54256
rect 49804 54253 49832 54284
rect 50890 54272 50896 54284
rect 50948 54272 50954 54324
rect 56134 54272 56140 54324
rect 56192 54312 56198 54324
rect 56873 54315 56931 54321
rect 56873 54312 56885 54315
rect 56192 54284 56885 54312
rect 56192 54272 56198 54284
rect 56873 54281 56885 54284
rect 56919 54281 56931 54315
rect 56873 54275 56931 54281
rect 49780 54247 49838 54253
rect 49780 54213 49792 54247
rect 49826 54213 49838 54247
rect 49780 54207 49838 54213
rect 43809 54179 43867 54185
rect 43809 54145 43821 54179
rect 43855 54145 43867 54179
rect 43809 54139 43867 54145
rect 44076 54179 44134 54185
rect 44076 54145 44088 54179
rect 44122 54176 44134 54179
rect 44818 54176 44824 54188
rect 44122 54148 44824 54176
rect 44122 54145 44134 54148
rect 44076 54139 44134 54145
rect 44818 54136 44824 54148
rect 44876 54136 44882 54188
rect 47848 54179 47906 54185
rect 47848 54145 47860 54179
rect 47894 54176 47906 54179
rect 48958 54176 48964 54188
rect 47894 54148 48964 54176
rect 47894 54145 47906 54148
rect 47848 54139 47906 54145
rect 48958 54136 48964 54148
rect 49016 54136 49022 54188
rect 49513 54179 49571 54185
rect 49513 54145 49525 54179
rect 49559 54176 49571 54179
rect 50154 54176 50160 54188
rect 49559 54148 50160 54176
rect 49559 54145 49571 54148
rect 49513 54139 49571 54145
rect 50154 54136 50160 54148
rect 50212 54136 50218 54188
rect 52454 54136 52460 54188
rect 52512 54176 52518 54188
rect 52989 54179 53047 54185
rect 52989 54176 53001 54179
rect 52512 54148 53001 54176
rect 52512 54136 52518 54148
rect 52989 54145 53001 54148
rect 53035 54145 53047 54179
rect 52989 54139 53047 54145
rect 55398 54136 55404 54188
rect 55456 54176 55462 54188
rect 55749 54179 55807 54185
rect 55749 54176 55761 54179
rect 55456 54148 55761 54176
rect 55456 54136 55462 54148
rect 55749 54145 55761 54148
rect 55795 54145 55807 54179
rect 55749 54139 55807 54145
rect 2866 54108 2872 54120
rect 2827 54080 2872 54108
rect 2866 54068 2872 54080
rect 2924 54068 2930 54120
rect 11517 54111 11575 54117
rect 11517 54077 11529 54111
rect 11563 54077 11575 54111
rect 11517 54071 11575 54077
rect 20441 54111 20499 54117
rect 20441 54077 20453 54111
rect 20487 54108 20499 54111
rect 20806 54108 20812 54120
rect 20487 54080 20812 54108
rect 20487 54077 20499 54080
rect 20441 54071 20499 54077
rect 4249 53975 4307 53981
rect 4249 53941 4261 53975
rect 4295 53972 4307 53975
rect 4614 53972 4620 53984
rect 4295 53944 4620 53972
rect 4295 53941 4307 53944
rect 4249 53935 4307 53941
rect 4614 53932 4620 53944
rect 4672 53932 4678 53984
rect 10962 53972 10968 53984
rect 10923 53944 10968 53972
rect 10962 53932 10968 53944
rect 11020 53932 11026 53984
rect 11532 53972 11560 54071
rect 20806 54068 20812 54080
rect 20864 54068 20870 54120
rect 21818 54108 21824 54120
rect 21779 54080 21824 54108
rect 21818 54068 21824 54080
rect 21876 54068 21882 54120
rect 33962 54108 33968 54120
rect 33923 54080 33968 54108
rect 33962 54068 33968 54080
rect 34020 54068 34026 54120
rect 40494 54108 40500 54120
rect 40455 54080 40500 54108
rect 40494 54068 40500 54080
rect 40552 54068 40558 54120
rect 45278 54068 45284 54120
rect 45336 54108 45342 54120
rect 45649 54111 45707 54117
rect 45649 54108 45661 54111
rect 45336 54080 45661 54108
rect 45336 54068 45342 54080
rect 45649 54077 45661 54080
rect 45695 54077 45707 54111
rect 47578 54108 47584 54120
rect 47539 54080 47584 54108
rect 45649 54071 45707 54077
rect 47578 54068 47584 54080
rect 47636 54068 47642 54120
rect 52730 54108 52736 54120
rect 52643 54080 52736 54108
rect 52730 54068 52736 54080
rect 52788 54068 52794 54120
rect 55490 54108 55496 54120
rect 55451 54080 55496 54108
rect 55490 54068 55496 54080
rect 55548 54068 55554 54120
rect 11698 53972 11704 53984
rect 11532 53944 11704 53972
rect 11698 53932 11704 53944
rect 11756 53932 11762 53984
rect 12894 53972 12900 53984
rect 12855 53944 12900 53972
rect 12894 53932 12900 53944
rect 12952 53932 12958 53984
rect 16022 53972 16028 53984
rect 15983 53944 16028 53972
rect 16022 53932 16028 53944
rect 16080 53932 16086 53984
rect 18046 53972 18052 53984
rect 18007 53944 18052 53972
rect 18046 53932 18052 53944
rect 18104 53932 18110 53984
rect 33226 53932 33232 53984
rect 33284 53972 33290 53984
rect 35345 53975 35403 53981
rect 35345 53972 35357 53975
rect 33284 53944 35357 53972
rect 33284 53932 33290 53944
rect 35345 53941 35357 53944
rect 35391 53941 35403 53975
rect 35345 53935 35403 53941
rect 38654 53932 38660 53984
rect 38712 53972 38718 53984
rect 40037 53975 40095 53981
rect 40037 53972 40049 53975
rect 38712 53944 40049 53972
rect 38712 53932 38718 53944
rect 40037 53941 40049 53944
rect 40083 53941 40095 53975
rect 40037 53935 40095 53941
rect 41414 53932 41420 53984
rect 41472 53972 41478 53984
rect 41877 53975 41935 53981
rect 41877 53972 41889 53975
rect 41472 53944 41889 53972
rect 41472 53932 41478 53944
rect 41877 53941 41889 53944
rect 41923 53941 41935 53975
rect 45186 53972 45192 53984
rect 45147 53944 45192 53972
rect 41877 53935 41935 53941
rect 45186 53932 45192 53944
rect 45244 53932 45250 53984
rect 47026 53972 47032 53984
rect 46987 53944 47032 53972
rect 47026 53932 47032 53944
rect 47084 53932 47090 53984
rect 52748 53972 52776 54068
rect 52914 53972 52920 53984
rect 52748 53944 52920 53972
rect 52914 53932 52920 53944
rect 52972 53932 52978 53984
rect 54110 53972 54116 53984
rect 54071 53944 54116 53972
rect 54110 53932 54116 53944
rect 54168 53932 54174 53984
rect 1104 53882 59340 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 59340 53882
rect 1104 53808 59340 53830
rect 11238 53768 11244 53780
rect 11199 53740 11244 53768
rect 11238 53728 11244 53740
rect 11296 53728 11302 53780
rect 15933 53771 15991 53777
rect 15933 53737 15945 53771
rect 15979 53768 15991 53771
rect 16206 53768 16212 53780
rect 15979 53740 16212 53768
rect 15979 53737 15991 53740
rect 15933 53731 15991 53737
rect 16206 53728 16212 53740
rect 16264 53728 16270 53780
rect 17770 53768 17776 53780
rect 17731 53740 17776 53768
rect 17770 53728 17776 53740
rect 17828 53728 17834 53780
rect 21082 53728 21088 53780
rect 21140 53768 21146 53780
rect 22465 53771 22523 53777
rect 22465 53768 22477 53771
rect 21140 53740 22477 53768
rect 21140 53728 21146 53740
rect 22465 53737 22477 53740
rect 22511 53737 22523 53771
rect 22465 53731 22523 53737
rect 27246 53728 27252 53780
rect 27304 53768 27310 53780
rect 27341 53771 27399 53777
rect 27341 53768 27353 53771
rect 27304 53740 27353 53768
rect 27304 53728 27310 53740
rect 27341 53737 27353 53740
rect 27387 53737 27399 53771
rect 32766 53768 32772 53780
rect 32727 53740 32772 53768
rect 27341 53731 27399 53737
rect 32766 53728 32772 53740
rect 32824 53728 32830 53780
rect 39298 53768 39304 53780
rect 39259 53740 39304 53768
rect 39298 53728 39304 53740
rect 39356 53728 39362 53780
rect 42610 53768 42616 53780
rect 42571 53740 42616 53768
rect 42610 53728 42616 53740
rect 42668 53728 42674 53780
rect 52454 53768 52460 53780
rect 52415 53740 52460 53768
rect 52454 53728 52460 53740
rect 52512 53728 52518 53780
rect 2866 53592 2872 53644
rect 2924 53632 2930 53644
rect 3786 53632 3792 53644
rect 2924 53604 3792 53632
rect 2924 53592 2930 53604
rect 3786 53592 3792 53604
rect 3844 53592 3850 53644
rect 5626 53632 5632 53644
rect 5587 53604 5632 53632
rect 5626 53592 5632 53604
rect 5684 53592 5690 53644
rect 14553 53635 14611 53641
rect 14553 53601 14565 53635
rect 14599 53632 14611 53635
rect 43070 53632 43076 53644
rect 14599 53604 14688 53632
rect 43031 53604 43076 53632
rect 14599 53601 14611 53604
rect 14553 53595 14611 53601
rect 4056 53567 4114 53573
rect 4056 53533 4068 53567
rect 4102 53564 4114 53567
rect 4614 53564 4620 53576
rect 4102 53536 4620 53564
rect 4102 53533 4114 53536
rect 4056 53527 4114 53533
rect 4614 53524 4620 53536
rect 4672 53524 4678 53576
rect 9490 53524 9496 53576
rect 9548 53564 9554 53576
rect 9861 53567 9919 53573
rect 9861 53564 9873 53567
rect 9548 53536 9873 53564
rect 9548 53524 9554 53536
rect 9861 53533 9873 53536
rect 9907 53533 9919 53567
rect 9861 53527 9919 53533
rect 10128 53567 10186 53573
rect 10128 53533 10140 53567
rect 10174 53564 10186 53567
rect 10962 53564 10968 53576
rect 10174 53536 10968 53564
rect 10174 53533 10186 53536
rect 10128 53527 10186 53533
rect 5874 53499 5932 53505
rect 5874 53496 5886 53499
rect 5184 53468 5886 53496
rect 5184 53437 5212 53468
rect 5874 53465 5886 53468
rect 5920 53465 5932 53499
rect 9876 53496 9904 53527
rect 10962 53524 10968 53536
rect 11020 53524 11026 53576
rect 11698 53564 11704 53576
rect 11659 53536 11704 53564
rect 11698 53524 11704 53536
rect 11756 53524 11762 53576
rect 11968 53567 12026 53573
rect 11968 53533 11980 53567
rect 12014 53564 12026 53567
rect 12894 53564 12900 53576
rect 12014 53536 12900 53564
rect 12014 53533 12026 53536
rect 11968 53527 12026 53533
rect 12894 53524 12900 53536
rect 12952 53524 12958 53576
rect 11716 53496 11744 53524
rect 14660 53508 14688 53604
rect 43070 53592 43076 53604
rect 43128 53592 43134 53644
rect 50154 53592 50160 53644
rect 50212 53632 50218 53644
rect 51077 53635 51135 53641
rect 51077 53632 51089 53635
rect 50212 53604 51089 53632
rect 50212 53592 50218 53604
rect 51077 53601 51089 53604
rect 51123 53601 51135 53635
rect 51077 53595 51135 53601
rect 14820 53567 14878 53573
rect 14820 53533 14832 53567
rect 14866 53564 14878 53567
rect 16022 53564 16028 53576
rect 14866 53536 16028 53564
rect 14866 53533 14878 53536
rect 14820 53527 14878 53533
rect 16022 53524 16028 53536
rect 16080 53524 16086 53576
rect 16666 53573 16672 53576
rect 16393 53567 16451 53573
rect 16393 53533 16405 53567
rect 16439 53533 16451 53567
rect 16660 53564 16672 53573
rect 16627 53536 16672 53564
rect 16393 53527 16451 53533
rect 16660 53527 16672 53536
rect 9876 53468 11744 53496
rect 5874 53459 5932 53465
rect 14642 53456 14648 53508
rect 14700 53496 14706 53508
rect 16408 53496 16436 53527
rect 16666 53524 16672 53527
rect 16724 53524 16730 53576
rect 17862 53524 17868 53576
rect 17920 53564 17926 53576
rect 18506 53564 18512 53576
rect 17920 53536 18512 53564
rect 17920 53524 17926 53536
rect 18506 53524 18512 53536
rect 18564 53564 18570 53576
rect 19245 53567 19303 53573
rect 19245 53564 19257 53567
rect 18564 53536 19257 53564
rect 18564 53524 18570 53536
rect 19245 53533 19257 53536
rect 19291 53564 19303 53567
rect 20806 53564 20812 53576
rect 19291 53536 20812 53564
rect 19291 53533 19303 53536
rect 19245 53527 19303 53533
rect 20806 53524 20812 53536
rect 20864 53524 20870 53576
rect 21085 53567 21143 53573
rect 21085 53533 21097 53567
rect 21131 53564 21143 53567
rect 21818 53564 21824 53576
rect 21131 53536 21824 53564
rect 21131 53533 21143 53536
rect 21085 53527 21143 53533
rect 21818 53524 21824 53536
rect 21876 53524 21882 53576
rect 25038 53524 25044 53576
rect 25096 53564 25102 53576
rect 25961 53567 26019 53573
rect 25961 53564 25973 53567
rect 25096 53536 25973 53564
rect 25096 53524 25102 53536
rect 25961 53533 25973 53536
rect 26007 53564 26019 53567
rect 26970 53564 26976 53576
rect 26007 53536 26976 53564
rect 26007 53533 26019 53536
rect 25961 53527 26019 53533
rect 26970 53524 26976 53536
rect 27028 53524 27034 53576
rect 29546 53564 29552 53576
rect 29459 53536 29552 53564
rect 29546 53524 29552 53536
rect 29604 53524 29610 53576
rect 29822 53573 29828 53576
rect 29816 53527 29828 53573
rect 29880 53564 29886 53576
rect 31389 53567 31447 53573
rect 31389 53564 31401 53567
rect 29880 53536 29916 53564
rect 30024 53536 31401 53564
rect 29822 53524 29828 53527
rect 29880 53524 29886 53536
rect 14700 53468 16436 53496
rect 19512 53499 19570 53505
rect 14700 53456 14706 53468
rect 19512 53465 19524 53499
rect 19558 53496 19570 53499
rect 19978 53496 19984 53508
rect 19558 53468 19984 53496
rect 19558 53465 19570 53468
rect 19512 53459 19570 53465
rect 19978 53456 19984 53468
rect 20036 53456 20042 53508
rect 20714 53456 20720 53508
rect 20772 53496 20778 53508
rect 21330 53499 21388 53505
rect 21330 53496 21342 53499
rect 20772 53468 21342 53496
rect 20772 53456 20778 53468
rect 21330 53465 21342 53468
rect 21376 53465 21388 53499
rect 21330 53459 21388 53465
rect 26228 53499 26286 53505
rect 26228 53465 26240 53499
rect 26274 53496 26286 53499
rect 26418 53496 26424 53508
rect 26274 53468 26424 53496
rect 26274 53465 26286 53468
rect 26228 53459 26286 53465
rect 26418 53456 26424 53468
rect 26476 53456 26482 53508
rect 29564 53496 29592 53524
rect 30024 53496 30052 53536
rect 31389 53533 31401 53536
rect 31435 53564 31447 53567
rect 32122 53564 32128 53576
rect 31435 53536 32128 53564
rect 31435 53533 31447 53536
rect 31389 53527 31447 53533
rect 32122 53524 32128 53536
rect 32180 53524 32186 53576
rect 34698 53564 34704 53576
rect 34659 53536 34704 53564
rect 34698 53524 34704 53536
rect 34756 53524 34762 53576
rect 37918 53564 37924 53576
rect 37879 53536 37924 53564
rect 37918 53524 37924 53536
rect 37976 53524 37982 53576
rect 38188 53567 38246 53573
rect 38188 53533 38200 53567
rect 38234 53564 38246 53567
rect 38654 53564 38660 53576
rect 38234 53536 38660 53564
rect 38234 53533 38246 53536
rect 38188 53527 38246 53533
rect 38654 53524 38660 53536
rect 38712 53524 38718 53576
rect 40494 53524 40500 53576
rect 40552 53564 40558 53576
rect 41233 53567 41291 53573
rect 41233 53564 41245 53567
rect 40552 53536 41245 53564
rect 40552 53524 40558 53536
rect 41233 53533 41245 53536
rect 41279 53564 41291 53567
rect 43088 53564 43116 53592
rect 45278 53564 45284 53576
rect 41279 53536 43116 53564
rect 45239 53536 45284 53564
rect 41279 53533 41291 53536
rect 41233 53527 41291 53533
rect 45278 53524 45284 53536
rect 45336 53524 45342 53576
rect 45548 53567 45606 53573
rect 45548 53533 45560 53567
rect 45594 53564 45606 53567
rect 47026 53564 47032 53576
rect 45594 53536 47032 53564
rect 45594 53533 45606 53536
rect 45548 53527 45606 53533
rect 47026 53524 47032 53536
rect 47084 53524 47090 53576
rect 47118 53524 47124 53576
rect 47176 53564 47182 53576
rect 51344 53567 51402 53573
rect 47176 53536 47221 53564
rect 47176 53524 47182 53536
rect 51344 53533 51356 53567
rect 51390 53564 51402 53567
rect 52546 53564 52552 53576
rect 51390 53536 52552 53564
rect 51390 53533 51402 53536
rect 51344 53527 51402 53533
rect 52546 53524 52552 53536
rect 52604 53524 52610 53576
rect 52914 53564 52920 53576
rect 52875 53536 52920 53564
rect 52914 53524 52920 53536
rect 52972 53524 52978 53576
rect 53184 53567 53242 53573
rect 53184 53533 53196 53567
rect 53230 53564 53242 53567
rect 54110 53564 54116 53576
rect 53230 53536 54116 53564
rect 53230 53533 53242 53536
rect 53184 53527 53242 53533
rect 54110 53524 54116 53536
rect 54168 53524 54174 53576
rect 55950 53524 55956 53576
rect 56008 53564 56014 53576
rect 56781 53567 56839 53573
rect 56781 53564 56793 53567
rect 56008 53536 56793 53564
rect 56008 53524 56014 53536
rect 56781 53533 56793 53536
rect 56827 53533 56839 53567
rect 56781 53527 56839 53533
rect 29564 53468 30052 53496
rect 30834 53456 30840 53508
rect 30892 53496 30898 53508
rect 31634 53499 31692 53505
rect 31634 53496 31646 53499
rect 30892 53468 31646 53496
rect 30892 53456 30898 53468
rect 31634 53465 31646 53468
rect 31680 53465 31692 53499
rect 31634 53459 31692 53465
rect 34054 53456 34060 53508
rect 34112 53496 34118 53508
rect 34946 53499 35004 53505
rect 34946 53496 34958 53499
rect 34112 53468 34958 53496
rect 34112 53456 34118 53468
rect 34946 53465 34958 53468
rect 34992 53465 35004 53499
rect 34946 53459 35004 53465
rect 41500 53499 41558 53505
rect 41500 53465 41512 53499
rect 41546 53496 41558 53499
rect 41874 53496 41880 53508
rect 41546 53468 41880 53496
rect 41546 53465 41558 53468
rect 41500 53459 41558 53465
rect 41874 53456 41880 53468
rect 41932 53456 41938 53508
rect 43340 53499 43398 53505
rect 43340 53465 43352 53499
rect 43386 53496 43398 53499
rect 44358 53496 44364 53508
rect 43386 53468 44364 53496
rect 43386 53465 43398 53468
rect 43340 53459 43398 53465
rect 44358 53456 44364 53468
rect 44416 53456 44422 53508
rect 57048 53499 57106 53505
rect 57048 53465 57060 53499
rect 57094 53496 57106 53499
rect 57698 53496 57704 53508
rect 57094 53468 57704 53496
rect 57094 53465 57106 53468
rect 57048 53459 57106 53465
rect 57698 53456 57704 53468
rect 57756 53456 57762 53508
rect 5169 53431 5227 53437
rect 5169 53397 5181 53431
rect 5215 53397 5227 53431
rect 7006 53428 7012 53440
rect 6967 53400 7012 53428
rect 5169 53391 5227 53397
rect 7006 53388 7012 53400
rect 7064 53388 7070 53440
rect 13078 53428 13084 53440
rect 13039 53400 13084 53428
rect 13078 53388 13084 53400
rect 13136 53388 13142 53440
rect 20622 53428 20628 53440
rect 20583 53400 20628 53428
rect 20622 53388 20628 53400
rect 20680 53388 20686 53440
rect 30926 53428 30932 53440
rect 30887 53400 30932 53428
rect 30926 53388 30932 53400
rect 30984 53388 30990 53440
rect 36078 53428 36084 53440
rect 36039 53400 36084 53428
rect 36078 53388 36084 53400
rect 36136 53388 36142 53440
rect 44450 53428 44456 53440
rect 44411 53400 44456 53428
rect 44450 53388 44456 53400
rect 44508 53388 44514 53440
rect 46658 53428 46664 53440
rect 46619 53400 46664 53428
rect 46658 53388 46664 53400
rect 46716 53388 46722 53440
rect 47578 53388 47584 53440
rect 47636 53428 47642 53440
rect 48409 53431 48467 53437
rect 48409 53428 48421 53431
rect 47636 53400 48421 53428
rect 47636 53388 47642 53400
rect 48409 53397 48421 53400
rect 48455 53397 48467 53431
rect 48409 53391 48467 53397
rect 51350 53388 51356 53440
rect 51408 53428 51414 53440
rect 54297 53431 54355 53437
rect 54297 53428 54309 53431
rect 51408 53400 54309 53428
rect 51408 53388 51414 53400
rect 54297 53397 54309 53400
rect 54343 53397 54355 53431
rect 58158 53428 58164 53440
rect 58119 53400 58164 53428
rect 54297 53391 54355 53397
rect 58158 53388 58164 53400
rect 58216 53388 58222 53440
rect 1104 53338 59340 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 59340 53338
rect 1104 53264 59340 53286
rect 3513 53227 3571 53233
rect 3513 53193 3525 53227
rect 3559 53193 3571 53227
rect 5350 53224 5356 53236
rect 5311 53196 5356 53224
rect 3513 53187 3571 53193
rect 2866 53156 2872 53168
rect 2148 53128 2872 53156
rect 2148 53097 2176 53128
rect 2866 53116 2872 53128
rect 2924 53156 2930 53168
rect 3528 53156 3556 53187
rect 5350 53184 5356 53196
rect 5408 53184 5414 53236
rect 7926 53224 7932 53236
rect 7887 53196 7932 53224
rect 7926 53184 7932 53196
rect 7984 53184 7990 53236
rect 19889 53227 19947 53233
rect 19889 53193 19901 53227
rect 19935 53224 19947 53227
rect 19978 53224 19984 53236
rect 19935 53196 19984 53224
rect 19935 53193 19947 53196
rect 19889 53187 19947 53193
rect 19978 53184 19984 53196
rect 20036 53184 20042 53236
rect 26418 53224 26424 53236
rect 26379 53196 26424 53224
rect 26418 53184 26424 53196
rect 26476 53184 26482 53236
rect 30374 53224 30380 53236
rect 27816 53196 30380 53224
rect 4218 53159 4276 53165
rect 4218 53156 4230 53159
rect 2924 53128 3464 53156
rect 3528 53128 4230 53156
rect 2924 53116 2930 53128
rect 2133 53091 2191 53097
rect 2133 53057 2145 53091
rect 2179 53057 2191 53091
rect 2133 53051 2191 53057
rect 2400 53091 2458 53097
rect 2400 53057 2412 53091
rect 2446 53088 2458 53091
rect 3234 53088 3240 53100
rect 2446 53060 3240 53088
rect 2446 53057 2458 53060
rect 2400 53051 2458 53057
rect 3234 53048 3240 53060
rect 3292 53048 3298 53100
rect 3436 53088 3464 53128
rect 4218 53125 4230 53128
rect 4264 53125 4276 53159
rect 4218 53119 4276 53125
rect 6816 53159 6874 53165
rect 6816 53125 6828 53159
rect 6862 53156 6874 53159
rect 7558 53156 7564 53168
rect 6862 53128 7564 53156
rect 6862 53125 6874 53128
rect 6816 53119 6874 53125
rect 7558 53116 7564 53128
rect 7616 53116 7622 53168
rect 13081 53159 13139 53165
rect 13081 53125 13093 53159
rect 13127 53156 13139 53159
rect 13354 53156 13360 53168
rect 13127 53128 13360 53156
rect 13127 53125 13139 53128
rect 13081 53119 13139 53125
rect 13354 53116 13360 53128
rect 13412 53156 13418 53168
rect 13814 53156 13820 53168
rect 13412 53128 13820 53156
rect 13412 53116 13418 53128
rect 13814 53116 13820 53128
rect 13872 53116 13878 53168
rect 14642 53156 14648 53168
rect 14603 53128 14648 53156
rect 14642 53116 14648 53128
rect 14700 53116 14706 53168
rect 16936 53159 16994 53165
rect 16936 53125 16948 53159
rect 16982 53156 16994 53159
rect 18046 53156 18052 53168
rect 16982 53128 18052 53156
rect 16982 53125 16994 53128
rect 16936 53119 16994 53125
rect 18046 53116 18052 53128
rect 18104 53116 18110 53168
rect 23468 53159 23526 53165
rect 23468 53125 23480 53159
rect 23514 53156 23526 53159
rect 27816 53156 27844 53196
rect 30374 53184 30380 53196
rect 30432 53184 30438 53236
rect 30834 53224 30840 53236
rect 30795 53196 30840 53224
rect 30834 53184 30840 53196
rect 30892 53184 30898 53236
rect 33134 53184 33140 53236
rect 33192 53224 33198 53236
rect 33505 53227 33563 53233
rect 33505 53224 33517 53227
rect 33192 53196 33517 53224
rect 33192 53184 33198 53196
rect 33505 53193 33517 53196
rect 33551 53193 33563 53227
rect 40034 53224 40040 53236
rect 39995 53196 40040 53224
rect 33505 53187 33563 53193
rect 40034 53184 40040 53196
rect 40092 53184 40098 53236
rect 41874 53224 41880 53236
rect 41835 53196 41880 53224
rect 41874 53184 41880 53196
rect 41932 53184 41938 53236
rect 44818 53224 44824 53236
rect 44779 53196 44824 53224
rect 44818 53184 44824 53196
rect 44876 53184 44882 53236
rect 48958 53224 48964 53236
rect 48919 53196 48964 53224
rect 48958 53184 48964 53196
rect 49016 53184 49022 53236
rect 55033 53227 55091 53233
rect 55033 53193 55045 53227
rect 55079 53224 55091 53227
rect 55398 53224 55404 53236
rect 55079 53196 55404 53224
rect 55079 53193 55091 53196
rect 55033 53187 55091 53193
rect 55398 53184 55404 53196
rect 55456 53184 55462 53236
rect 57330 53224 57336 53236
rect 57291 53196 57336 53224
rect 57330 53184 57336 53196
rect 57388 53184 57394 53236
rect 23514 53128 27844 53156
rect 29724 53159 29782 53165
rect 23514 53125 23526 53128
rect 23468 53119 23526 53125
rect 29724 53125 29736 53159
rect 29770 53156 29782 53159
rect 30926 53156 30932 53168
rect 29770 53128 30932 53156
rect 29770 53125 29782 53128
rect 29724 53119 29782 53125
rect 30926 53116 30932 53128
rect 30984 53116 30990 53168
rect 32398 53165 32404 53168
rect 32392 53156 32404 53165
rect 32359 53128 32404 53156
rect 32392 53119 32404 53128
rect 32398 53116 32404 53119
rect 32456 53116 32462 53168
rect 34232 53159 34290 53165
rect 34232 53125 34244 53159
rect 34278 53156 34290 53159
rect 36078 53156 36084 53168
rect 34278 53128 36084 53156
rect 34278 53125 34290 53128
rect 34232 53119 34290 53125
rect 36078 53116 36084 53128
rect 36136 53116 36142 53168
rect 38930 53165 38936 53168
rect 38924 53156 38936 53165
rect 38891 53128 38936 53156
rect 38924 53119 38936 53128
rect 38930 53116 38936 53119
rect 38988 53116 38994 53168
rect 40764 53159 40822 53165
rect 40764 53125 40776 53159
rect 40810 53156 40822 53159
rect 44174 53156 44180 53168
rect 40810 53128 44180 53156
rect 40810 53125 40822 53128
rect 40764 53119 40822 53125
rect 44174 53116 44180 53128
rect 44232 53116 44238 53168
rect 45548 53159 45606 53165
rect 45548 53125 45560 53159
rect 45594 53156 45606 53159
rect 46658 53156 46664 53168
rect 45594 53128 46664 53156
rect 45594 53125 45606 53128
rect 45548 53119 45606 53125
rect 46658 53116 46664 53128
rect 46716 53116 46722 53168
rect 56220 53159 56278 53165
rect 56220 53125 56232 53159
rect 56266 53156 56278 53159
rect 58158 53156 58164 53168
rect 56266 53128 58164 53156
rect 56266 53125 56278 53128
rect 56220 53119 56278 53125
rect 58158 53116 58164 53128
rect 58216 53116 58222 53168
rect 3973 53091 4031 53097
rect 3973 53088 3985 53091
rect 3436 53060 3985 53088
rect 3973 53057 3985 53060
rect 4019 53057 4031 53091
rect 3973 53051 4031 53057
rect 6270 53048 6276 53100
rect 6328 53088 6334 53100
rect 6549 53091 6607 53097
rect 6549 53088 6561 53091
rect 6328 53060 6561 53088
rect 6328 53048 6334 53060
rect 6549 53057 6561 53060
rect 6595 53057 6607 53091
rect 6549 53051 6607 53057
rect 16669 53091 16727 53097
rect 16669 53057 16681 53091
rect 16715 53088 16727 53091
rect 18506 53088 18512 53100
rect 16715 53060 18512 53088
rect 16715 53057 16727 53060
rect 16669 53051 16727 53057
rect 18506 53048 18512 53060
rect 18564 53048 18570 53100
rect 18598 53048 18604 53100
rect 18656 53088 18662 53100
rect 18765 53091 18823 53097
rect 18765 53088 18777 53091
rect 18656 53060 18777 53088
rect 18656 53048 18662 53060
rect 18765 53057 18777 53060
rect 18811 53057 18823 53091
rect 18765 53051 18823 53057
rect 23201 53091 23259 53097
rect 23201 53057 23213 53091
rect 23247 53088 23259 53091
rect 24854 53088 24860 53100
rect 23247 53060 24860 53088
rect 23247 53057 23259 53060
rect 23201 53051 23259 53057
rect 24854 53048 24860 53060
rect 24912 53048 24918 53100
rect 25038 53088 25044 53100
rect 24999 53060 25044 53088
rect 25038 53048 25044 53060
rect 25096 53048 25102 53100
rect 25308 53091 25366 53097
rect 25308 53057 25320 53091
rect 25354 53088 25366 53091
rect 26234 53088 26240 53100
rect 25354 53060 26240 53088
rect 25354 53057 25366 53060
rect 25308 53051 25366 53057
rect 26234 53048 26240 53060
rect 26292 53048 26298 53100
rect 29454 53088 29460 53100
rect 29415 53060 29460 53088
rect 29454 53048 29460 53060
rect 29512 53048 29518 53100
rect 32125 53091 32183 53097
rect 32125 53057 32137 53091
rect 32171 53088 32183 53091
rect 33962 53088 33968 53100
rect 32171 53060 33968 53088
rect 32171 53057 32183 53060
rect 32125 53051 32183 53057
rect 33962 53048 33968 53060
rect 34020 53088 34026 53100
rect 34698 53088 34704 53100
rect 34020 53060 34704 53088
rect 34020 53048 34026 53060
rect 34698 53048 34704 53060
rect 34756 53048 34762 53100
rect 37918 53048 37924 53100
rect 37976 53088 37982 53100
rect 38657 53091 38715 53097
rect 38657 53088 38669 53091
rect 37976 53060 38669 53088
rect 37976 53048 37982 53060
rect 38657 53057 38669 53060
rect 38703 53088 38715 53091
rect 40494 53088 40500 53100
rect 38703 53060 40500 53088
rect 38703 53057 38715 53060
rect 38657 53051 38715 53057
rect 40494 53048 40500 53060
rect 40552 53048 40558 53100
rect 43708 53091 43766 53097
rect 43708 53057 43720 53091
rect 43754 53088 43766 53091
rect 47848 53091 47906 53097
rect 43754 53060 46704 53088
rect 43754 53057 43766 53060
rect 43708 53051 43766 53057
rect 43441 53023 43499 53029
rect 43441 52989 43453 53023
rect 43487 52989 43499 53023
rect 45278 53020 45284 53032
rect 45191 52992 45284 53020
rect 43441 52983 43499 52989
rect 17402 52844 17408 52896
rect 17460 52884 17466 52896
rect 18049 52887 18107 52893
rect 18049 52884 18061 52887
rect 17460 52856 18061 52884
rect 17460 52844 17466 52856
rect 18049 52853 18061 52856
rect 18095 52853 18107 52887
rect 18049 52847 18107 52853
rect 24581 52887 24639 52893
rect 24581 52853 24593 52887
rect 24627 52884 24639 52887
rect 26786 52884 26792 52896
rect 24627 52856 26792 52884
rect 24627 52853 24639 52856
rect 24581 52847 24639 52853
rect 26786 52844 26792 52856
rect 26844 52844 26850 52896
rect 35342 52884 35348 52896
rect 35303 52856 35348 52884
rect 35342 52844 35348 52856
rect 35400 52844 35406 52896
rect 43070 52844 43076 52896
rect 43128 52884 43134 52896
rect 43456 52884 43484 52983
rect 45278 52980 45284 52992
rect 45336 52980 45342 53032
rect 45296 52884 45324 52980
rect 46676 52961 46704 53060
rect 47848 53057 47860 53091
rect 47894 53088 47906 53091
rect 48314 53088 48320 53100
rect 47894 53060 48320 53088
rect 47894 53057 47906 53060
rect 47848 53051 47906 53057
rect 48314 53048 48320 53060
rect 48372 53048 48378 53100
rect 52914 53048 52920 53100
rect 52972 53088 52978 53100
rect 53653 53091 53711 53097
rect 53653 53088 53665 53091
rect 52972 53060 53665 53088
rect 52972 53048 52978 53060
rect 53653 53057 53665 53060
rect 53699 53057 53711 53091
rect 53653 53051 53711 53057
rect 53920 53091 53978 53097
rect 53920 53057 53932 53091
rect 53966 53088 53978 53091
rect 54754 53088 54760 53100
rect 53966 53060 54760 53088
rect 53966 53057 53978 53060
rect 53920 53051 53978 53057
rect 54754 53048 54760 53060
rect 54812 53048 54818 53100
rect 55950 53088 55956 53100
rect 55911 53060 55956 53088
rect 55950 53048 55956 53060
rect 56008 53048 56014 53100
rect 47578 53020 47584 53032
rect 47539 52992 47584 53020
rect 47578 52980 47584 52992
rect 47636 52980 47642 53032
rect 46661 52955 46719 52961
rect 46661 52921 46673 52955
rect 46707 52921 46719 52955
rect 46661 52915 46719 52921
rect 45462 52884 45468 52896
rect 43128 52856 45468 52884
rect 43128 52844 43134 52856
rect 45462 52844 45468 52856
rect 45520 52844 45526 52896
rect 1104 52794 59340 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 59340 52794
rect 1104 52720 59340 52742
rect 3234 52680 3240 52692
rect 3195 52652 3240 52680
rect 3234 52640 3240 52652
rect 3292 52640 3298 52692
rect 5810 52680 5816 52692
rect 5771 52652 5816 52680
rect 5810 52640 5816 52652
rect 5868 52640 5874 52692
rect 9490 52680 9496 52692
rect 9140 52652 9496 52680
rect 9140 52553 9168 52652
rect 9490 52640 9496 52652
rect 9548 52640 9554 52692
rect 18509 52683 18567 52689
rect 18509 52649 18521 52683
rect 18555 52680 18567 52683
rect 18598 52680 18604 52692
rect 18555 52652 18604 52680
rect 18555 52649 18567 52652
rect 18509 52643 18567 52649
rect 18598 52640 18604 52652
rect 18656 52640 18662 52692
rect 26234 52640 26240 52692
rect 26292 52680 26298 52692
rect 34054 52680 34060 52692
rect 26292 52652 26337 52680
rect 34015 52652 34060 52680
rect 26292 52640 26298 52652
rect 34054 52640 34060 52652
rect 34112 52640 34118 52692
rect 41782 52680 41788 52692
rect 41743 52652 41788 52680
rect 41782 52640 41788 52652
rect 41840 52640 41846 52692
rect 44358 52640 44364 52692
rect 44416 52680 44422 52692
rect 44453 52683 44511 52689
rect 44453 52680 44465 52683
rect 44416 52652 44465 52680
rect 44416 52640 44422 52652
rect 44453 52649 44465 52652
rect 44499 52649 44511 52683
rect 48314 52680 48320 52692
rect 48275 52652 48320 52680
rect 44453 52643 44511 52649
rect 48314 52640 48320 52652
rect 48372 52640 48378 52692
rect 54754 52680 54760 52692
rect 54715 52652 54760 52680
rect 54754 52640 54760 52652
rect 54812 52640 54818 52692
rect 57698 52680 57704 52692
rect 57659 52652 57704 52680
rect 57698 52640 57704 52652
rect 57756 52640 57762 52692
rect 10134 52572 10140 52624
rect 10192 52612 10198 52624
rect 10505 52615 10563 52621
rect 10505 52612 10517 52615
rect 10192 52584 10517 52612
rect 10192 52572 10198 52584
rect 10505 52581 10517 52584
rect 10551 52581 10563 52615
rect 10505 52575 10563 52581
rect 23014 52572 23020 52624
rect 23072 52612 23078 52624
rect 23201 52615 23259 52621
rect 23201 52612 23213 52615
rect 23072 52584 23213 52612
rect 23072 52572 23078 52584
rect 23201 52581 23213 52584
rect 23247 52581 23259 52615
rect 23201 52575 23259 52581
rect 9125 52547 9183 52553
rect 9125 52513 9137 52547
rect 9171 52513 9183 52547
rect 24854 52544 24860 52556
rect 24815 52516 24860 52544
rect 9125 52507 9183 52513
rect 24854 52504 24860 52516
rect 24912 52504 24918 52556
rect 43070 52544 43076 52556
rect 43031 52516 43076 52544
rect 43070 52504 43076 52516
rect 43128 52504 43134 52556
rect 55950 52504 55956 52556
rect 56008 52544 56014 52556
rect 56321 52547 56379 52553
rect 56321 52544 56333 52547
rect 56008 52516 56333 52544
rect 56008 52504 56014 52516
rect 56321 52513 56333 52516
rect 56367 52513 56379 52547
rect 56321 52507 56379 52513
rect 1578 52436 1584 52488
rect 1636 52476 1642 52488
rect 1857 52479 1915 52485
rect 1857 52476 1869 52479
rect 1636 52448 1869 52476
rect 1636 52436 1642 52448
rect 1857 52445 1869 52448
rect 1903 52445 1915 52479
rect 1857 52439 1915 52445
rect 2124 52479 2182 52485
rect 2124 52445 2136 52479
rect 2170 52476 2182 52479
rect 3418 52476 3424 52488
rect 2170 52448 3424 52476
rect 2170 52445 2182 52448
rect 2124 52439 2182 52445
rect 3418 52436 3424 52448
rect 3476 52436 3482 52488
rect 4433 52479 4491 52485
rect 4433 52445 4445 52479
rect 4479 52476 4491 52479
rect 4700 52479 4758 52485
rect 4479 52448 4660 52476
rect 4479 52445 4491 52448
rect 4433 52439 4491 52445
rect 4632 52420 4660 52448
rect 4700 52445 4712 52479
rect 4746 52476 4758 52479
rect 7006 52476 7012 52488
rect 4746 52448 7012 52476
rect 4746 52445 4758 52448
rect 4700 52439 4758 52445
rect 7006 52436 7012 52448
rect 7064 52436 7070 52488
rect 9392 52479 9450 52485
rect 9392 52445 9404 52479
rect 9438 52476 9450 52479
rect 10962 52476 10968 52488
rect 9438 52448 10968 52476
rect 9438 52445 9450 52448
rect 9392 52439 9450 52445
rect 10962 52436 10968 52448
rect 11020 52436 11026 52488
rect 11517 52479 11575 52485
rect 11517 52445 11529 52479
rect 11563 52476 11575 52479
rect 11606 52476 11612 52488
rect 11563 52448 11612 52476
rect 11563 52445 11575 52448
rect 11517 52439 11575 52445
rect 11606 52436 11612 52448
rect 11664 52436 11670 52488
rect 11784 52479 11842 52485
rect 11784 52445 11796 52479
rect 11830 52476 11842 52479
rect 13078 52476 13084 52488
rect 11830 52448 13084 52476
rect 11830 52445 11842 52448
rect 11784 52439 11842 52445
rect 13078 52436 13084 52448
rect 13136 52436 13142 52488
rect 14090 52476 14096 52488
rect 14003 52448 14096 52476
rect 14090 52436 14096 52448
rect 14148 52476 14154 52488
rect 14642 52476 14648 52488
rect 14148 52448 14648 52476
rect 14148 52436 14154 52448
rect 14642 52436 14648 52448
rect 14700 52436 14706 52488
rect 16666 52436 16672 52488
rect 16724 52476 16730 52488
rect 17402 52485 17408 52488
rect 17129 52479 17187 52485
rect 17129 52476 17141 52479
rect 16724 52448 17141 52476
rect 16724 52436 16730 52448
rect 17129 52445 17141 52448
rect 17175 52445 17187 52479
rect 17396 52476 17408 52485
rect 17363 52448 17408 52476
rect 17129 52439 17187 52445
rect 17396 52439 17408 52448
rect 17402 52436 17408 52439
rect 17460 52436 17466 52488
rect 19981 52479 20039 52485
rect 19981 52445 19993 52479
rect 20027 52476 20039 52479
rect 20248 52479 20306 52485
rect 20027 52448 20208 52476
rect 20027 52445 20039 52448
rect 19981 52439 20039 52445
rect 4614 52368 4620 52420
rect 4672 52368 4678 52420
rect 13814 52368 13820 52420
rect 13872 52408 13878 52420
rect 14338 52411 14396 52417
rect 14338 52408 14350 52411
rect 13872 52380 14350 52408
rect 13872 52368 13878 52380
rect 14338 52377 14350 52380
rect 14384 52377 14396 52411
rect 20180 52408 20208 52448
rect 20248 52445 20260 52479
rect 20294 52476 20306 52479
rect 20622 52476 20628 52488
rect 20294 52448 20628 52476
rect 20294 52445 20306 52448
rect 20248 52439 20306 52445
rect 20622 52436 20628 52448
rect 20680 52436 20686 52488
rect 21726 52436 21732 52488
rect 21784 52476 21790 52488
rect 21821 52479 21879 52485
rect 21821 52476 21833 52479
rect 21784 52448 21833 52476
rect 21784 52436 21790 52448
rect 21821 52445 21833 52448
rect 21867 52445 21879 52479
rect 21821 52439 21879 52445
rect 22088 52479 22146 52485
rect 22088 52445 22100 52479
rect 22134 52476 22146 52479
rect 23750 52476 23756 52488
rect 22134 52448 23756 52476
rect 22134 52445 22146 52448
rect 22088 52439 22146 52445
rect 23750 52436 23756 52448
rect 23808 52436 23814 52488
rect 25124 52479 25182 52485
rect 25124 52445 25136 52479
rect 25170 52476 25182 52479
rect 25682 52476 25688 52488
rect 25170 52448 25688 52476
rect 25170 52445 25182 52448
rect 25124 52439 25182 52445
rect 25682 52436 25688 52448
rect 25740 52436 25746 52488
rect 26697 52479 26755 52485
rect 26697 52445 26709 52479
rect 26743 52445 26755 52479
rect 26697 52439 26755 52445
rect 20806 52408 20812 52420
rect 20180 52380 20812 52408
rect 14338 52371 14396 52377
rect 20806 52368 20812 52380
rect 20864 52368 20870 52420
rect 24854 52368 24860 52420
rect 24912 52408 24918 52420
rect 26712 52408 26740 52439
rect 26786 52436 26792 52488
rect 26844 52476 26850 52488
rect 26953 52479 27011 52485
rect 26953 52476 26965 52479
rect 26844 52448 26965 52476
rect 26844 52436 26850 52448
rect 26953 52445 26965 52448
rect 26999 52445 27011 52479
rect 26953 52439 27011 52445
rect 32677 52479 32735 52485
rect 32677 52445 32689 52479
rect 32723 52445 32735 52479
rect 32677 52439 32735 52445
rect 32944 52479 33002 52485
rect 32944 52445 32956 52479
rect 32990 52476 33002 52479
rect 33226 52476 33232 52488
rect 32990 52448 33232 52476
rect 32990 52445 33002 52448
rect 32944 52439 33002 52445
rect 32692 52408 32720 52439
rect 33226 52436 33232 52448
rect 33284 52436 33290 52488
rect 39850 52436 39856 52488
rect 39908 52476 39914 52488
rect 40405 52479 40463 52485
rect 40405 52476 40417 52479
rect 39908 52448 40417 52476
rect 39908 52436 39914 52448
rect 40405 52445 40417 52448
rect 40451 52445 40463 52479
rect 40405 52439 40463 52445
rect 40672 52479 40730 52485
rect 40672 52445 40684 52479
rect 40718 52476 40730 52479
rect 41414 52476 41420 52488
rect 40718 52448 41420 52476
rect 40718 52445 40730 52448
rect 40672 52439 40730 52445
rect 41414 52436 41420 52448
rect 41472 52436 41478 52488
rect 43340 52479 43398 52485
rect 43340 52445 43352 52479
rect 43386 52476 43398 52479
rect 45186 52476 45192 52488
rect 43386 52448 45192 52476
rect 43386 52445 43398 52448
rect 43340 52439 43398 52445
rect 45186 52436 45192 52448
rect 45244 52436 45250 52488
rect 45462 52436 45468 52488
rect 45520 52476 45526 52488
rect 46937 52479 46995 52485
rect 45520 52436 45554 52476
rect 46937 52445 46949 52479
rect 46983 52445 46995 52479
rect 46937 52439 46995 52445
rect 47204 52479 47262 52485
rect 47204 52445 47216 52479
rect 47250 52476 47262 52479
rect 48958 52476 48964 52488
rect 47250 52448 48964 52476
rect 47250 52445 47262 52448
rect 47204 52439 47262 52445
rect 45526 52408 45554 52436
rect 46952 52408 46980 52439
rect 48958 52436 48964 52448
rect 49016 52436 49022 52488
rect 51350 52485 51356 52488
rect 51077 52479 51135 52485
rect 51077 52445 51089 52479
rect 51123 52476 51135 52479
rect 51344 52476 51356 52485
rect 51123 52448 51212 52476
rect 51311 52448 51356 52476
rect 51123 52445 51135 52448
rect 51077 52439 51135 52445
rect 47578 52408 47584 52420
rect 24912 52380 27016 52408
rect 32692 52380 33272 52408
rect 45526 52380 47584 52408
rect 24912 52368 24918 52380
rect 26988 52352 27016 52380
rect 33244 52352 33272 52380
rect 47578 52368 47584 52380
rect 47636 52368 47642 52420
rect 51184 52408 51212 52448
rect 51344 52439 51356 52448
rect 51350 52436 51356 52439
rect 51408 52436 51414 52488
rect 53098 52476 53104 52488
rect 51460 52448 53104 52476
rect 51460 52408 51488 52448
rect 53098 52436 53104 52448
rect 53156 52476 53162 52488
rect 53377 52479 53435 52485
rect 53377 52476 53389 52479
rect 53156 52448 53389 52476
rect 53156 52436 53162 52448
rect 53377 52445 53389 52448
rect 53423 52445 53435 52479
rect 53377 52439 53435 52445
rect 53644 52479 53702 52485
rect 53644 52445 53656 52479
rect 53690 52476 53702 52479
rect 54478 52476 54484 52488
rect 53690 52448 54484 52476
rect 53690 52445 53702 52448
rect 53644 52439 53702 52445
rect 54478 52436 54484 52448
rect 54536 52436 54542 52488
rect 51184 52380 51488 52408
rect 56588 52411 56646 52417
rect 56588 52377 56600 52411
rect 56634 52408 56646 52411
rect 57330 52408 57336 52420
rect 56634 52380 57336 52408
rect 56634 52377 56646 52380
rect 56588 52371 56646 52377
rect 57330 52368 57336 52380
rect 57388 52368 57394 52420
rect 12894 52340 12900 52352
rect 12855 52312 12900 52340
rect 12894 52300 12900 52312
rect 12952 52300 12958 52352
rect 15194 52300 15200 52352
rect 15252 52340 15258 52352
rect 15473 52343 15531 52349
rect 15473 52340 15485 52343
rect 15252 52312 15485 52340
rect 15252 52300 15258 52312
rect 15473 52309 15485 52312
rect 15519 52309 15531 52343
rect 21358 52340 21364 52352
rect 21319 52312 21364 52340
rect 15473 52303 15531 52309
rect 21358 52300 21364 52312
rect 21416 52300 21422 52352
rect 26970 52300 26976 52352
rect 27028 52300 27034 52352
rect 28074 52340 28080 52352
rect 28035 52312 28080 52340
rect 28074 52300 28080 52312
rect 28132 52300 28138 52352
rect 33226 52300 33232 52352
rect 33284 52300 33290 52352
rect 52454 52340 52460 52352
rect 52415 52312 52460 52340
rect 52454 52300 52460 52312
rect 52512 52300 52518 52352
rect 1104 52250 59340 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 59340 52250
rect 1104 52176 59340 52198
rect 3418 52136 3424 52148
rect 3379 52108 3424 52136
rect 3418 52096 3424 52108
rect 3476 52096 3482 52148
rect 10962 52136 10968 52148
rect 10923 52108 10968 52136
rect 10962 52096 10968 52108
rect 11020 52096 11026 52148
rect 13354 52136 13360 52148
rect 13315 52108 13360 52136
rect 13354 52096 13360 52108
rect 13412 52096 13418 52148
rect 20625 52139 20683 52145
rect 20625 52105 20637 52139
rect 20671 52136 20683 52139
rect 20714 52136 20720 52148
rect 20671 52108 20720 52136
rect 20671 52105 20683 52108
rect 20625 52099 20683 52105
rect 20714 52096 20720 52108
rect 20772 52096 20778 52148
rect 40310 52136 40316 52148
rect 40223 52108 40316 52136
rect 40310 52096 40316 52108
rect 40368 52136 40374 52148
rect 41690 52136 41696 52148
rect 40368 52108 41696 52136
rect 40368 52096 40374 52108
rect 41690 52096 41696 52108
rect 41748 52136 41754 52148
rect 43070 52136 43076 52148
rect 41748 52108 43076 52136
rect 41748 52096 41754 52108
rect 43070 52096 43076 52108
rect 43128 52096 43134 52148
rect 44542 52136 44548 52148
rect 44503 52108 44548 52136
rect 44542 52096 44548 52108
rect 44600 52096 44606 52148
rect 46845 52139 46903 52145
rect 46845 52105 46857 52139
rect 46891 52136 46903 52139
rect 47118 52136 47124 52148
rect 46891 52108 47124 52136
rect 46891 52105 46903 52108
rect 46845 52099 46903 52105
rect 47118 52096 47124 52108
rect 47176 52096 47182 52148
rect 48958 52136 48964 52148
rect 48919 52108 48964 52136
rect 48958 52096 48964 52108
rect 49016 52096 49022 52148
rect 54478 52136 54484 52148
rect 54439 52108 54484 52136
rect 54478 52096 54484 52108
rect 54536 52096 54542 52148
rect 57330 52136 57336 52148
rect 57291 52108 57336 52136
rect 57330 52096 57336 52108
rect 57388 52096 57394 52148
rect 7006 52068 7012 52080
rect 6564 52040 7012 52068
rect 2308 52003 2366 52009
rect 2308 51969 2320 52003
rect 2354 52000 2366 52003
rect 3234 52000 3240 52012
rect 2354 51972 3240 52000
rect 2354 51969 2366 51972
rect 2308 51963 2366 51969
rect 3234 51960 3240 51972
rect 3292 51960 3298 52012
rect 6564 52009 6592 52040
rect 7006 52028 7012 52040
rect 7064 52028 7070 52080
rect 11784 52071 11842 52077
rect 9600 52040 11560 52068
rect 6549 52003 6607 52009
rect 6549 51969 6561 52003
rect 6595 51969 6607 52003
rect 6549 51963 6607 51969
rect 6816 52003 6874 52009
rect 6816 51969 6828 52003
rect 6862 52000 6874 52003
rect 8386 52000 8392 52012
rect 6862 51972 8392 52000
rect 6862 51969 6874 51972
rect 6816 51963 6874 51969
rect 8386 51960 8392 51972
rect 8444 51960 8450 52012
rect 9600 52009 9628 52040
rect 9585 52003 9643 52009
rect 9585 51969 9597 52003
rect 9631 51969 9643 52003
rect 9585 51963 9643 51969
rect 9852 52003 9910 52009
rect 9852 51969 9864 52003
rect 9898 52000 9910 52003
rect 10962 52000 10968 52012
rect 9898 51972 10968 52000
rect 9898 51969 9910 51972
rect 9852 51963 9910 51969
rect 10962 51960 10968 51972
rect 11020 51960 11026 52012
rect 11532 52009 11560 52040
rect 11784 52037 11796 52071
rect 11830 52068 11842 52071
rect 12894 52068 12900 52080
rect 11830 52040 12900 52068
rect 11830 52037 11842 52040
rect 11784 52031 11842 52037
rect 12894 52028 12900 52040
rect 12952 52028 12958 52080
rect 19512 52071 19570 52077
rect 19512 52037 19524 52071
rect 19558 52068 19570 52071
rect 21358 52068 21364 52080
rect 19558 52040 21364 52068
rect 19558 52037 19570 52040
rect 19512 52031 19570 52037
rect 21358 52028 21364 52040
rect 21416 52028 21422 52080
rect 27240 52071 27298 52077
rect 27240 52037 27252 52071
rect 27286 52068 27298 52071
rect 28074 52068 28080 52080
rect 27286 52040 28080 52068
rect 27286 52037 27298 52040
rect 27240 52031 27298 52037
rect 28074 52028 28080 52040
rect 28132 52028 28138 52080
rect 33404 52071 33462 52077
rect 33404 52037 33416 52071
rect 33450 52068 33462 52071
rect 35342 52068 35348 52080
rect 33450 52040 35348 52068
rect 33450 52037 33462 52040
rect 33404 52031 33462 52037
rect 35342 52028 35348 52040
rect 35400 52028 35406 52080
rect 43432 52071 43490 52077
rect 43432 52037 43444 52071
rect 43478 52068 43490 52071
rect 44450 52068 44456 52080
rect 43478 52040 44456 52068
rect 43478 52037 43490 52040
rect 43432 52031 43490 52037
rect 44450 52028 44456 52040
rect 44508 52028 44514 52080
rect 51068 52071 51126 52077
rect 51068 52037 51080 52071
rect 51114 52068 51126 52071
rect 52454 52068 52460 52080
rect 51114 52040 52460 52068
rect 51114 52037 51126 52040
rect 51068 52031 51126 52037
rect 52454 52028 52460 52040
rect 52512 52028 52518 52080
rect 53116 52040 55214 52068
rect 53116 52012 53144 52040
rect 11517 52003 11575 52009
rect 11517 51969 11529 52003
rect 11563 52000 11575 52003
rect 11606 52000 11612 52012
rect 11563 51972 11612 52000
rect 11563 51969 11575 51972
rect 11517 51963 11575 51969
rect 11606 51960 11612 51972
rect 11664 51960 11670 52012
rect 13541 52003 13599 52009
rect 13541 51969 13553 52003
rect 13587 51969 13599 52003
rect 13541 51963 13599 51969
rect 1578 51892 1584 51944
rect 1636 51932 1642 51944
rect 2041 51935 2099 51941
rect 2041 51932 2053 51935
rect 1636 51904 2053 51932
rect 1636 51892 1642 51904
rect 2041 51901 2053 51904
rect 2087 51901 2099 51935
rect 13556 51932 13584 51963
rect 13630 51960 13636 52012
rect 13688 52000 13694 52012
rect 14349 52003 14407 52009
rect 14349 52000 14361 52003
rect 13688 51972 14361 52000
rect 13688 51960 13694 51972
rect 14349 51969 14361 51972
rect 14395 51969 14407 52003
rect 16666 52000 16672 52012
rect 16627 51972 16672 52000
rect 14349 51963 14407 51969
rect 16666 51960 16672 51972
rect 16724 51960 16730 52012
rect 16936 52003 16994 52009
rect 16936 51969 16948 52003
rect 16982 52000 16994 52003
rect 18046 52000 18052 52012
rect 16982 51972 18052 52000
rect 16982 51969 16994 51972
rect 16936 51963 16994 51969
rect 18046 51960 18052 51972
rect 18104 51960 18110 52012
rect 22088 52003 22146 52009
rect 22088 51969 22100 52003
rect 22134 52000 22146 52003
rect 23198 52000 23204 52012
rect 22134 51972 23204 52000
rect 22134 51969 22146 51972
rect 22088 51963 22146 51969
rect 23198 51960 23204 51972
rect 23256 51960 23262 52012
rect 23928 52003 23986 52009
rect 23928 51969 23940 52003
rect 23974 52000 23986 52003
rect 24486 52000 24492 52012
rect 23974 51972 24492 52000
rect 23974 51969 23986 51972
rect 23928 51963 23986 51969
rect 24486 51960 24492 51972
rect 24544 51960 24550 52012
rect 28813 52003 28871 52009
rect 28813 51969 28825 52003
rect 28859 52000 28871 52003
rect 28902 52000 28908 52012
rect 28859 51972 28908 52000
rect 28859 51969 28871 51972
rect 28813 51963 28871 51969
rect 28902 51960 28908 51972
rect 28960 51960 28966 52012
rect 29080 52003 29138 52009
rect 29080 51969 29092 52003
rect 29126 52000 29138 52003
rect 29914 52000 29920 52012
rect 29126 51972 29920 52000
rect 29126 51969 29138 51972
rect 29080 51963 29138 51969
rect 29914 51960 29920 51972
rect 29972 51960 29978 52012
rect 33137 52003 33195 52009
rect 33137 51969 33149 52003
rect 33183 52000 33195 52003
rect 33226 52000 33232 52012
rect 33183 51972 33232 52000
rect 33183 51969 33195 51972
rect 33137 51963 33195 51969
rect 33226 51960 33232 51972
rect 33284 51960 33290 52012
rect 34698 51960 34704 52012
rect 34756 52000 34762 52012
rect 35161 52003 35219 52009
rect 35161 52000 35173 52003
rect 34756 51972 35173 52000
rect 34756 51960 34762 51972
rect 35161 51969 35173 51972
rect 35207 51969 35219 52003
rect 35161 51963 35219 51969
rect 35428 52003 35486 52009
rect 35428 51969 35440 52003
rect 35474 52000 35486 52003
rect 35986 52000 35992 52012
rect 35474 51972 35992 52000
rect 35474 51969 35486 51972
rect 35428 51963 35486 51969
rect 35986 51960 35992 51972
rect 36044 51960 36050 52012
rect 38004 52003 38062 52009
rect 38004 51969 38016 52003
rect 38050 52000 38062 52003
rect 39942 52000 39948 52012
rect 38050 51972 39948 52000
rect 38050 51969 38062 51972
rect 38004 51963 38062 51969
rect 39942 51960 39948 51972
rect 40000 51960 40006 52012
rect 40497 52003 40555 52009
rect 40497 51969 40509 52003
rect 40543 52000 40555 52003
rect 40954 52000 40960 52012
rect 40543 51972 40960 52000
rect 40543 51969 40555 51972
rect 40497 51963 40555 51969
rect 40954 51960 40960 51972
rect 41012 52000 41018 52012
rect 47029 52003 47087 52009
rect 47029 52000 47041 52003
rect 41012 51972 47041 52000
rect 41012 51960 41018 51972
rect 47029 51969 47041 51972
rect 47075 51969 47087 52003
rect 47029 51963 47087 51969
rect 47848 52003 47906 52009
rect 47848 51969 47860 52003
rect 47894 52000 47906 52003
rect 49050 52000 49056 52012
rect 47894 51972 49056 52000
rect 47894 51969 47906 51972
rect 47848 51963 47906 51969
rect 49050 51960 49056 51972
rect 49108 51960 49114 52012
rect 53098 52000 53104 52012
rect 53059 51972 53104 52000
rect 53098 51960 53104 51972
rect 53156 51960 53162 52012
rect 53368 52003 53426 52009
rect 53368 51969 53380 52003
rect 53414 52000 53426 52003
rect 54294 52000 54300 52012
rect 53414 51972 54300 52000
rect 53414 51969 53426 51972
rect 53368 51963 53426 51969
rect 54294 51960 54300 51972
rect 54352 51960 54358 52012
rect 55186 52000 55214 52040
rect 55950 52000 55956 52012
rect 55186 51972 55956 52000
rect 55950 51960 55956 51972
rect 56008 51960 56014 52012
rect 56220 52003 56278 52009
rect 56220 51969 56232 52003
rect 56266 52000 56278 52003
rect 57146 52000 57152 52012
rect 56266 51972 57152 52000
rect 56266 51969 56278 51972
rect 56220 51963 56278 51969
rect 57146 51960 57152 51972
rect 57204 51960 57210 52012
rect 13998 51932 14004 51944
rect 13556 51904 14004 51932
rect 2041 51895 2099 51901
rect 13998 51892 14004 51904
rect 14056 51892 14062 51944
rect 14090 51892 14096 51944
rect 14148 51932 14154 51944
rect 19242 51932 19248 51944
rect 14148 51904 14193 51932
rect 19203 51904 19248 51932
rect 14148 51892 14154 51904
rect 19242 51892 19248 51904
rect 19300 51892 19306 51944
rect 21818 51932 21824 51944
rect 21779 51904 21824 51932
rect 21818 51892 21824 51904
rect 21876 51892 21882 51944
rect 23658 51932 23664 51944
rect 23619 51904 23664 51932
rect 23658 51892 23664 51904
rect 23716 51892 23722 51944
rect 26970 51932 26976 51944
rect 26931 51904 26976 51932
rect 26970 51892 26976 51904
rect 27028 51892 27034 51944
rect 37182 51892 37188 51944
rect 37240 51932 37246 51944
rect 37737 51935 37795 51941
rect 37737 51932 37749 51935
rect 37240 51904 37749 51932
rect 37240 51892 37246 51904
rect 37737 51901 37749 51904
rect 37783 51901 37795 51935
rect 43162 51932 43168 51944
rect 43123 51904 43168 51932
rect 37737 51895 37795 51901
rect 43162 51892 43168 51904
rect 43220 51892 43226 51944
rect 47578 51932 47584 51944
rect 47539 51904 47584 51932
rect 47578 51892 47584 51904
rect 47636 51892 47642 51944
rect 48774 51892 48780 51944
rect 48832 51932 48838 51944
rect 50801 51935 50859 51941
rect 50801 51932 50813 51935
rect 48832 51904 50813 51932
rect 48832 51892 48838 51904
rect 50801 51901 50813 51904
rect 50847 51901 50859 51935
rect 50801 51895 50859 51901
rect 12897 51867 12955 51873
rect 12897 51833 12909 51867
rect 12943 51864 12955 51867
rect 13814 51864 13820 51876
rect 12943 51836 13820 51864
rect 12943 51833 12955 51836
rect 12897 51827 12955 51833
rect 13814 51824 13820 51836
rect 13872 51824 13878 51876
rect 7926 51796 7932 51808
rect 7887 51768 7932 51796
rect 7926 51756 7932 51768
rect 7984 51756 7990 51808
rect 15470 51796 15476 51808
rect 15431 51768 15476 51796
rect 15470 51756 15476 51768
rect 15528 51756 15534 51808
rect 17770 51756 17776 51808
rect 17828 51796 17834 51808
rect 18049 51799 18107 51805
rect 18049 51796 18061 51799
rect 17828 51768 18061 51796
rect 17828 51756 17834 51768
rect 18049 51765 18061 51768
rect 18095 51765 18107 51799
rect 18049 51759 18107 51765
rect 23201 51799 23259 51805
rect 23201 51765 23213 51799
rect 23247 51796 23259 51799
rect 23934 51796 23940 51808
rect 23247 51768 23940 51796
rect 23247 51765 23259 51768
rect 23201 51759 23259 51765
rect 23934 51756 23940 51768
rect 23992 51756 23998 51808
rect 24946 51756 24952 51808
rect 25004 51796 25010 51808
rect 25041 51799 25099 51805
rect 25041 51796 25053 51799
rect 25004 51768 25053 51796
rect 25004 51756 25010 51768
rect 25041 51765 25053 51768
rect 25087 51765 25099 51799
rect 28350 51796 28356 51808
rect 28311 51768 28356 51796
rect 25041 51759 25099 51765
rect 28350 51756 28356 51768
rect 28408 51756 28414 51808
rect 30190 51796 30196 51808
rect 30151 51768 30196 51796
rect 30190 51756 30196 51768
rect 30248 51756 30254 51808
rect 33042 51756 33048 51808
rect 33100 51796 33106 51808
rect 34517 51799 34575 51805
rect 34517 51796 34529 51799
rect 33100 51768 34529 51796
rect 33100 51756 33106 51768
rect 34517 51765 34529 51768
rect 34563 51765 34575 51799
rect 34517 51759 34575 51765
rect 36541 51799 36599 51805
rect 36541 51765 36553 51799
rect 36587 51796 36599 51799
rect 36630 51796 36636 51808
rect 36587 51768 36636 51796
rect 36587 51765 36599 51768
rect 36541 51759 36599 51765
rect 36630 51756 36636 51768
rect 36688 51756 36694 51808
rect 39117 51799 39175 51805
rect 39117 51765 39129 51799
rect 39163 51796 39175 51799
rect 40126 51796 40132 51808
rect 39163 51768 40132 51796
rect 39163 51765 39175 51768
rect 39117 51759 39175 51765
rect 40126 51756 40132 51768
rect 40184 51756 40190 51808
rect 52178 51796 52184 51808
rect 52139 51768 52184 51796
rect 52178 51756 52184 51768
rect 52236 51756 52242 51808
rect 1104 51706 59340 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 59340 51706
rect 1104 51632 59340 51654
rect 3234 51592 3240 51604
rect 3195 51564 3240 51592
rect 3234 51552 3240 51564
rect 3292 51552 3298 51604
rect 8386 51592 8392 51604
rect 8347 51564 8392 51592
rect 8386 51552 8392 51564
rect 8444 51552 8450 51604
rect 13449 51595 13507 51601
rect 13449 51561 13461 51595
rect 13495 51592 13507 51595
rect 13630 51592 13636 51604
rect 13495 51564 13636 51592
rect 13495 51561 13507 51564
rect 13449 51555 13507 51561
rect 13630 51552 13636 51564
rect 13688 51552 13694 51604
rect 13998 51552 14004 51604
rect 14056 51592 14062 51604
rect 24762 51592 24768 51604
rect 14056 51564 20199 51592
rect 14056 51552 14062 51564
rect 19334 51484 19340 51536
rect 19392 51524 19398 51536
rect 19981 51527 20039 51533
rect 19981 51524 19993 51527
rect 19392 51496 19993 51524
rect 19392 51484 19398 51496
rect 19981 51493 19993 51496
rect 20027 51524 20039 51527
rect 20070 51524 20076 51536
rect 20027 51496 20076 51524
rect 20027 51493 20039 51496
rect 19981 51487 20039 51493
rect 20070 51484 20076 51496
rect 20128 51484 20134 51536
rect 20171 51524 20199 51564
rect 24412 51564 24768 51592
rect 20714 51524 20720 51536
rect 20171 51496 20720 51524
rect 14090 51456 14096 51468
rect 13832 51428 14096 51456
rect 1578 51348 1584 51400
rect 1636 51388 1642 51400
rect 1857 51391 1915 51397
rect 1857 51388 1869 51391
rect 1636 51360 1869 51388
rect 1636 51348 1642 51360
rect 1857 51357 1869 51360
rect 1903 51388 1915 51391
rect 4430 51388 4436 51400
rect 1903 51360 4436 51388
rect 1903 51357 1915 51360
rect 1857 51351 1915 51357
rect 4430 51348 4436 51360
rect 4488 51388 4494 51400
rect 5166 51388 5172 51400
rect 4488 51360 5172 51388
rect 4488 51348 4494 51360
rect 5166 51348 5172 51360
rect 5224 51348 5230 51400
rect 7006 51388 7012 51400
rect 6967 51360 7012 51388
rect 7006 51348 7012 51360
rect 7064 51348 7070 51400
rect 10229 51391 10287 51397
rect 10229 51357 10241 51391
rect 10275 51388 10287 51391
rect 11698 51388 11704 51400
rect 10275 51360 11704 51388
rect 10275 51357 10287 51360
rect 10229 51351 10287 51357
rect 11698 51348 11704 51360
rect 11756 51388 11762 51400
rect 12069 51391 12127 51397
rect 12069 51388 12081 51391
rect 11756 51360 12081 51388
rect 11756 51348 11762 51360
rect 12069 51357 12081 51360
rect 12115 51388 12127 51391
rect 13832 51388 13860 51428
rect 14090 51416 14096 51428
rect 14148 51416 14154 51468
rect 12115 51360 13860 51388
rect 14360 51391 14418 51397
rect 12115 51357 12127 51360
rect 12069 51351 12127 51357
rect 14360 51357 14372 51391
rect 14406 51388 14418 51391
rect 15470 51388 15476 51400
rect 14406 51360 15476 51388
rect 14406 51357 14418 51360
rect 14360 51351 14418 51357
rect 15470 51348 15476 51360
rect 15528 51348 15534 51400
rect 15933 51391 15991 51397
rect 15933 51357 15945 51391
rect 15979 51388 15991 51391
rect 16666 51388 16672 51400
rect 15979 51360 16672 51388
rect 15979 51357 15991 51360
rect 15933 51351 15991 51357
rect 16666 51348 16672 51360
rect 16724 51348 16730 51400
rect 20171 51397 20199 51496
rect 20714 51484 20720 51496
rect 20772 51484 20778 51536
rect 24412 51465 24440 51564
rect 24762 51552 24768 51564
rect 24820 51552 24826 51604
rect 49050 51592 49056 51604
rect 49011 51564 49056 51592
rect 49050 51552 49056 51564
rect 49108 51552 49114 51604
rect 54294 51592 54300 51604
rect 54255 51564 54300 51592
rect 54294 51552 54300 51564
rect 54352 51552 54358 51604
rect 55950 51552 55956 51604
rect 56008 51592 56014 51604
rect 57149 51595 57207 51601
rect 57149 51592 57161 51595
rect 56008 51564 57161 51592
rect 56008 51552 56014 51564
rect 57149 51561 57161 51564
rect 57195 51561 57207 51595
rect 57149 51555 57207 51561
rect 24397 51459 24455 51465
rect 24397 51425 24409 51459
rect 24443 51425 24455 51459
rect 39850 51456 39856 51468
rect 39811 51428 39856 51456
rect 24397 51419 24455 51425
rect 39850 51416 39856 51428
rect 39908 51416 39914 51468
rect 45554 51416 45560 51468
rect 45612 51456 45618 51468
rect 45833 51459 45891 51465
rect 45833 51456 45845 51459
rect 45612 51428 45845 51456
rect 45612 51416 45618 51428
rect 45833 51425 45845 51428
rect 45879 51425 45891 51459
rect 45833 51419 45891 51425
rect 20165 51391 20223 51397
rect 20165 51357 20177 51391
rect 20211 51357 20223 51391
rect 20165 51351 20223 51357
rect 20717 51391 20775 51397
rect 20717 51357 20729 51391
rect 20763 51388 20775 51391
rect 20806 51388 20812 51400
rect 20763 51360 20812 51388
rect 20763 51357 20775 51360
rect 20717 51351 20775 51357
rect 20806 51348 20812 51360
rect 20864 51388 20870 51400
rect 21818 51388 21824 51400
rect 20864 51360 21824 51388
rect 20864 51348 20870 51360
rect 21818 51348 21824 51360
rect 21876 51348 21882 51400
rect 25774 51348 25780 51400
rect 25832 51388 25838 51400
rect 27249 51391 27307 51397
rect 27249 51388 27261 51391
rect 25832 51360 27261 51388
rect 25832 51348 25838 51360
rect 27249 51357 27261 51360
rect 27295 51388 27307 51391
rect 27614 51388 27620 51400
rect 27295 51360 27620 51388
rect 27295 51357 27307 51360
rect 27249 51351 27307 51357
rect 27614 51348 27620 51360
rect 27672 51348 27678 51400
rect 29549 51391 29607 51397
rect 29549 51357 29561 51391
rect 29595 51388 29607 51391
rect 30098 51388 30104 51400
rect 29595 51360 30104 51388
rect 29595 51357 29607 51360
rect 29549 51351 29607 51357
rect 30098 51348 30104 51360
rect 30156 51388 30162 51400
rect 33042 51397 33048 51400
rect 32769 51391 32827 51397
rect 32769 51388 32781 51391
rect 30156 51360 32781 51388
rect 30156 51348 30162 51360
rect 32769 51357 32781 51360
rect 32815 51357 32827 51391
rect 33036 51388 33048 51397
rect 33003 51360 33048 51388
rect 32769 51351 32827 51357
rect 33036 51351 33048 51360
rect 2124 51323 2182 51329
rect 2124 51289 2136 51323
rect 2170 51320 2182 51323
rect 3418 51320 3424 51332
rect 2170 51292 3424 51320
rect 2170 51289 2182 51292
rect 2124 51283 2182 51289
rect 3418 51280 3424 51292
rect 3476 51280 3482 51332
rect 5436 51323 5494 51329
rect 5436 51289 5448 51323
rect 5482 51320 5494 51323
rect 6178 51320 6184 51332
rect 5482 51292 6184 51320
rect 5482 51289 5494 51292
rect 5436 51283 5494 51289
rect 6178 51280 6184 51292
rect 6236 51280 6242 51332
rect 7276 51323 7334 51329
rect 7276 51289 7288 51323
rect 7322 51320 7334 51323
rect 9122 51320 9128 51332
rect 7322 51292 9128 51320
rect 7322 51289 7334 51292
rect 7276 51283 7334 51289
rect 9122 51280 9128 51292
rect 9180 51280 9186 51332
rect 10496 51323 10554 51329
rect 10496 51289 10508 51323
rect 10542 51320 10554 51323
rect 12158 51320 12164 51332
rect 10542 51292 12164 51320
rect 10542 51289 10554 51292
rect 10496 51283 10554 51289
rect 12158 51280 12164 51292
rect 12216 51280 12222 51332
rect 12336 51323 12394 51329
rect 12336 51289 12348 51323
rect 12382 51320 12394 51323
rect 15194 51320 15200 51332
rect 12382 51292 15200 51320
rect 12382 51289 12394 51292
rect 12336 51283 12394 51289
rect 15194 51280 15200 51292
rect 15252 51280 15258 51332
rect 15562 51280 15568 51332
rect 15620 51320 15626 51332
rect 16178 51323 16236 51329
rect 16178 51320 16190 51323
rect 15620 51292 16190 51320
rect 15620 51280 15626 51292
rect 16178 51289 16190 51292
rect 16224 51289 16236 51323
rect 16178 51283 16236 51289
rect 20984 51323 21042 51329
rect 20984 51289 20996 51323
rect 21030 51320 21042 51323
rect 21266 51320 21272 51332
rect 21030 51292 21272 51320
rect 21030 51289 21042 51292
rect 20984 51283 21042 51289
rect 21266 51280 21272 51292
rect 21324 51280 21330 51332
rect 24664 51323 24722 51329
rect 24664 51289 24676 51323
rect 24710 51320 24722 51323
rect 25038 51320 25044 51332
rect 24710 51292 25044 51320
rect 24710 51289 24722 51292
rect 24664 51283 24722 51289
rect 25038 51280 25044 51292
rect 25096 51280 25102 51332
rect 29816 51323 29874 51329
rect 29816 51289 29828 51323
rect 29862 51320 29874 51323
rect 30466 51320 30472 51332
rect 29862 51292 30472 51320
rect 29862 51289 29874 51292
rect 29816 51283 29874 51289
rect 30466 51280 30472 51292
rect 30524 51280 30530 51332
rect 32784 51320 32812 51351
rect 33042 51348 33048 51351
rect 33100 51348 33106 51400
rect 34701 51391 34759 51397
rect 34701 51388 34713 51391
rect 34532 51360 34713 51388
rect 33226 51320 33232 51332
rect 32784 51292 33232 51320
rect 33226 51280 33232 51292
rect 33284 51320 33290 51332
rect 34532 51320 34560 51360
rect 34701 51357 34713 51360
rect 34747 51357 34759 51391
rect 36538 51388 36544 51400
rect 36451 51360 36544 51388
rect 34701 51351 34759 51357
rect 36538 51348 36544 51360
rect 36596 51388 36602 51400
rect 37182 51388 37188 51400
rect 36596 51360 37188 51388
rect 36596 51348 36602 51360
rect 37182 51348 37188 51360
rect 37240 51348 37246 51400
rect 47578 51348 47584 51400
rect 47636 51388 47642 51400
rect 47673 51391 47731 51397
rect 47673 51388 47685 51391
rect 47636 51360 47685 51388
rect 47636 51348 47642 51360
rect 47673 51357 47685 51360
rect 47719 51357 47731 51391
rect 47673 51351 47731 51357
rect 50614 51348 50620 51400
rect 50672 51388 50678 51400
rect 50893 51391 50951 51397
rect 50893 51388 50905 51391
rect 50672 51360 50905 51388
rect 50672 51348 50678 51360
rect 50893 51357 50905 51360
rect 50939 51357 50951 51391
rect 50893 51351 50951 51357
rect 51160 51391 51218 51397
rect 51160 51357 51172 51391
rect 51206 51388 51218 51391
rect 52178 51388 52184 51400
rect 51206 51360 52184 51388
rect 51206 51357 51218 51360
rect 51160 51351 51218 51357
rect 52178 51348 52184 51360
rect 52236 51348 52242 51400
rect 52917 51391 52975 51397
rect 52917 51357 52929 51391
rect 52963 51388 52975 51391
rect 53006 51388 53012 51400
rect 52963 51360 53012 51388
rect 52963 51357 52975 51360
rect 52917 51351 52975 51357
rect 53006 51348 53012 51360
rect 53064 51348 53070 51400
rect 53184 51391 53242 51397
rect 53184 51357 53196 51391
rect 53230 51388 53242 51391
rect 58526 51388 58532 51400
rect 53230 51360 58532 51388
rect 53230 51357 53242 51360
rect 53184 51351 53242 51357
rect 58526 51348 58532 51360
rect 58584 51348 58590 51400
rect 33284 51292 34560 51320
rect 33284 51280 33290 51292
rect 34606 51280 34612 51332
rect 34664 51320 34670 51332
rect 34946 51323 35004 51329
rect 34946 51320 34958 51323
rect 34664 51292 34958 51320
rect 34664 51280 34670 51292
rect 34946 51289 34958 51292
rect 34992 51289 35004 51323
rect 34946 51283 35004 51289
rect 36808 51323 36866 51329
rect 36808 51289 36820 51323
rect 36854 51320 36866 51323
rect 37826 51320 37832 51332
rect 36854 51292 37832 51320
rect 36854 51289 36866 51292
rect 36808 51283 36866 51289
rect 37826 51280 37832 51292
rect 37884 51280 37890 51332
rect 40120 51323 40178 51329
rect 40120 51289 40132 51323
rect 40166 51320 40178 51323
rect 41138 51320 41144 51332
rect 40166 51292 41144 51320
rect 40166 51289 40178 51292
rect 40120 51283 40178 51289
rect 41138 51280 41144 51292
rect 41196 51280 41202 51332
rect 46100 51323 46158 51329
rect 46100 51289 46112 51323
rect 46146 51320 46158 51323
rect 47762 51320 47768 51332
rect 46146 51292 47768 51320
rect 46146 51289 46158 51292
rect 46100 51283 46158 51289
rect 47762 51280 47768 51292
rect 47820 51280 47826 51332
rect 47940 51323 47998 51329
rect 47940 51289 47952 51323
rect 47986 51320 47998 51323
rect 48958 51320 48964 51332
rect 47986 51292 48964 51320
rect 47986 51289 47998 51292
rect 47940 51283 47998 51289
rect 48958 51280 48964 51292
rect 49016 51280 49022 51332
rect 55861 51323 55919 51329
rect 55861 51289 55873 51323
rect 55907 51320 55919 51323
rect 56042 51320 56048 51332
rect 55907 51292 56048 51320
rect 55907 51289 55919 51292
rect 55861 51283 55919 51289
rect 56042 51280 56048 51292
rect 56100 51280 56106 51332
rect 6546 51252 6552 51264
rect 6507 51224 6552 51252
rect 6546 51212 6552 51224
rect 6604 51212 6610 51264
rect 11606 51252 11612 51264
rect 11567 51224 11612 51252
rect 11606 51212 11612 51224
rect 11664 51212 11670 51264
rect 15470 51252 15476 51264
rect 15431 51224 15476 51252
rect 15470 51212 15476 51224
rect 15528 51212 15534 51264
rect 17310 51252 17316 51264
rect 17271 51224 17316 51252
rect 17310 51212 17316 51224
rect 17368 51212 17374 51264
rect 20070 51212 20076 51264
rect 20128 51252 20134 51264
rect 21174 51252 21180 51264
rect 20128 51224 21180 51252
rect 20128 51212 20134 51224
rect 21174 51212 21180 51224
rect 21232 51212 21238 51264
rect 22094 51252 22100 51264
rect 22055 51224 22100 51252
rect 22094 51212 22100 51224
rect 22152 51212 22158 51264
rect 23474 51212 23480 51264
rect 23532 51252 23538 51264
rect 25777 51255 25835 51261
rect 25777 51252 25789 51255
rect 23532 51224 25789 51252
rect 23532 51212 23538 51224
rect 25777 51221 25789 51224
rect 25823 51221 25835 51255
rect 25777 51215 25835 51221
rect 28721 51255 28779 51261
rect 28721 51221 28733 51255
rect 28767 51252 28779 51255
rect 28902 51252 28908 51264
rect 28767 51224 28908 51252
rect 28767 51221 28779 51224
rect 28721 51215 28779 51221
rect 28902 51212 28908 51224
rect 28960 51212 28966 51264
rect 30282 51212 30288 51264
rect 30340 51252 30346 51264
rect 30929 51255 30987 51261
rect 30929 51252 30941 51255
rect 30340 51224 30941 51252
rect 30340 51212 30346 51224
rect 30929 51221 30941 51224
rect 30975 51221 30987 51255
rect 34146 51252 34152 51264
rect 34107 51224 34152 51252
rect 30929 51215 30987 51221
rect 34146 51212 34152 51224
rect 34204 51212 34210 51264
rect 36078 51252 36084 51264
rect 36039 51224 36084 51252
rect 36078 51212 36084 51224
rect 36136 51212 36142 51264
rect 37918 51252 37924 51264
rect 37879 51224 37924 51252
rect 37918 51212 37924 51224
rect 37976 51212 37982 51264
rect 41233 51255 41291 51261
rect 41233 51221 41245 51255
rect 41279 51252 41291 51255
rect 41782 51252 41788 51264
rect 41279 51224 41788 51252
rect 41279 51221 41291 51224
rect 41233 51215 41291 51221
rect 41782 51212 41788 51224
rect 41840 51212 41846 51264
rect 47210 51252 47216 51264
rect 47171 51224 47216 51252
rect 47210 51212 47216 51224
rect 47268 51212 47274 51264
rect 52270 51252 52276 51264
rect 52231 51224 52276 51252
rect 52270 51212 52276 51224
rect 52328 51212 52334 51264
rect 1104 51162 59340 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 59340 51162
rect 1104 51088 59340 51110
rect 3418 51048 3424 51060
rect 3379 51020 3424 51048
rect 3418 51008 3424 51020
rect 3476 51008 3482 51060
rect 9122 51048 9128 51060
rect 9083 51020 9128 51048
rect 9122 51008 9128 51020
rect 9180 51008 9186 51060
rect 10962 51048 10968 51060
rect 10923 51020 10968 51048
rect 10962 51008 10968 51020
rect 11020 51008 11026 51060
rect 12158 51008 12164 51060
rect 12216 51048 12222 51060
rect 13081 51051 13139 51057
rect 13081 51048 13093 51051
rect 12216 51020 13093 51048
rect 12216 51008 12222 51020
rect 13081 51017 13093 51020
rect 13127 51017 13139 51051
rect 18046 51048 18052 51060
rect 18007 51020 18052 51048
rect 13081 51011 13139 51017
rect 18046 51008 18052 51020
rect 18104 51008 18110 51060
rect 21266 51048 21272 51060
rect 21227 51020 21272 51048
rect 21266 51008 21272 51020
rect 21324 51008 21330 51060
rect 23198 51048 23204 51060
rect 23159 51020 23204 51048
rect 23198 51008 23204 51020
rect 23256 51008 23262 51060
rect 25038 51048 25044 51060
rect 24999 51020 25044 51048
rect 25038 51008 25044 51020
rect 25096 51008 25102 51060
rect 34606 51048 34612 51060
rect 34567 51020 34612 51048
rect 34606 51008 34612 51020
rect 34664 51008 34670 51060
rect 39942 51008 39948 51060
rect 40000 51048 40006 51060
rect 40497 51051 40555 51057
rect 40497 51048 40509 51051
rect 40000 51020 40509 51048
rect 40000 51008 40006 51020
rect 40497 51017 40509 51020
rect 40543 51017 40555 51051
rect 48958 51048 48964 51060
rect 48919 51020 48964 51048
rect 40497 51011 40555 51017
rect 48958 51008 48964 51020
rect 49016 51008 49022 51060
rect 57146 51048 57152 51060
rect 57107 51020 57152 51048
rect 57146 51008 57152 51020
rect 57204 51008 57210 51060
rect 4700 50983 4758 50989
rect 4700 50949 4712 50983
rect 4746 50980 4758 50983
rect 6546 50980 6552 50992
rect 4746 50952 6552 50980
rect 4746 50949 4758 50952
rect 4700 50943 4758 50949
rect 6546 50940 6552 50952
rect 6604 50940 6610 50992
rect 9852 50983 9910 50989
rect 9852 50949 9864 50983
rect 9898 50980 9910 50983
rect 11606 50980 11612 50992
rect 9898 50952 11612 50980
rect 9898 50949 9910 50952
rect 9852 50943 9910 50949
rect 11606 50940 11612 50952
rect 11664 50940 11670 50992
rect 14360 50983 14418 50989
rect 14360 50949 14372 50983
rect 14406 50980 14418 50983
rect 15470 50980 15476 50992
rect 14406 50952 15476 50980
rect 14406 50949 14418 50952
rect 14360 50943 14418 50949
rect 15470 50940 15476 50952
rect 15528 50940 15534 50992
rect 22094 50989 22100 50992
rect 22088 50980 22100 50989
rect 22055 50952 22100 50980
rect 22088 50943 22100 50952
rect 22094 50940 22100 50943
rect 22152 50940 22158 50992
rect 23934 50989 23940 50992
rect 23928 50980 23940 50989
rect 23895 50952 23940 50980
rect 23928 50943 23940 50952
rect 23934 50940 23940 50943
rect 23992 50940 23998 50992
rect 27240 50983 27298 50989
rect 27240 50949 27252 50983
rect 27286 50980 27298 50983
rect 28350 50980 28356 50992
rect 27286 50952 28356 50980
rect 27286 50949 27298 50952
rect 27240 50943 27298 50949
rect 28350 50940 28356 50952
rect 28408 50940 28414 50992
rect 30098 50980 30104 50992
rect 28828 50952 30104 50980
rect 2308 50915 2366 50921
rect 2308 50881 2320 50915
rect 2354 50912 2366 50915
rect 3234 50912 3240 50924
rect 2354 50884 3240 50912
rect 2354 50881 2366 50884
rect 2308 50875 2366 50881
rect 3234 50872 3240 50884
rect 3292 50872 3298 50924
rect 4430 50912 4436 50924
rect 4391 50884 4436 50912
rect 4430 50872 4436 50884
rect 4488 50872 4494 50924
rect 8012 50915 8070 50921
rect 8012 50881 8024 50915
rect 8058 50912 8070 50915
rect 10134 50912 10140 50924
rect 8058 50884 10140 50912
rect 8058 50881 8070 50884
rect 8012 50875 8070 50881
rect 10134 50872 10140 50884
rect 10192 50872 10198 50924
rect 11238 50872 11244 50924
rect 11296 50912 11302 50924
rect 11957 50915 12015 50921
rect 11957 50912 11969 50915
rect 11296 50884 11969 50912
rect 11296 50872 11302 50884
rect 11957 50881 11969 50884
rect 12003 50881 12015 50915
rect 11957 50875 12015 50881
rect 16936 50915 16994 50921
rect 16936 50881 16948 50915
rect 16982 50912 16994 50915
rect 17402 50912 17408 50924
rect 16982 50884 17408 50912
rect 16982 50881 16994 50884
rect 16936 50875 16994 50881
rect 17402 50872 17408 50884
rect 17460 50872 17466 50924
rect 20156 50915 20214 50921
rect 20156 50881 20168 50915
rect 20202 50912 20214 50915
rect 23106 50912 23112 50924
rect 20202 50884 23112 50912
rect 20202 50881 20214 50884
rect 20156 50875 20214 50881
rect 23106 50872 23112 50884
rect 23164 50872 23170 50924
rect 23658 50912 23664 50924
rect 23619 50884 23664 50912
rect 23658 50872 23664 50884
rect 23716 50872 23722 50924
rect 1578 50804 1584 50856
rect 1636 50844 1642 50856
rect 2041 50847 2099 50853
rect 2041 50844 2053 50847
rect 1636 50816 2053 50844
rect 1636 50804 1642 50816
rect 2041 50813 2053 50816
rect 2087 50813 2099 50847
rect 2041 50807 2099 50813
rect 7745 50847 7803 50853
rect 7745 50813 7757 50847
rect 7791 50813 7803 50847
rect 7745 50807 7803 50813
rect 9585 50847 9643 50853
rect 9585 50813 9597 50847
rect 9631 50813 9643 50847
rect 11698 50844 11704 50856
rect 11659 50816 11704 50844
rect 9585 50807 9643 50813
rect 5810 50708 5816 50720
rect 5771 50680 5816 50708
rect 5810 50668 5816 50680
rect 5868 50668 5874 50720
rect 7760 50708 7788 50807
rect 8110 50708 8116 50720
rect 7760 50680 8116 50708
rect 8110 50668 8116 50680
rect 8168 50708 8174 50720
rect 9600 50708 9628 50807
rect 11698 50804 11704 50816
rect 11756 50804 11762 50856
rect 14090 50844 14096 50856
rect 14051 50816 14096 50844
rect 14090 50804 14096 50816
rect 14148 50804 14154 50856
rect 16666 50844 16672 50856
rect 16579 50816 16672 50844
rect 16666 50804 16672 50816
rect 16724 50804 16730 50856
rect 19889 50847 19947 50853
rect 19889 50813 19901 50847
rect 19935 50813 19947 50847
rect 19889 50807 19947 50813
rect 21821 50847 21879 50853
rect 21821 50813 21833 50847
rect 21867 50813 21879 50847
rect 26970 50844 26976 50856
rect 26931 50816 26976 50844
rect 21821 50807 21879 50813
rect 15470 50708 15476 50720
rect 8168 50680 9628 50708
rect 15431 50680 15476 50708
rect 8168 50668 8174 50680
rect 15470 50668 15476 50680
rect 15528 50668 15534 50720
rect 16684 50708 16712 50804
rect 17034 50708 17040 50720
rect 16684 50680 17040 50708
rect 17034 50668 17040 50680
rect 17092 50708 17098 50720
rect 19242 50708 19248 50720
rect 17092 50680 19248 50708
rect 17092 50668 17098 50680
rect 19242 50668 19248 50680
rect 19300 50668 19306 50720
rect 19904 50708 19932 50807
rect 20070 50708 20076 50720
rect 19904 50680 20076 50708
rect 20070 50668 20076 50680
rect 20128 50708 20134 50720
rect 21836 50708 21864 50807
rect 26970 50804 26976 50816
rect 27028 50804 27034 50856
rect 28828 50853 28856 50952
rect 30098 50940 30104 50952
rect 30156 50940 30162 50992
rect 33496 50983 33554 50989
rect 33496 50949 33508 50983
rect 33542 50980 33554 50983
rect 34146 50980 34152 50992
rect 33542 50952 34152 50980
rect 33542 50949 33554 50952
rect 33496 50943 33554 50949
rect 34146 50940 34152 50952
rect 34204 50940 34210 50992
rect 35336 50983 35394 50989
rect 35336 50949 35348 50983
rect 35382 50980 35394 50983
rect 36078 50980 36084 50992
rect 35382 50952 36084 50980
rect 35382 50949 35394 50952
rect 35336 50943 35394 50949
rect 36078 50940 36084 50952
rect 36136 50940 36142 50992
rect 37544 50983 37602 50989
rect 37544 50949 37556 50983
rect 37590 50980 37602 50983
rect 37918 50980 37924 50992
rect 37590 50952 37924 50980
rect 37590 50949 37602 50952
rect 37544 50943 37602 50949
rect 37918 50940 37924 50952
rect 37976 50940 37982 50992
rect 43162 50980 43168 50992
rect 42444 50952 43168 50980
rect 28902 50872 28908 50924
rect 28960 50912 28966 50924
rect 29069 50915 29127 50921
rect 29069 50912 29081 50915
rect 28960 50884 29081 50912
rect 28960 50872 28966 50884
rect 29069 50881 29081 50884
rect 29115 50881 29127 50915
rect 33226 50912 33232 50924
rect 33187 50884 33232 50912
rect 29069 50875 29127 50881
rect 33226 50872 33232 50884
rect 33284 50872 33290 50924
rect 35069 50915 35127 50921
rect 35069 50881 35081 50915
rect 35115 50912 35127 50915
rect 36538 50912 36544 50924
rect 35115 50884 36544 50912
rect 35115 50881 35127 50884
rect 35069 50875 35127 50881
rect 36538 50872 36544 50884
rect 36596 50872 36602 50924
rect 37182 50872 37188 50924
rect 37240 50912 37246 50924
rect 37277 50915 37335 50921
rect 37277 50912 37289 50915
rect 37240 50884 37289 50912
rect 37240 50872 37246 50884
rect 37277 50881 37289 50884
rect 37323 50881 37335 50915
rect 37277 50875 37335 50881
rect 38746 50872 38752 50924
rect 38804 50912 38810 50924
rect 39373 50915 39431 50921
rect 39373 50912 39385 50915
rect 38804 50884 39385 50912
rect 38804 50872 38810 50884
rect 39373 50881 39385 50884
rect 39419 50881 39431 50915
rect 39373 50875 39431 50881
rect 28813 50847 28871 50853
rect 28813 50813 28825 50847
rect 28859 50813 28871 50847
rect 28813 50807 28871 50813
rect 39117 50847 39175 50853
rect 39117 50813 39129 50847
rect 39163 50813 39175 50847
rect 39117 50807 39175 50813
rect 22462 50708 22468 50720
rect 20128 50680 22468 50708
rect 20128 50668 20134 50680
rect 22462 50668 22468 50680
rect 22520 50708 22526 50720
rect 23658 50708 23664 50720
rect 22520 50680 23664 50708
rect 22520 50668 22526 50680
rect 23658 50668 23664 50680
rect 23716 50668 23722 50720
rect 28350 50708 28356 50720
rect 28311 50680 28356 50708
rect 28350 50668 28356 50680
rect 28408 50668 28414 50720
rect 29086 50668 29092 50720
rect 29144 50708 29150 50720
rect 30193 50711 30251 50717
rect 30193 50708 30205 50711
rect 29144 50680 30205 50708
rect 29144 50668 29150 50680
rect 30193 50677 30205 50680
rect 30239 50677 30251 50711
rect 36446 50708 36452 50720
rect 36407 50680 36452 50708
rect 30193 50671 30251 50677
rect 36446 50668 36452 50680
rect 36504 50668 36510 50720
rect 38654 50708 38660 50720
rect 38615 50680 38660 50708
rect 38654 50668 38660 50680
rect 38712 50668 38718 50720
rect 39132 50708 39160 50807
rect 41690 50804 41696 50856
rect 41748 50844 41754 50856
rect 42444 50853 42472 50952
rect 43162 50940 43168 50952
rect 43220 50980 43226 50992
rect 43220 50952 44312 50980
rect 43220 50940 43226 50952
rect 44284 50924 44312 50952
rect 47210 50940 47216 50992
rect 47268 50980 47274 50992
rect 47826 50983 47884 50989
rect 47826 50980 47838 50983
rect 47268 50952 47838 50980
rect 47268 50940 47274 50952
rect 47826 50949 47838 50952
rect 47872 50949 47884 50983
rect 47826 50943 47884 50949
rect 51068 50983 51126 50989
rect 51068 50949 51080 50983
rect 51114 50980 51126 50983
rect 52270 50980 52276 50992
rect 51114 50952 52276 50980
rect 51114 50949 51126 50952
rect 51068 50943 51126 50949
rect 52270 50940 52276 50952
rect 52328 50940 52334 50992
rect 55950 50940 55956 50992
rect 56008 50940 56014 50992
rect 42696 50915 42754 50921
rect 42696 50881 42708 50915
rect 42742 50912 42754 50915
rect 43714 50912 43720 50924
rect 42742 50884 43720 50912
rect 42742 50881 42754 50884
rect 42696 50875 42754 50881
rect 43714 50872 43720 50884
rect 43772 50872 43778 50924
rect 44266 50912 44272 50924
rect 44179 50884 44272 50912
rect 44266 50872 44272 50884
rect 44324 50872 44330 50924
rect 44536 50915 44594 50921
rect 44536 50881 44548 50915
rect 44582 50912 44594 50915
rect 46382 50912 46388 50924
rect 44582 50884 46388 50912
rect 44582 50881 44594 50884
rect 44536 50875 44594 50881
rect 46382 50872 46388 50884
rect 46440 50872 46446 50924
rect 55769 50915 55827 50921
rect 55769 50881 55781 50915
rect 55815 50912 55827 50915
rect 55968 50912 55996 50940
rect 55815 50884 55996 50912
rect 56036 50915 56094 50921
rect 55815 50881 55827 50884
rect 55769 50875 55827 50881
rect 56036 50881 56048 50915
rect 56082 50912 56094 50915
rect 57422 50912 57428 50924
rect 56082 50884 57428 50912
rect 56082 50881 56094 50884
rect 56036 50875 56094 50881
rect 57422 50872 57428 50884
rect 57480 50872 57486 50924
rect 42429 50847 42487 50853
rect 42429 50844 42441 50847
rect 41748 50816 42441 50844
rect 41748 50804 41754 50816
rect 42429 50813 42441 50816
rect 42475 50813 42487 50847
rect 47578 50844 47584 50856
rect 47539 50816 47584 50844
rect 42429 50807 42487 50813
rect 47578 50804 47584 50816
rect 47636 50804 47642 50856
rect 50614 50804 50620 50856
rect 50672 50844 50678 50856
rect 50801 50847 50859 50853
rect 50801 50844 50813 50847
rect 50672 50816 50813 50844
rect 50672 50804 50678 50816
rect 50801 50813 50813 50816
rect 50847 50813 50859 50847
rect 50801 50807 50859 50813
rect 39850 50708 39856 50720
rect 39132 50680 39856 50708
rect 39850 50668 39856 50680
rect 39908 50668 39914 50720
rect 43806 50708 43812 50720
rect 43767 50680 43812 50708
rect 43806 50668 43812 50680
rect 43864 50668 43870 50720
rect 45646 50708 45652 50720
rect 45607 50680 45652 50708
rect 45646 50668 45652 50680
rect 45704 50668 45710 50720
rect 52178 50708 52184 50720
rect 52139 50680 52184 50708
rect 52178 50668 52184 50680
rect 52236 50668 52242 50720
rect 1104 50618 59340 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 59340 50618
rect 1104 50544 59340 50566
rect 3234 50504 3240 50516
rect 3195 50476 3240 50504
rect 3234 50464 3240 50476
rect 3292 50464 3298 50516
rect 5166 50464 5172 50516
rect 5224 50504 5230 50516
rect 5445 50507 5503 50513
rect 5445 50504 5457 50507
rect 5224 50476 5457 50504
rect 5224 50464 5230 50476
rect 5445 50473 5457 50476
rect 5491 50473 5503 50507
rect 5445 50467 5503 50473
rect 6178 50464 6184 50516
rect 6236 50504 6242 50516
rect 7745 50507 7803 50513
rect 7745 50504 7757 50507
rect 6236 50476 7757 50504
rect 6236 50464 6242 50476
rect 7745 50473 7757 50476
rect 7791 50473 7803 50507
rect 11238 50504 11244 50516
rect 11199 50476 11244 50504
rect 7745 50467 7803 50473
rect 11238 50464 11244 50476
rect 11296 50464 11302 50516
rect 14090 50464 14096 50516
rect 14148 50504 14154 50516
rect 15562 50504 15568 50516
rect 14148 50476 15148 50504
rect 15523 50476 15568 50504
rect 14148 50464 14154 50476
rect 14200 50377 14228 50476
rect 15120 50436 15148 50476
rect 15562 50464 15568 50476
rect 15620 50464 15626 50516
rect 17402 50504 17408 50516
rect 17363 50476 17408 50504
rect 17402 50464 17408 50476
rect 17460 50464 17466 50516
rect 23106 50504 23112 50516
rect 23067 50476 23112 50504
rect 23106 50464 23112 50476
rect 23164 50464 23170 50516
rect 25682 50464 25688 50516
rect 25740 50504 25746 50516
rect 25777 50507 25835 50513
rect 25777 50504 25789 50507
rect 25740 50476 25789 50504
rect 25740 50464 25746 50476
rect 25777 50473 25789 50476
rect 25823 50473 25835 50507
rect 25777 50467 25835 50473
rect 30466 50464 30472 50516
rect 30524 50504 30530 50516
rect 30929 50507 30987 50513
rect 30929 50504 30941 50507
rect 30524 50476 30941 50504
rect 30524 50464 30530 50476
rect 30929 50473 30941 50476
rect 30975 50473 30987 50507
rect 30929 50467 30987 50473
rect 37826 50464 37832 50516
rect 37884 50504 37890 50516
rect 37921 50507 37979 50513
rect 37921 50504 37933 50507
rect 37884 50476 37933 50504
rect 37884 50464 37890 50476
rect 37921 50473 37933 50476
rect 37967 50473 37979 50507
rect 37921 50467 37979 50473
rect 47762 50464 47768 50516
rect 47820 50504 47826 50516
rect 48225 50507 48283 50513
rect 48225 50504 48237 50507
rect 47820 50476 48237 50504
rect 47820 50464 47826 50476
rect 48225 50473 48237 50476
rect 48271 50473 48283 50507
rect 57422 50504 57428 50516
rect 57383 50476 57428 50504
rect 48225 50467 48283 50473
rect 57422 50464 57428 50476
rect 57480 50464 57486 50516
rect 15120 50408 16068 50436
rect 16040 50377 16068 50408
rect 6365 50371 6423 50377
rect 6365 50337 6377 50371
rect 6411 50368 6423 50371
rect 14185 50371 14243 50377
rect 6411 50340 6500 50368
rect 6411 50337 6423 50340
rect 6365 50331 6423 50337
rect 1578 50260 1584 50312
rect 1636 50300 1642 50312
rect 1857 50303 1915 50309
rect 1857 50300 1869 50303
rect 1636 50272 1869 50300
rect 1636 50260 1642 50272
rect 1857 50269 1869 50272
rect 1903 50269 1915 50303
rect 1857 50263 1915 50269
rect 4157 50303 4215 50309
rect 4157 50269 4169 50303
rect 4203 50300 4215 50303
rect 5534 50300 5540 50312
rect 4203 50272 5540 50300
rect 4203 50269 4215 50272
rect 4157 50263 4215 50269
rect 5534 50260 5540 50272
rect 5592 50260 5598 50312
rect 2124 50235 2182 50241
rect 2124 50201 2136 50235
rect 2170 50232 2182 50235
rect 2866 50232 2872 50244
rect 2170 50204 2872 50232
rect 2170 50201 2182 50204
rect 2124 50195 2182 50201
rect 2866 50192 2872 50204
rect 2924 50192 2930 50244
rect 6472 50232 6500 50340
rect 14185 50337 14197 50371
rect 14231 50337 14243 50371
rect 14185 50331 14243 50337
rect 16025 50371 16083 50377
rect 16025 50337 16037 50371
rect 16071 50337 16083 50371
rect 16025 50331 16083 50337
rect 19242 50328 19248 50380
rect 19300 50368 19306 50380
rect 19889 50371 19947 50377
rect 19889 50368 19901 50371
rect 19300 50340 19901 50368
rect 19300 50328 19306 50340
rect 19889 50337 19901 50340
rect 19935 50337 19947 50371
rect 21726 50368 21732 50380
rect 21687 50340 21732 50368
rect 19889 50331 19947 50337
rect 21726 50328 21732 50340
rect 21784 50328 21790 50380
rect 36538 50368 36544 50380
rect 36499 50340 36544 50368
rect 36538 50328 36544 50340
rect 36596 50328 36602 50380
rect 39850 50368 39856 50380
rect 39811 50340 39856 50368
rect 39850 50328 39856 50340
rect 39908 50328 39914 50380
rect 55950 50328 55956 50380
rect 56008 50368 56014 50380
rect 56045 50371 56103 50377
rect 56045 50368 56057 50371
rect 56008 50340 56057 50368
rect 56008 50328 56014 50340
rect 56045 50337 56057 50340
rect 56091 50337 56103 50371
rect 56045 50331 56103 50337
rect 6632 50303 6690 50309
rect 6632 50269 6644 50303
rect 6678 50300 6690 50303
rect 7926 50300 7932 50312
rect 6678 50272 7932 50300
rect 6678 50269 6690 50272
rect 6632 50263 6690 50269
rect 7926 50260 7932 50272
rect 7984 50260 7990 50312
rect 8938 50260 8944 50312
rect 8996 50300 9002 50312
rect 9861 50303 9919 50309
rect 9861 50300 9873 50303
rect 8996 50272 9873 50300
rect 8996 50260 9002 50272
rect 9861 50269 9873 50272
rect 9907 50269 9919 50303
rect 9861 50263 9919 50269
rect 12161 50303 12219 50309
rect 12161 50269 12173 50303
rect 12207 50300 12219 50303
rect 13814 50300 13820 50312
rect 12207 50272 13820 50300
rect 12207 50269 12219 50272
rect 12161 50263 12219 50269
rect 13814 50260 13820 50272
rect 13872 50260 13878 50312
rect 14452 50303 14510 50309
rect 14452 50269 14464 50303
rect 14498 50300 14510 50303
rect 15470 50300 15476 50312
rect 14498 50272 15476 50300
rect 14498 50269 14510 50272
rect 14452 50263 14510 50269
rect 15470 50260 15476 50272
rect 15528 50260 15534 50312
rect 16292 50303 16350 50309
rect 16292 50269 16304 50303
rect 16338 50300 16350 50303
rect 17310 50300 17316 50312
rect 16338 50272 17316 50300
rect 16338 50269 16350 50272
rect 16292 50263 16350 50269
rect 17310 50260 17316 50272
rect 17368 50260 17374 50312
rect 21744 50300 21772 50328
rect 24397 50303 24455 50309
rect 24397 50300 24409 50303
rect 21744 50272 24409 50300
rect 24397 50269 24409 50272
rect 24443 50269 24455 50303
rect 24397 50263 24455 50269
rect 24664 50303 24722 50309
rect 24664 50269 24676 50303
rect 24710 50300 24722 50303
rect 24946 50300 24952 50312
rect 24710 50272 24952 50300
rect 24710 50269 24722 50272
rect 24664 50263 24722 50269
rect 7006 50232 7012 50244
rect 6472 50204 7012 50232
rect 6362 50124 6368 50176
rect 6420 50164 6426 50176
rect 6472 50164 6500 50204
rect 7006 50192 7012 50204
rect 7064 50232 7070 50244
rect 8110 50232 8116 50244
rect 7064 50204 8116 50232
rect 7064 50192 7070 50204
rect 8110 50192 8116 50204
rect 8168 50192 8174 50244
rect 10128 50235 10186 50241
rect 10128 50201 10140 50235
rect 10174 50232 10186 50235
rect 10778 50232 10784 50244
rect 10174 50204 10784 50232
rect 10174 50201 10186 50204
rect 10128 50195 10186 50201
rect 10778 50192 10784 50204
rect 10836 50192 10842 50244
rect 12428 50235 12486 50241
rect 12428 50201 12440 50235
rect 12474 50232 12486 50235
rect 16114 50232 16120 50244
rect 12474 50204 16120 50232
rect 12474 50201 12486 50204
rect 12428 50195 12486 50201
rect 16114 50192 16120 50204
rect 16172 50192 16178 50244
rect 20156 50235 20214 50241
rect 20156 50201 20168 50235
rect 20202 50232 20214 50235
rect 21082 50232 21088 50244
rect 20202 50204 21088 50232
rect 20202 50201 20214 50204
rect 20156 50195 20214 50201
rect 21082 50192 21088 50204
rect 21140 50192 21146 50244
rect 21974 50235 22032 50241
rect 21974 50232 21986 50235
rect 21284 50204 21986 50232
rect 13538 50164 13544 50176
rect 6420 50136 6500 50164
rect 13499 50136 13544 50164
rect 6420 50124 6426 50136
rect 13538 50124 13544 50136
rect 13596 50124 13602 50176
rect 21284 50173 21312 50204
rect 21974 50201 21986 50204
rect 22020 50201 22032 50235
rect 24412 50232 24440 50263
rect 24946 50260 24952 50272
rect 25004 50260 25010 50312
rect 26970 50300 26976 50312
rect 26931 50272 26976 50300
rect 26970 50260 26976 50272
rect 27028 50260 27034 50312
rect 27240 50303 27298 50309
rect 27240 50269 27252 50303
rect 27286 50300 27298 50303
rect 28350 50300 28356 50312
rect 27286 50272 28356 50300
rect 27286 50269 27298 50272
rect 27240 50263 27298 50269
rect 28350 50260 28356 50272
rect 28408 50260 28414 50312
rect 28994 50260 29000 50312
rect 29052 50300 29058 50312
rect 29546 50300 29552 50312
rect 29052 50272 29552 50300
rect 29052 50260 29058 50272
rect 29546 50260 29552 50272
rect 29604 50260 29610 50312
rect 29816 50303 29874 50309
rect 29816 50269 29828 50303
rect 29862 50300 29874 50303
rect 30190 50300 30196 50312
rect 29862 50272 30196 50300
rect 29862 50269 29874 50272
rect 29816 50263 29874 50269
rect 30190 50260 30196 50272
rect 30248 50260 30254 50312
rect 31389 50303 31447 50309
rect 31389 50300 31401 50303
rect 31220 50272 31401 50300
rect 24854 50232 24860 50244
rect 24412 50204 24860 50232
rect 21974 50195 22032 50201
rect 24854 50192 24860 50204
rect 24912 50192 24918 50244
rect 30098 50192 30104 50244
rect 30156 50232 30162 50244
rect 31220 50232 31248 50272
rect 31389 50269 31401 50272
rect 31435 50269 31447 50303
rect 34698 50300 34704 50312
rect 34659 50272 34704 50300
rect 31389 50263 31447 50269
rect 34698 50260 34704 50272
rect 34756 50260 34762 50312
rect 34968 50303 35026 50309
rect 34968 50269 34980 50303
rect 35014 50300 35026 50303
rect 36446 50300 36452 50312
rect 35014 50272 36452 50300
rect 35014 50269 35026 50272
rect 34968 50263 35026 50269
rect 36446 50260 36452 50272
rect 36504 50260 36510 50312
rect 36630 50260 36636 50312
rect 36688 50300 36694 50312
rect 40126 50309 40132 50312
rect 36797 50303 36855 50309
rect 36797 50300 36809 50303
rect 36688 50272 36809 50300
rect 36688 50260 36694 50272
rect 36797 50269 36809 50272
rect 36843 50269 36855 50303
rect 40120 50300 40132 50309
rect 40087 50272 40132 50300
rect 36797 50263 36855 50269
rect 40120 50263 40132 50272
rect 40126 50260 40132 50263
rect 40184 50260 40190 50312
rect 41690 50300 41696 50312
rect 41651 50272 41696 50300
rect 41690 50260 41696 50272
rect 41748 50260 41754 50312
rect 41782 50260 41788 50312
rect 41840 50300 41846 50312
rect 41949 50303 42007 50309
rect 41949 50300 41961 50303
rect 41840 50272 41961 50300
rect 41840 50260 41846 50272
rect 41949 50269 41961 50272
rect 41995 50269 42007 50303
rect 41949 50263 42007 50269
rect 44266 50260 44272 50312
rect 44324 50300 44330 50312
rect 45005 50303 45063 50309
rect 45005 50300 45017 50303
rect 44324 50272 45017 50300
rect 44324 50260 44330 50272
rect 45005 50269 45017 50272
rect 45051 50269 45063 50303
rect 45005 50263 45063 50269
rect 46845 50303 46903 50309
rect 46845 50269 46857 50303
rect 46891 50300 46903 50303
rect 47578 50300 47584 50312
rect 46891 50272 47584 50300
rect 46891 50269 46903 50272
rect 46845 50263 46903 50269
rect 47578 50260 47584 50272
rect 47636 50260 47642 50312
rect 50614 50260 50620 50312
rect 50672 50300 50678 50312
rect 50709 50303 50767 50309
rect 50709 50300 50721 50303
rect 50672 50272 50721 50300
rect 50672 50260 50678 50272
rect 50709 50269 50721 50272
rect 50755 50269 50767 50303
rect 50709 50263 50767 50269
rect 50976 50303 51034 50309
rect 50976 50269 50988 50303
rect 51022 50300 51034 50303
rect 52178 50300 52184 50312
rect 51022 50272 52184 50300
rect 51022 50269 51034 50272
rect 50976 50263 51034 50269
rect 52178 50260 52184 50272
rect 52236 50260 52242 50312
rect 30156 50204 31248 50232
rect 30156 50192 30162 50204
rect 31294 50192 31300 50244
rect 31352 50232 31358 50244
rect 31634 50235 31692 50241
rect 31634 50232 31646 50235
rect 31352 50204 31646 50232
rect 31352 50192 31358 50204
rect 31634 50201 31646 50204
rect 31680 50201 31692 50235
rect 31634 50195 31692 50201
rect 45272 50235 45330 50241
rect 45272 50201 45284 50235
rect 45318 50232 45330 50235
rect 46290 50232 46296 50244
rect 45318 50204 46296 50232
rect 45318 50201 45330 50204
rect 45272 50195 45330 50201
rect 46290 50192 46296 50204
rect 46348 50192 46354 50244
rect 47090 50235 47148 50241
rect 47090 50232 47102 50235
rect 46400 50204 47102 50232
rect 21269 50167 21327 50173
rect 21269 50133 21281 50167
rect 21315 50133 21327 50167
rect 28350 50164 28356 50176
rect 28311 50136 28356 50164
rect 21269 50127 21327 50133
rect 28350 50124 28356 50136
rect 28408 50124 28414 50176
rect 32766 50164 32772 50176
rect 32727 50136 32772 50164
rect 32766 50124 32772 50136
rect 32824 50124 32830 50176
rect 36078 50164 36084 50176
rect 36039 50136 36084 50164
rect 36078 50124 36084 50136
rect 36136 50124 36142 50176
rect 41230 50164 41236 50176
rect 41191 50136 41236 50164
rect 41230 50124 41236 50136
rect 41288 50124 41294 50176
rect 41414 50124 41420 50176
rect 41472 50164 41478 50176
rect 46400 50173 46428 50204
rect 47090 50201 47102 50204
rect 47136 50201 47148 50235
rect 47090 50195 47148 50201
rect 56312 50235 56370 50241
rect 56312 50201 56324 50235
rect 56358 50232 56370 50235
rect 56594 50232 56600 50244
rect 56358 50204 56600 50232
rect 56358 50201 56370 50204
rect 56312 50195 56370 50201
rect 56594 50192 56600 50204
rect 56652 50192 56658 50244
rect 43073 50167 43131 50173
rect 43073 50164 43085 50167
rect 41472 50136 43085 50164
rect 41472 50124 41478 50136
rect 43073 50133 43085 50136
rect 43119 50133 43131 50167
rect 43073 50127 43131 50133
rect 46385 50167 46443 50173
rect 46385 50133 46397 50167
rect 46431 50133 46443 50167
rect 52086 50164 52092 50176
rect 52047 50136 52092 50164
rect 46385 50127 46443 50133
rect 52086 50124 52092 50136
rect 52144 50124 52150 50176
rect 1104 50074 59340 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 59340 50074
rect 1104 50000 59340 50022
rect 16114 49960 16120 49972
rect 16075 49932 16120 49960
rect 16114 49920 16120 49932
rect 16172 49920 16178 49972
rect 21082 49960 21088 49972
rect 21043 49932 21088 49960
rect 21082 49920 21088 49932
rect 21140 49920 21146 49972
rect 24486 49960 24492 49972
rect 24447 49932 24492 49960
rect 24486 49920 24492 49932
rect 24544 49920 24550 49972
rect 26234 49920 26240 49972
rect 26292 49960 26298 49972
rect 26329 49963 26387 49969
rect 26329 49960 26341 49963
rect 26292 49932 26341 49960
rect 26292 49920 26298 49932
rect 26329 49929 26341 49932
rect 26375 49929 26387 49963
rect 26329 49923 26387 49929
rect 29914 49920 29920 49972
rect 29972 49960 29978 49972
rect 30193 49963 30251 49969
rect 30193 49960 30205 49963
rect 29972 49932 30205 49960
rect 29972 49920 29978 49932
rect 30193 49929 30205 49932
rect 30239 49929 30251 49963
rect 30193 49923 30251 49929
rect 33226 49920 33232 49972
rect 33284 49960 33290 49972
rect 33781 49963 33839 49969
rect 33781 49960 33793 49963
rect 33284 49932 33793 49960
rect 33284 49920 33290 49932
rect 33781 49929 33793 49932
rect 33827 49929 33839 49963
rect 33781 49923 33839 49929
rect 44266 49920 44272 49972
rect 44324 49960 44330 49972
rect 44453 49963 44511 49969
rect 44453 49960 44465 49963
rect 44324 49932 44465 49960
rect 44324 49920 44330 49932
rect 44453 49929 44465 49932
rect 44499 49929 44511 49963
rect 51997 49963 52055 49969
rect 51997 49960 52009 49963
rect 44453 49923 44511 49929
rect 50264 49932 52009 49960
rect 5810 49852 5816 49904
rect 5868 49892 5874 49904
rect 6610 49895 6668 49901
rect 6610 49892 6622 49895
rect 5868 49864 6622 49892
rect 5868 49852 5874 49864
rect 6610 49861 6622 49864
rect 6656 49861 6668 49895
rect 6610 49855 6668 49861
rect 13164 49895 13222 49901
rect 13164 49861 13176 49895
rect 13210 49892 13222 49895
rect 16022 49892 16028 49904
rect 13210 49864 16028 49892
rect 13210 49861 13222 49864
rect 13164 49855 13222 49861
rect 16022 49852 16028 49864
rect 16080 49852 16086 49904
rect 18785 49895 18843 49901
rect 18785 49861 18797 49895
rect 18831 49892 18843 49895
rect 19242 49892 19248 49904
rect 18831 49864 19248 49892
rect 18831 49861 18843 49864
rect 18785 49855 18843 49861
rect 19242 49852 19248 49864
rect 19300 49852 19306 49904
rect 20070 49892 20076 49904
rect 19720 49864 20076 49892
rect 19720 49836 19748 49864
rect 20070 49852 20076 49864
rect 20128 49852 20134 49904
rect 23376 49895 23434 49901
rect 23376 49861 23388 49895
rect 23422 49892 23434 49895
rect 23474 49892 23480 49904
rect 23422 49864 23480 49892
rect 23422 49861 23434 49864
rect 23376 49855 23434 49861
rect 23474 49852 23480 49864
rect 23532 49852 23538 49904
rect 27240 49895 27298 49901
rect 27240 49861 27252 49895
rect 27286 49892 27298 49895
rect 28350 49892 28356 49904
rect 27286 49864 28356 49892
rect 27286 49861 27298 49864
rect 27240 49855 27298 49861
rect 28350 49852 28356 49864
rect 28408 49852 28414 49904
rect 29086 49901 29092 49904
rect 29080 49892 29092 49901
rect 29047 49864 29092 49892
rect 29080 49855 29092 49864
rect 29086 49852 29092 49855
rect 29144 49852 29150 49904
rect 32490 49892 32496 49904
rect 32451 49864 32496 49892
rect 32490 49852 32496 49864
rect 32548 49892 32554 49904
rect 34790 49892 34796 49904
rect 32548 49864 34796 49892
rect 32548 49852 32554 49864
rect 34790 49852 34796 49864
rect 34848 49852 34854 49904
rect 34968 49895 35026 49901
rect 34968 49861 34980 49895
rect 35014 49892 35026 49895
rect 36078 49892 36084 49904
rect 35014 49864 36084 49892
rect 35014 49861 35026 49864
rect 34968 49855 35026 49861
rect 36078 49852 36084 49864
rect 36136 49852 36142 49904
rect 37544 49895 37602 49901
rect 37544 49861 37556 49895
rect 37590 49892 37602 49895
rect 38654 49892 38660 49904
rect 37590 49864 38660 49892
rect 37590 49861 37602 49864
rect 37544 49855 37602 49861
rect 38654 49852 38660 49864
rect 38712 49852 38718 49904
rect 39384 49895 39442 49901
rect 39384 49861 39396 49895
rect 39430 49892 39442 49895
rect 41230 49892 41236 49904
rect 39430 49864 41236 49892
rect 39430 49861 39442 49864
rect 39384 49855 39442 49861
rect 41230 49852 41236 49864
rect 41288 49852 41294 49904
rect 43070 49852 43076 49904
rect 43128 49892 43134 49904
rect 43165 49895 43223 49901
rect 43165 49892 43177 49895
rect 43128 49864 43177 49892
rect 43128 49852 43134 49864
rect 43165 49861 43177 49864
rect 43211 49861 43223 49895
rect 43165 49855 43223 49861
rect 43806 49852 43812 49904
rect 43864 49892 43870 49904
rect 45618 49895 45676 49901
rect 45618 49892 45630 49895
rect 43864 49864 45630 49892
rect 43864 49852 43870 49864
rect 45618 49861 45630 49864
rect 45664 49861 45676 49895
rect 45618 49855 45676 49861
rect 49044 49895 49102 49901
rect 49044 49861 49056 49895
rect 49090 49892 49102 49895
rect 50264 49892 50292 49932
rect 51997 49929 52009 49932
rect 52043 49929 52055 49963
rect 51997 49923 52055 49929
rect 54481 49963 54539 49969
rect 54481 49929 54493 49963
rect 54527 49960 54539 49963
rect 55398 49960 55404 49972
rect 54527 49932 55404 49960
rect 54527 49929 54539 49932
rect 54481 49923 54539 49929
rect 55398 49920 55404 49932
rect 55456 49920 55462 49972
rect 49090 49864 50292 49892
rect 50884 49895 50942 49901
rect 49090 49861 49102 49864
rect 49044 49855 49102 49861
rect 50884 49861 50896 49895
rect 50930 49892 50942 49895
rect 52086 49892 52092 49904
rect 50930 49864 52092 49892
rect 50930 49861 50942 49864
rect 50884 49855 50942 49861
rect 52086 49852 52092 49864
rect 52144 49852 52150 49904
rect 53116 49864 54984 49892
rect 1848 49827 1906 49833
rect 1848 49793 1860 49827
rect 1894 49824 1906 49827
rect 3510 49824 3516 49836
rect 1894 49796 3516 49824
rect 1894 49793 1906 49796
rect 1848 49787 1906 49793
rect 3510 49784 3516 49796
rect 3568 49784 3574 49836
rect 4700 49827 4758 49833
rect 4700 49793 4712 49827
rect 4746 49824 4758 49827
rect 6454 49824 6460 49836
rect 4746 49796 6460 49824
rect 4746 49793 4758 49796
rect 4700 49787 4758 49793
rect 6454 49784 6460 49796
rect 6512 49784 6518 49836
rect 9300 49827 9358 49833
rect 9300 49793 9312 49827
rect 9346 49824 9358 49827
rect 10226 49824 10232 49836
rect 9346 49796 10232 49824
rect 9346 49793 9358 49796
rect 9300 49787 9358 49793
rect 10226 49784 10232 49796
rect 10284 49784 10290 49836
rect 12897 49827 12955 49833
rect 12897 49793 12909 49827
rect 12943 49824 12955 49827
rect 13722 49824 13728 49836
rect 12943 49796 13728 49824
rect 12943 49793 12955 49796
rect 12897 49787 12955 49793
rect 13722 49784 13728 49796
rect 13780 49784 13786 49836
rect 13906 49784 13912 49836
rect 13964 49824 13970 49836
rect 14993 49827 15051 49833
rect 14993 49824 15005 49827
rect 13964 49796 15005 49824
rect 13964 49784 13970 49796
rect 14993 49793 15005 49796
rect 15039 49793 15051 49827
rect 14993 49787 15051 49793
rect 17037 49827 17095 49833
rect 17037 49793 17049 49827
rect 17083 49824 17095 49827
rect 19334 49824 19340 49836
rect 17083 49796 19340 49824
rect 17083 49793 17095 49796
rect 17037 49787 17095 49793
rect 19334 49784 19340 49796
rect 19392 49784 19398 49836
rect 19702 49824 19708 49836
rect 19615 49796 19708 49824
rect 19702 49784 19708 49796
rect 19760 49784 19766 49836
rect 19972 49827 20030 49833
rect 19972 49793 19984 49827
rect 20018 49824 20030 49827
rect 21082 49824 21088 49836
rect 20018 49796 21088 49824
rect 20018 49793 20030 49796
rect 19972 49787 20030 49793
rect 21082 49784 21088 49796
rect 21140 49784 21146 49836
rect 24854 49784 24860 49836
rect 24912 49824 24918 49836
rect 24949 49827 25007 49833
rect 24949 49824 24961 49827
rect 24912 49796 24961 49824
rect 24912 49784 24918 49796
rect 24949 49793 24961 49796
rect 24995 49793 25007 49827
rect 24949 49787 25007 49793
rect 25216 49827 25274 49833
rect 25216 49793 25228 49827
rect 25262 49824 25274 49827
rect 26418 49824 26424 49836
rect 25262 49796 26424 49824
rect 25262 49793 25274 49796
rect 25216 49787 25274 49793
rect 26418 49784 26424 49796
rect 26476 49784 26482 49836
rect 26970 49824 26976 49836
rect 26883 49796 26976 49824
rect 26970 49784 26976 49796
rect 27028 49824 27034 49836
rect 28813 49827 28871 49833
rect 28813 49824 28825 49827
rect 27028 49796 28825 49824
rect 27028 49784 27034 49796
rect 28813 49793 28825 49796
rect 28859 49824 28871 49827
rect 29546 49824 29552 49836
rect 28859 49796 29552 49824
rect 28859 49793 28871 49796
rect 28813 49787 28871 49793
rect 29546 49784 29552 49796
rect 29604 49784 29610 49836
rect 34698 49824 34704 49836
rect 34611 49796 34704 49824
rect 34698 49784 34704 49796
rect 34756 49824 34762 49836
rect 36538 49824 36544 49836
rect 34756 49796 36544 49824
rect 34756 49784 34762 49796
rect 36538 49784 36544 49796
rect 36596 49784 36602 49836
rect 37274 49824 37280 49836
rect 37187 49796 37280 49824
rect 37274 49784 37280 49796
rect 37332 49824 37338 49836
rect 39117 49827 39175 49833
rect 39117 49824 39129 49827
rect 37332 49796 39129 49824
rect 37332 49784 37338 49796
rect 39117 49793 39129 49796
rect 39163 49824 39175 49827
rect 48774 49824 48780 49836
rect 39163 49796 40163 49824
rect 48735 49796 48780 49824
rect 39163 49793 39175 49796
rect 39117 49787 39175 49793
rect 1578 49756 1584 49768
rect 1539 49728 1584 49756
rect 1578 49716 1584 49728
rect 1636 49716 1642 49768
rect 4433 49759 4491 49765
rect 4433 49725 4445 49759
rect 4479 49725 4491 49759
rect 6362 49756 6368 49768
rect 6323 49728 6368 49756
rect 4433 49719 4491 49725
rect 2958 49620 2964 49632
rect 2919 49592 2964 49620
rect 2958 49580 2964 49592
rect 3016 49580 3022 49632
rect 4448 49620 4476 49719
rect 6362 49716 6368 49728
rect 6420 49716 6426 49768
rect 8938 49716 8944 49768
rect 8996 49756 9002 49768
rect 9033 49759 9091 49765
rect 9033 49756 9045 49759
rect 8996 49728 9045 49756
rect 8996 49716 9002 49728
rect 9033 49725 9045 49728
rect 9079 49725 9091 49759
rect 14734 49756 14740 49768
rect 14695 49728 14740 49756
rect 9033 49719 9091 49725
rect 14734 49716 14740 49728
rect 14792 49716 14798 49768
rect 21726 49716 21732 49768
rect 21784 49756 21790 49768
rect 23109 49759 23167 49765
rect 23109 49756 23121 49759
rect 21784 49728 23121 49756
rect 21784 49716 21790 49728
rect 23109 49725 23121 49728
rect 23155 49725 23167 49759
rect 28718 49756 28724 49768
rect 23109 49719 23167 49725
rect 28368 49728 28724 49756
rect 5442 49648 5448 49700
rect 5500 49688 5506 49700
rect 6380 49688 6408 49716
rect 28368 49697 28396 49728
rect 28718 49716 28724 49728
rect 28776 49716 28782 49768
rect 35986 49716 35992 49768
rect 36044 49756 36050 49768
rect 38746 49756 38752 49768
rect 36044 49728 36124 49756
rect 36044 49716 36050 49728
rect 36096 49697 36124 49728
rect 38672 49728 38752 49756
rect 38672 49697 38700 49728
rect 38746 49716 38752 49728
rect 38804 49716 38810 49768
rect 5500 49660 6408 49688
rect 28353 49691 28411 49697
rect 5500 49648 5506 49660
rect 28353 49657 28365 49691
rect 28399 49657 28411 49691
rect 28353 49651 28411 49657
rect 36081 49691 36139 49697
rect 36081 49657 36093 49691
rect 36127 49657 36139 49691
rect 36081 49651 36139 49657
rect 38657 49691 38715 49697
rect 38657 49657 38669 49691
rect 38703 49657 38715 49691
rect 40135 49688 40163 49796
rect 48774 49784 48780 49796
rect 48832 49784 48838 49836
rect 45002 49716 45008 49768
rect 45060 49756 45066 49768
rect 45373 49759 45431 49765
rect 45373 49756 45385 49759
rect 45060 49728 45385 49756
rect 45060 49716 45066 49728
rect 45373 49725 45385 49728
rect 45419 49725 45431 49759
rect 50614 49756 50620 49768
rect 50575 49728 50620 49756
rect 45373 49719 45431 49725
rect 50614 49716 50620 49728
rect 50672 49716 50678 49768
rect 52730 49716 52736 49768
rect 52788 49756 52794 49768
rect 53116 49765 53144 49864
rect 53368 49827 53426 49833
rect 53368 49793 53380 49827
rect 53414 49824 53426 49827
rect 53926 49824 53932 49836
rect 53414 49796 53932 49824
rect 53414 49793 53426 49796
rect 53368 49787 53426 49793
rect 53926 49784 53932 49796
rect 53984 49784 53990 49836
rect 54956 49833 54984 49864
rect 54941 49827 54999 49833
rect 54941 49793 54953 49827
rect 54987 49793 54999 49827
rect 54941 49787 54999 49793
rect 55208 49827 55266 49833
rect 55208 49793 55220 49827
rect 55254 49824 55266 49827
rect 56778 49824 56784 49836
rect 55254 49796 56784 49824
rect 55254 49793 55266 49796
rect 55208 49787 55266 49793
rect 56778 49784 56784 49796
rect 56836 49784 56842 49836
rect 53101 49759 53159 49765
rect 53101 49756 53113 49759
rect 52788 49728 53113 49756
rect 52788 49716 52794 49728
rect 53101 49725 53113 49728
rect 53147 49725 53159 49759
rect 53101 49719 53159 49725
rect 40402 49688 40408 49700
rect 40135 49660 40408 49688
rect 38657 49651 38715 49657
rect 40402 49648 40408 49660
rect 40460 49648 40466 49700
rect 5460 49620 5488 49648
rect 5810 49620 5816 49632
rect 4448 49592 5488 49620
rect 5771 49592 5816 49620
rect 5810 49580 5816 49592
rect 5868 49580 5874 49632
rect 7742 49620 7748 49632
rect 7703 49592 7748 49620
rect 7742 49580 7748 49592
rect 7800 49580 7806 49632
rect 10410 49620 10416 49632
rect 10371 49592 10416 49620
rect 10410 49580 10416 49592
rect 10468 49580 10474 49632
rect 14277 49623 14335 49629
rect 14277 49589 14289 49623
rect 14323 49620 14335 49623
rect 14366 49620 14372 49632
rect 14323 49592 14372 49620
rect 14323 49589 14335 49592
rect 14277 49583 14335 49589
rect 14366 49580 14372 49592
rect 14424 49580 14430 49632
rect 40494 49620 40500 49632
rect 40455 49592 40500 49620
rect 40494 49580 40500 49592
rect 40552 49580 40558 49632
rect 46750 49620 46756 49632
rect 46711 49592 46756 49620
rect 46750 49580 46756 49592
rect 46808 49580 46814 49632
rect 50154 49620 50160 49632
rect 50115 49592 50160 49620
rect 50154 49580 50160 49592
rect 50212 49580 50218 49632
rect 56318 49620 56324 49632
rect 56279 49592 56324 49620
rect 56318 49580 56324 49592
rect 56376 49580 56382 49632
rect 1104 49530 59340 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 59340 49530
rect 1104 49456 59340 49478
rect 2866 49376 2872 49428
rect 2924 49416 2930 49428
rect 2961 49419 3019 49425
rect 2961 49416 2973 49419
rect 2924 49388 2973 49416
rect 2924 49376 2930 49388
rect 2961 49385 2973 49388
rect 3007 49385 3019 49419
rect 2961 49379 3019 49385
rect 6454 49376 6460 49428
rect 6512 49416 6518 49428
rect 6825 49419 6883 49425
rect 6825 49416 6837 49419
rect 6512 49388 6837 49416
rect 6512 49376 6518 49388
rect 6825 49385 6837 49388
rect 6871 49385 6883 49419
rect 6825 49379 6883 49385
rect 13541 49419 13599 49425
rect 13541 49385 13553 49419
rect 13587 49416 13599 49419
rect 13906 49416 13912 49428
rect 13587 49388 13912 49416
rect 13587 49385 13599 49388
rect 13541 49379 13599 49385
rect 13906 49376 13912 49388
rect 13964 49376 13970 49428
rect 14734 49416 14740 49428
rect 14108 49388 14740 49416
rect 13814 49308 13820 49360
rect 13872 49348 13878 49360
rect 14108 49348 14136 49388
rect 14734 49376 14740 49388
rect 14792 49376 14798 49428
rect 21082 49416 21088 49428
rect 21043 49388 21088 49416
rect 21082 49376 21088 49388
rect 21140 49376 21146 49428
rect 26418 49416 26424 49428
rect 26379 49388 26424 49416
rect 26418 49376 26424 49388
rect 26476 49376 26482 49428
rect 31294 49416 31300 49428
rect 31255 49388 31300 49416
rect 31294 49376 31300 49388
rect 31352 49376 31358 49428
rect 36538 49376 36544 49428
rect 36596 49416 36602 49428
rect 36817 49419 36875 49425
rect 36817 49416 36829 49419
rect 36596 49388 36829 49416
rect 36596 49376 36602 49388
rect 36817 49385 36829 49388
rect 36863 49385 36875 49419
rect 36817 49379 36875 49385
rect 41138 49376 41144 49428
rect 41196 49416 41202 49428
rect 41233 49419 41291 49425
rect 41233 49416 41245 49419
rect 41196 49388 41245 49416
rect 41196 49376 41202 49388
rect 41233 49385 41245 49388
rect 41279 49385 41291 49419
rect 41233 49379 41291 49385
rect 46290 49376 46296 49428
rect 46348 49416 46354 49428
rect 46385 49419 46443 49425
rect 46385 49416 46397 49419
rect 46348 49388 46397 49416
rect 46348 49376 46354 49388
rect 46385 49385 46397 49388
rect 46431 49385 46443 49419
rect 55950 49416 55956 49428
rect 46385 49379 46443 49385
rect 55324 49388 55956 49416
rect 13872 49320 14136 49348
rect 13872 49308 13878 49320
rect 4982 49240 4988 49292
rect 5040 49280 5046 49292
rect 5442 49280 5448 49292
rect 5040 49252 5448 49280
rect 5040 49240 5046 49252
rect 5442 49240 5448 49252
rect 5500 49240 5506 49292
rect 14108 49289 14136 49320
rect 55324 49292 55352 49388
rect 55950 49376 55956 49388
rect 56008 49416 56014 49428
rect 58526 49416 58532 49428
rect 56008 49388 57192 49416
rect 58487 49388 58532 49416
rect 56008 49376 56014 49388
rect 14093 49283 14151 49289
rect 14093 49249 14105 49283
rect 14139 49249 14151 49283
rect 14093 49243 14151 49249
rect 17034 49240 17040 49292
rect 17092 49280 17098 49292
rect 17221 49283 17279 49289
rect 17221 49280 17233 49283
rect 17092 49252 17233 49280
rect 17092 49240 17098 49252
rect 17221 49249 17233 49252
rect 17267 49249 17279 49283
rect 17221 49243 17279 49249
rect 19426 49240 19432 49292
rect 19484 49280 19490 49292
rect 19702 49280 19708 49292
rect 19484 49252 19708 49280
rect 19484 49240 19490 49252
rect 19702 49240 19708 49252
rect 19760 49240 19766 49292
rect 21726 49240 21732 49292
rect 21784 49280 21790 49292
rect 22465 49283 22523 49289
rect 22465 49280 22477 49283
rect 21784 49252 22477 49280
rect 21784 49240 21790 49252
rect 22465 49249 22477 49252
rect 22511 49249 22523 49283
rect 22465 49243 22523 49249
rect 24854 49240 24860 49292
rect 24912 49280 24918 49292
rect 25041 49283 25099 49289
rect 25041 49280 25053 49283
rect 24912 49252 25053 49280
rect 24912 49240 24918 49252
rect 25041 49249 25053 49252
rect 25087 49249 25099 49283
rect 25041 49243 25099 49249
rect 29546 49240 29552 49292
rect 29604 49280 29610 49292
rect 29917 49283 29975 49289
rect 29917 49280 29929 49283
rect 29604 49252 29929 49280
rect 29604 49240 29610 49252
rect 29917 49249 29929 49252
rect 29963 49249 29975 49283
rect 39850 49280 39856 49292
rect 39811 49252 39856 49280
rect 29917 49243 29975 49249
rect 39850 49240 39856 49252
rect 39908 49240 39914 49292
rect 48222 49280 48228 49292
rect 48135 49252 48228 49280
rect 48222 49240 48228 49252
rect 48280 49280 48286 49292
rect 55306 49280 55312 49292
rect 48280 49252 48360 49280
rect 55219 49252 55312 49280
rect 48280 49240 48286 49252
rect 1578 49212 1584 49224
rect 1491 49184 1584 49212
rect 1578 49172 1584 49184
rect 1636 49172 1642 49224
rect 1848 49215 1906 49221
rect 1848 49181 1860 49215
rect 1894 49212 1906 49215
rect 2958 49212 2964 49224
rect 1894 49184 2964 49212
rect 1894 49181 1906 49184
rect 1848 49175 1906 49181
rect 2958 49172 2964 49184
rect 3016 49172 3022 49224
rect 5712 49215 5770 49221
rect 5712 49181 5724 49215
rect 5758 49212 5770 49215
rect 7742 49212 7748 49224
rect 5758 49184 7748 49212
rect 5758 49181 5770 49184
rect 5712 49175 5770 49181
rect 7742 49172 7748 49184
rect 7800 49172 7806 49224
rect 8938 49212 8944 49224
rect 8899 49184 8944 49212
rect 8938 49172 8944 49184
rect 8996 49172 9002 49224
rect 12158 49212 12164 49224
rect 12119 49184 12164 49212
rect 12158 49172 12164 49184
rect 12216 49172 12222 49224
rect 13538 49212 13544 49224
rect 12268 49184 13544 49212
rect 1596 49144 1624 49172
rect 9208 49147 9266 49153
rect 1596 49116 1900 49144
rect 1872 49088 1900 49116
rect 9208 49113 9220 49147
rect 9254 49144 9266 49147
rect 12268 49144 12296 49184
rect 13538 49172 13544 49184
rect 13596 49172 13602 49224
rect 14366 49221 14372 49224
rect 14360 49212 14372 49221
rect 14327 49184 14372 49212
rect 14360 49175 14372 49184
rect 14366 49172 14372 49175
rect 14424 49172 14430 49224
rect 17488 49215 17546 49221
rect 17488 49181 17500 49215
rect 17534 49212 17546 49215
rect 17770 49212 17776 49224
rect 17534 49184 17776 49212
rect 17534 49181 17546 49184
rect 17488 49175 17546 49181
rect 17770 49172 17776 49184
rect 17828 49172 17834 49224
rect 31754 49212 31760 49224
rect 31715 49184 31760 49212
rect 31754 49172 31760 49184
rect 31812 49172 31818 49224
rect 32024 49215 32082 49221
rect 32024 49181 32036 49215
rect 32070 49212 32082 49215
rect 32766 49212 32772 49224
rect 32070 49184 32772 49212
rect 32070 49181 32082 49184
rect 32024 49175 32082 49181
rect 32766 49172 32772 49184
rect 32824 49172 32830 49224
rect 34790 49172 34796 49224
rect 34848 49212 34854 49224
rect 35529 49215 35587 49221
rect 35529 49212 35541 49215
rect 34848 49184 35541 49212
rect 34848 49172 34854 49184
rect 35529 49181 35541 49184
rect 35575 49212 35587 49215
rect 35575 49184 35894 49212
rect 35575 49181 35587 49184
rect 35529 49175 35587 49181
rect 9254 49116 12296 49144
rect 12428 49147 12486 49153
rect 9254 49113 9266 49116
rect 9208 49107 9266 49113
rect 12428 49113 12440 49147
rect 12474 49144 12486 49147
rect 19972 49147 20030 49153
rect 12474 49116 15516 49144
rect 12474 49113 12486 49116
rect 12428 49107 12486 49113
rect 1854 49036 1860 49088
rect 1912 49036 1918 49088
rect 10318 49076 10324 49088
rect 10279 49048 10324 49076
rect 10318 49036 10324 49048
rect 10376 49036 10382 49088
rect 15488 49085 15516 49116
rect 19972 49113 19984 49147
rect 20018 49144 20030 49147
rect 20990 49144 20996 49156
rect 20018 49116 20996 49144
rect 20018 49113 20030 49116
rect 19972 49107 20030 49113
rect 20990 49104 20996 49116
rect 21048 49104 21054 49156
rect 22732 49147 22790 49153
rect 22732 49113 22744 49147
rect 22778 49144 22790 49147
rect 24026 49144 24032 49156
rect 22778 49116 24032 49144
rect 22778 49113 22790 49116
rect 22732 49107 22790 49113
rect 24026 49104 24032 49116
rect 24084 49104 24090 49156
rect 25308 49147 25366 49153
rect 25308 49113 25320 49147
rect 25354 49144 25366 49147
rect 26326 49144 26332 49156
rect 25354 49116 26332 49144
rect 25354 49113 25366 49116
rect 25308 49107 25366 49113
rect 26326 49104 26332 49116
rect 26384 49104 26390 49156
rect 30184 49147 30242 49153
rect 30184 49113 30196 49147
rect 30230 49144 30242 49147
rect 30282 49144 30288 49156
rect 30230 49116 30288 49144
rect 30230 49113 30242 49116
rect 30184 49107 30242 49113
rect 30282 49104 30288 49116
rect 30340 49104 30346 49156
rect 15473 49079 15531 49085
rect 15473 49045 15485 49079
rect 15519 49045 15531 49079
rect 18598 49076 18604 49088
rect 18559 49048 18604 49076
rect 15473 49039 15531 49045
rect 18598 49036 18604 49048
rect 18656 49036 18662 49088
rect 23106 49036 23112 49088
rect 23164 49076 23170 49088
rect 23845 49079 23903 49085
rect 23845 49076 23857 49079
rect 23164 49048 23857 49076
rect 23164 49036 23170 49048
rect 23845 49045 23857 49048
rect 23891 49045 23903 49079
rect 33134 49076 33140 49088
rect 33095 49048 33140 49076
rect 23845 49039 23903 49045
rect 33134 49036 33140 49048
rect 33192 49036 33198 49088
rect 35866 49076 35894 49184
rect 39868 49144 39896 49240
rect 40120 49215 40178 49221
rect 40120 49181 40132 49215
rect 40166 49212 40178 49215
rect 40494 49212 40500 49224
rect 40166 49184 40500 49212
rect 40166 49181 40178 49184
rect 40120 49175 40178 49181
rect 40494 49172 40500 49184
rect 40552 49172 40558 49224
rect 41690 49212 41696 49224
rect 41603 49184 41696 49212
rect 41690 49172 41696 49184
rect 41748 49172 41754 49224
rect 45002 49212 45008 49224
rect 44963 49184 45008 49212
rect 45002 49172 45008 49184
rect 45060 49172 45066 49224
rect 45272 49215 45330 49221
rect 45272 49181 45284 49215
rect 45318 49212 45330 49215
rect 45646 49212 45652 49224
rect 45318 49184 45652 49212
rect 45318 49181 45330 49184
rect 45272 49175 45330 49181
rect 45646 49172 45652 49184
rect 45704 49172 45710 49224
rect 48332 49212 48360 49252
rect 55306 49240 55312 49252
rect 55364 49240 55370 49292
rect 57164 49289 57192 49388
rect 58526 49376 58532 49388
rect 58584 49376 58590 49428
rect 57149 49283 57207 49289
rect 57149 49249 57161 49283
rect 57195 49249 57207 49283
rect 57149 49243 57207 49249
rect 48492 49215 48550 49221
rect 48332 49184 48452 49212
rect 41708 49144 41736 49172
rect 39868 49116 41736 49144
rect 41782 49104 41788 49156
rect 41840 49144 41846 49156
rect 41938 49147 41996 49153
rect 41938 49144 41950 49147
rect 41840 49116 41950 49144
rect 41840 49104 41846 49116
rect 41938 49113 41950 49116
rect 41984 49113 41996 49147
rect 48424 49144 48452 49184
rect 48492 49181 48504 49215
rect 48538 49212 48550 49215
rect 50062 49212 50068 49224
rect 48538 49184 50068 49212
rect 48538 49181 48550 49184
rect 48492 49175 48550 49181
rect 50062 49172 50068 49184
rect 50120 49172 50126 49224
rect 50157 49215 50215 49221
rect 50157 49181 50169 49215
rect 50203 49212 50215 49215
rect 52730 49212 52736 49224
rect 50203 49184 50660 49212
rect 52691 49184 52736 49212
rect 50203 49181 50215 49184
rect 50157 49175 50215 49181
rect 50632 49156 50660 49184
rect 52730 49172 52736 49184
rect 52788 49172 52794 49224
rect 55576 49215 55634 49221
rect 55576 49181 55588 49215
rect 55622 49212 55634 49215
rect 56318 49212 56324 49224
rect 55622 49184 56324 49212
rect 55622 49181 55634 49184
rect 55576 49175 55634 49181
rect 56318 49172 56324 49184
rect 56376 49172 56382 49224
rect 57416 49215 57474 49221
rect 57416 49181 57428 49215
rect 57462 49212 57474 49215
rect 59449 49215 59507 49221
rect 59449 49212 59461 49215
rect 57462 49184 59461 49212
rect 57462 49181 57474 49184
rect 57416 49175 57474 49181
rect 59449 49181 59461 49184
rect 59495 49181 59507 49215
rect 59449 49175 59507 49181
rect 48774 49144 48780 49156
rect 48424 49116 48780 49144
rect 41938 49107 41996 49113
rect 48774 49104 48780 49116
rect 48832 49104 48838 49156
rect 50402 49147 50460 49153
rect 50402 49144 50414 49147
rect 49620 49116 50414 49144
rect 40310 49076 40316 49088
rect 35866 49048 40316 49076
rect 40310 49036 40316 49048
rect 40368 49036 40374 49088
rect 43070 49076 43076 49088
rect 43031 49048 43076 49076
rect 43070 49036 43076 49048
rect 43128 49036 43134 49088
rect 49620 49085 49648 49116
rect 50402 49113 50414 49116
rect 50448 49113 50460 49147
rect 50402 49107 50460 49113
rect 50614 49104 50620 49156
rect 50672 49104 50678 49156
rect 53000 49147 53058 49153
rect 53000 49113 53012 49147
rect 53046 49144 53058 49147
rect 53374 49144 53380 49156
rect 53046 49116 53380 49144
rect 53046 49113 53058 49116
rect 53000 49107 53058 49113
rect 53374 49104 53380 49116
rect 53432 49104 53438 49156
rect 49605 49079 49663 49085
rect 49605 49045 49617 49079
rect 49651 49045 49663 49079
rect 49605 49039 49663 49045
rect 49786 49036 49792 49088
rect 49844 49076 49850 49088
rect 51537 49079 51595 49085
rect 51537 49076 51549 49079
rect 49844 49048 51549 49076
rect 49844 49036 49850 49048
rect 51537 49045 51549 49048
rect 51583 49045 51595 49079
rect 51537 49039 51595 49045
rect 53834 49036 53840 49088
rect 53892 49076 53898 49088
rect 54113 49079 54171 49085
rect 54113 49076 54125 49079
rect 53892 49048 54125 49076
rect 53892 49036 53898 49048
rect 54113 49045 54125 49048
rect 54159 49045 54171 49079
rect 56686 49076 56692 49088
rect 56647 49048 56692 49076
rect 54113 49039 54171 49045
rect 56686 49036 56692 49048
rect 56744 49036 56750 49088
rect 1104 48986 59340 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 59340 48986
rect 1104 48912 59340 48934
rect 3510 48872 3516 48884
rect 3471 48844 3516 48872
rect 3510 48832 3516 48844
rect 3568 48832 3574 48884
rect 5353 48875 5411 48881
rect 5353 48872 5365 48875
rect 3896 48844 5365 48872
rect 2400 48807 2458 48813
rect 2400 48773 2412 48807
rect 2446 48804 2458 48807
rect 3896 48804 3924 48844
rect 5353 48841 5365 48844
rect 5399 48841 5411 48875
rect 5353 48835 5411 48841
rect 10226 48832 10232 48884
rect 10284 48872 10290 48884
rect 10413 48875 10471 48881
rect 10413 48872 10425 48875
rect 10284 48844 10425 48872
rect 10284 48832 10290 48844
rect 10413 48841 10425 48844
rect 10459 48841 10471 48875
rect 20990 48872 20996 48884
rect 20951 48844 20996 48872
rect 10413 48835 10471 48841
rect 20990 48832 20996 48844
rect 21048 48832 21054 48884
rect 26326 48832 26332 48884
rect 26384 48872 26390 48884
rect 26421 48875 26479 48881
rect 26421 48872 26433 48875
rect 26384 48844 26433 48872
rect 26384 48832 26390 48844
rect 26421 48841 26433 48844
rect 26467 48841 26479 48875
rect 41782 48872 41788 48884
rect 41743 48844 41788 48872
rect 26421 48835 26479 48841
rect 41782 48832 41788 48844
rect 41840 48832 41846 48884
rect 46382 48872 46388 48884
rect 46343 48844 46388 48872
rect 46382 48832 46388 48844
rect 46440 48832 46446 48884
rect 56778 48872 56784 48884
rect 56739 48844 56784 48872
rect 56778 48832 56784 48844
rect 56836 48832 56842 48884
rect 2446 48776 3924 48804
rect 4240 48807 4298 48813
rect 2446 48773 2458 48776
rect 2400 48767 2458 48773
rect 4240 48773 4252 48807
rect 4286 48804 4298 48807
rect 5810 48804 5816 48816
rect 4286 48776 5816 48804
rect 4286 48773 4298 48776
rect 4240 48767 4298 48773
rect 5810 48764 5816 48776
rect 5868 48764 5874 48816
rect 9300 48807 9358 48813
rect 9300 48773 9312 48807
rect 9346 48804 9358 48807
rect 10318 48804 10324 48816
rect 9346 48776 10324 48804
rect 9346 48773 9358 48776
rect 9300 48767 9358 48773
rect 10318 48764 10324 48776
rect 10376 48764 10382 48816
rect 12158 48804 12164 48816
rect 11716 48776 12164 48804
rect 2133 48739 2191 48745
rect 2133 48705 2145 48739
rect 2179 48736 2191 48739
rect 4982 48736 4988 48748
rect 2179 48708 4988 48736
rect 2179 48705 2191 48708
rect 2133 48699 2191 48705
rect 4982 48696 4988 48708
rect 5040 48696 5046 48748
rect 5534 48696 5540 48748
rect 5592 48736 5598 48748
rect 6825 48739 6883 48745
rect 6825 48736 6837 48739
rect 5592 48708 6837 48736
rect 5592 48696 5598 48708
rect 6825 48705 6837 48708
rect 6871 48705 6883 48739
rect 6825 48699 6883 48705
rect 3973 48671 4031 48677
rect 3973 48637 3985 48671
rect 4019 48637 4031 48671
rect 6840 48668 6868 48699
rect 8110 48696 8116 48748
rect 8168 48736 8174 48748
rect 11716 48745 11744 48776
rect 12158 48764 12164 48776
rect 12216 48804 12222 48816
rect 17212 48807 17270 48813
rect 12216 48776 13584 48804
rect 12216 48764 12222 48776
rect 8573 48739 8631 48745
rect 8573 48736 8585 48739
rect 8168 48708 8585 48736
rect 8168 48696 8174 48708
rect 8573 48705 8585 48708
rect 8619 48736 8631 48739
rect 9033 48739 9091 48745
rect 9033 48736 9045 48739
rect 8619 48708 9045 48736
rect 8619 48705 8631 48708
rect 8573 48699 8631 48705
rect 9033 48705 9045 48708
rect 9079 48705 9091 48739
rect 9033 48699 9091 48705
rect 11701 48739 11759 48745
rect 11701 48705 11713 48739
rect 11747 48705 11759 48739
rect 11701 48699 11759 48705
rect 11968 48739 12026 48745
rect 11968 48705 11980 48739
rect 12014 48736 12026 48739
rect 12894 48736 12900 48748
rect 12014 48708 12900 48736
rect 12014 48705 12026 48708
rect 11968 48699 12026 48705
rect 12894 48696 12900 48708
rect 12952 48696 12958 48748
rect 13556 48745 13584 48776
rect 17212 48773 17224 48807
rect 17258 48804 17270 48807
rect 18598 48804 18604 48816
rect 17258 48776 18604 48804
rect 17258 48773 17270 48776
rect 17212 48767 17270 48773
rect 18598 48764 18604 48776
rect 18656 48764 18662 48816
rect 32392 48807 32450 48813
rect 32392 48773 32404 48807
rect 32438 48804 32450 48807
rect 33134 48804 33140 48816
rect 32438 48776 33140 48804
rect 32438 48773 32450 48776
rect 32392 48767 32450 48773
rect 33134 48764 33140 48776
rect 33192 48764 33198 48816
rect 34330 48804 34336 48816
rect 33980 48776 34336 48804
rect 13541 48739 13599 48745
rect 13541 48705 13553 48739
rect 13587 48736 13599 48739
rect 13630 48736 13636 48748
rect 13587 48708 13636 48736
rect 13587 48705 13599 48708
rect 13541 48699 13599 48705
rect 13630 48696 13636 48708
rect 13688 48696 13694 48748
rect 13808 48739 13866 48745
rect 13808 48705 13820 48739
rect 13854 48736 13866 48739
rect 15470 48736 15476 48748
rect 13854 48708 15476 48736
rect 13854 48705 13866 48708
rect 13808 48699 13866 48705
rect 15470 48696 15476 48708
rect 15528 48696 15534 48748
rect 16945 48739 17003 48745
rect 16945 48705 16957 48739
rect 16991 48736 17003 48739
rect 17034 48736 17040 48748
rect 16991 48708 17040 48736
rect 16991 48705 17003 48708
rect 16945 48699 17003 48705
rect 17034 48696 17040 48708
rect 17092 48696 17098 48748
rect 19426 48696 19432 48748
rect 19484 48736 19490 48748
rect 19613 48739 19671 48745
rect 19613 48736 19625 48739
rect 19484 48708 19625 48736
rect 19484 48696 19490 48708
rect 19613 48705 19625 48708
rect 19659 48705 19671 48739
rect 19613 48699 19671 48705
rect 19880 48739 19938 48745
rect 19880 48705 19892 48739
rect 19926 48736 19938 48739
rect 20806 48736 20812 48748
rect 19926 48708 20812 48736
rect 19926 48705 19938 48708
rect 19880 48699 19938 48705
rect 20806 48696 20812 48708
rect 20864 48696 20870 48748
rect 22462 48736 22468 48748
rect 22423 48708 22468 48736
rect 22462 48696 22468 48708
rect 22520 48696 22526 48748
rect 22732 48739 22790 48745
rect 22732 48705 22744 48739
rect 22778 48736 22790 48739
rect 24394 48736 24400 48748
rect 22778 48708 24400 48736
rect 22778 48705 22790 48708
rect 22732 48699 22790 48705
rect 24394 48696 24400 48708
rect 24452 48696 24458 48748
rect 24854 48696 24860 48748
rect 24912 48736 24918 48748
rect 25041 48739 25099 48745
rect 25041 48736 25053 48739
rect 24912 48708 25053 48736
rect 24912 48696 24918 48708
rect 25041 48705 25053 48708
rect 25087 48705 25099 48739
rect 25041 48699 25099 48705
rect 25308 48739 25366 48745
rect 25308 48705 25320 48739
rect 25354 48736 25366 48739
rect 26418 48736 26424 48748
rect 25354 48708 26424 48736
rect 25354 48705 25366 48708
rect 25308 48699 25366 48705
rect 26418 48696 26424 48708
rect 26476 48696 26482 48748
rect 30460 48739 30518 48745
rect 30460 48705 30472 48739
rect 30506 48736 30518 48739
rect 32950 48736 32956 48748
rect 30506 48708 32956 48736
rect 30506 48705 30518 48708
rect 30460 48699 30518 48705
rect 32950 48696 32956 48708
rect 33008 48696 33014 48748
rect 33980 48745 34008 48776
rect 34330 48764 34336 48776
rect 34388 48764 34394 48816
rect 40672 48807 40730 48813
rect 40672 48773 40684 48807
rect 40718 48804 40730 48807
rect 41414 48804 41420 48816
rect 40718 48776 41420 48804
rect 40718 48773 40730 48776
rect 40672 48767 40730 48773
rect 41414 48764 41420 48776
rect 41472 48764 41478 48816
rect 43070 48764 43076 48816
rect 43128 48804 43134 48816
rect 43410 48807 43468 48813
rect 43410 48804 43422 48807
rect 43128 48776 43422 48804
rect 43128 48764 43134 48776
rect 43410 48773 43422 48776
rect 43456 48773 43468 48807
rect 43410 48767 43468 48773
rect 49044 48807 49102 48813
rect 49044 48773 49056 48807
rect 49090 48804 49102 48807
rect 50154 48804 50160 48816
rect 49090 48776 50160 48804
rect 49090 48773 49102 48776
rect 49044 48767 49102 48773
rect 50154 48764 50160 48776
rect 50212 48764 50218 48816
rect 55398 48764 55404 48816
rect 55456 48804 55462 48816
rect 55646 48807 55704 48813
rect 55646 48804 55658 48807
rect 55456 48776 55658 48804
rect 55456 48764 55462 48776
rect 55646 48773 55658 48776
rect 55692 48773 55704 48807
rect 55646 48767 55704 48773
rect 33965 48739 34023 48745
rect 33965 48705 33977 48739
rect 34011 48705 34023 48739
rect 33965 48699 34023 48705
rect 34232 48739 34290 48745
rect 34232 48705 34244 48739
rect 34278 48736 34290 48739
rect 35618 48736 35624 48748
rect 34278 48708 35624 48736
rect 34278 48705 34290 48708
rect 34232 48699 34290 48705
rect 35618 48696 35624 48708
rect 35676 48696 35682 48748
rect 37274 48736 37280 48748
rect 37235 48708 37280 48736
rect 37274 48696 37280 48708
rect 37332 48696 37338 48748
rect 37544 48739 37602 48745
rect 37544 48705 37556 48739
rect 37590 48736 37602 48739
rect 38746 48736 38752 48748
rect 37590 48708 38752 48736
rect 37590 48705 37602 48708
rect 37544 48699 37602 48705
rect 38746 48696 38752 48708
rect 38804 48696 38810 48748
rect 41690 48696 41696 48748
rect 41748 48736 41754 48748
rect 42426 48736 42432 48748
rect 41748 48708 42432 48736
rect 41748 48696 41754 48708
rect 42426 48696 42432 48708
rect 42484 48736 42490 48748
rect 43165 48739 43223 48745
rect 43165 48736 43177 48739
rect 42484 48708 43177 48736
rect 42484 48696 42490 48708
rect 43165 48705 43177 48708
rect 43211 48736 43223 48739
rect 43211 48708 44220 48736
rect 43211 48705 43223 48708
rect 43165 48699 43223 48705
rect 6840 48640 8984 48668
rect 3973 48631 4031 48637
rect 1854 48492 1860 48544
rect 1912 48532 1918 48544
rect 3988 48532 4016 48631
rect 1912 48504 4016 48532
rect 8956 48532 8984 48640
rect 30098 48628 30104 48680
rect 30156 48668 30162 48680
rect 30193 48671 30251 48677
rect 30193 48668 30205 48671
rect 30156 48640 30205 48668
rect 30156 48628 30162 48640
rect 30193 48637 30205 48640
rect 30239 48637 30251 48671
rect 31754 48668 31760 48680
rect 30193 48631 30251 48637
rect 31404 48640 31760 48668
rect 11882 48532 11888 48544
rect 8956 48504 11888 48532
rect 1912 48492 1918 48504
rect 11882 48492 11888 48504
rect 11940 48492 11946 48544
rect 13081 48535 13139 48541
rect 13081 48501 13093 48535
rect 13127 48532 13139 48535
rect 14182 48532 14188 48544
rect 13127 48504 14188 48532
rect 13127 48501 13139 48504
rect 13081 48495 13139 48501
rect 14182 48492 14188 48504
rect 14240 48492 14246 48544
rect 14918 48532 14924 48544
rect 14879 48504 14924 48532
rect 14918 48492 14924 48504
rect 14976 48492 14982 48544
rect 18322 48532 18328 48544
rect 18283 48504 18328 48532
rect 18322 48492 18328 48504
rect 18380 48492 18386 48544
rect 23842 48532 23848 48544
rect 23803 48504 23848 48532
rect 23842 48492 23848 48504
rect 23900 48492 23906 48544
rect 30208 48532 30236 48631
rect 31404 48532 31432 48640
rect 31754 48628 31760 48640
rect 31812 48668 31818 48680
rect 32125 48671 32183 48677
rect 32125 48668 32137 48671
rect 31812 48640 32137 48668
rect 31812 48628 31818 48640
rect 32125 48637 32137 48640
rect 32171 48637 32183 48671
rect 40402 48668 40408 48680
rect 40363 48640 40408 48668
rect 32125 48631 32183 48637
rect 40402 48628 40408 48640
rect 40460 48628 40466 48680
rect 44192 48668 44220 48708
rect 44450 48696 44456 48748
rect 44508 48736 44514 48748
rect 45261 48739 45319 48745
rect 45261 48736 45273 48739
rect 44508 48708 45273 48736
rect 44508 48696 44514 48708
rect 45261 48705 45273 48708
rect 45307 48705 45319 48739
rect 48774 48736 48780 48748
rect 48735 48708 48780 48736
rect 45261 48699 45319 48705
rect 48774 48696 48780 48708
rect 48832 48696 48838 48748
rect 53190 48736 53196 48748
rect 53151 48708 53196 48736
rect 53190 48696 53196 48708
rect 53248 48736 53254 48748
rect 56042 48736 56048 48748
rect 53248 48708 56048 48736
rect 53248 48696 53254 48708
rect 56042 48696 56048 48708
rect 56100 48696 56106 48748
rect 45002 48668 45008 48680
rect 44192 48640 45008 48668
rect 45002 48628 45008 48640
rect 45060 48628 45066 48680
rect 55306 48628 55312 48680
rect 55364 48668 55370 48680
rect 55401 48671 55459 48677
rect 55401 48668 55413 48671
rect 55364 48640 55413 48668
rect 55364 48628 55370 48640
rect 55401 48637 55413 48640
rect 55447 48637 55459 48671
rect 55401 48631 55459 48637
rect 50062 48560 50068 48612
rect 50120 48600 50126 48612
rect 50157 48603 50215 48609
rect 50157 48600 50169 48603
rect 50120 48572 50169 48600
rect 50120 48560 50126 48572
rect 50157 48569 50169 48572
rect 50203 48569 50215 48603
rect 50157 48563 50215 48569
rect 31570 48532 31576 48544
rect 30208 48504 31432 48532
rect 31531 48504 31576 48532
rect 31570 48492 31576 48504
rect 31628 48492 31634 48544
rect 33502 48532 33508 48544
rect 33463 48504 33508 48532
rect 33502 48492 33508 48504
rect 33560 48492 33566 48544
rect 34238 48492 34244 48544
rect 34296 48532 34302 48544
rect 35345 48535 35403 48541
rect 35345 48532 35357 48535
rect 34296 48504 35357 48532
rect 34296 48492 34302 48504
rect 35345 48501 35357 48504
rect 35391 48501 35403 48535
rect 35345 48495 35403 48501
rect 38010 48492 38016 48544
rect 38068 48532 38074 48544
rect 38657 48535 38715 48541
rect 38657 48532 38669 48535
rect 38068 48504 38669 48532
rect 38068 48492 38074 48504
rect 38657 48501 38669 48504
rect 38703 48501 38715 48535
rect 38657 48495 38715 48501
rect 42978 48492 42984 48544
rect 43036 48532 43042 48544
rect 44545 48535 44603 48541
rect 44545 48532 44557 48535
rect 43036 48504 44557 48532
rect 43036 48492 43042 48504
rect 44545 48501 44557 48504
rect 44591 48501 44603 48535
rect 44545 48495 44603 48501
rect 52730 48492 52736 48544
rect 52788 48532 52794 48544
rect 54481 48535 54539 48541
rect 54481 48532 54493 48535
rect 52788 48504 54493 48532
rect 52788 48492 52794 48504
rect 54481 48501 54493 48504
rect 54527 48501 54539 48535
rect 54481 48495 54539 48501
rect 1104 48442 59340 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 59340 48442
rect 1104 48368 59340 48390
rect 14826 48288 14832 48340
rect 14884 48328 14890 48340
rect 17034 48328 17040 48340
rect 14884 48300 17040 48328
rect 14884 48288 14890 48300
rect 17034 48288 17040 48300
rect 17092 48288 17098 48340
rect 22462 48288 22468 48340
rect 22520 48328 22526 48340
rect 22557 48331 22615 48337
rect 22557 48328 22569 48331
rect 22520 48300 22569 48328
rect 22520 48288 22526 48300
rect 22557 48297 22569 48300
rect 22603 48297 22615 48331
rect 22557 48291 22615 48297
rect 24854 48288 24860 48340
rect 24912 48328 24918 48340
rect 24912 48300 26234 48328
rect 24912 48288 24918 48300
rect 10778 48260 10784 48272
rect 10739 48232 10784 48260
rect 10778 48220 10784 48232
rect 10836 48220 10842 48272
rect 12894 48260 12900 48272
rect 12855 48232 12900 48260
rect 12894 48220 12900 48232
rect 12952 48220 12958 48272
rect 16022 48260 16028 48272
rect 15983 48232 16028 48260
rect 16022 48220 16028 48232
rect 16080 48220 16086 48272
rect 4982 48192 4988 48204
rect 4943 48164 4988 48192
rect 4982 48152 4988 48164
rect 5040 48152 5046 48204
rect 17052 48201 17080 48288
rect 20806 48260 20812 48272
rect 20767 48232 20812 48260
rect 20806 48220 20812 48232
rect 20864 48220 20870 48272
rect 26206 48260 26234 48300
rect 32950 48288 32956 48340
rect 33008 48328 33014 48340
rect 33008 48300 33180 48328
rect 33008 48288 33014 48300
rect 26973 48263 27031 48269
rect 26973 48260 26985 48263
rect 26206 48232 26985 48260
rect 26973 48229 26985 48232
rect 27019 48229 27031 48263
rect 33152 48260 33180 48300
rect 48222 48288 48228 48340
rect 48280 48328 48286 48340
rect 53374 48328 53380 48340
rect 48280 48300 49648 48328
rect 53335 48300 53380 48328
rect 48280 48288 48286 48300
rect 33597 48263 33655 48269
rect 33597 48260 33609 48263
rect 33152 48232 33609 48260
rect 26973 48223 27031 48229
rect 33597 48229 33609 48232
rect 33643 48229 33655 48263
rect 33597 48223 33655 48229
rect 43714 48220 43720 48272
rect 43772 48260 43778 48272
rect 43809 48263 43867 48269
rect 43809 48260 43821 48263
rect 43772 48232 43821 48260
rect 43772 48220 43778 48232
rect 43809 48229 43821 48232
rect 43855 48229 43867 48263
rect 49620 48260 49648 48300
rect 53374 48288 53380 48300
rect 53432 48288 53438 48340
rect 50062 48260 50068 48272
rect 49620 48232 50068 48260
rect 43809 48223 43867 48229
rect 50062 48220 50068 48232
rect 50120 48260 50126 48272
rect 50120 48232 50200 48260
rect 50120 48220 50126 48232
rect 17037 48195 17095 48201
rect 17037 48161 17049 48195
rect 17083 48161 17095 48195
rect 19426 48192 19432 48204
rect 19387 48164 19432 48192
rect 17037 48155 17095 48161
rect 19426 48152 19432 48164
rect 19484 48152 19490 48204
rect 36538 48192 36544 48204
rect 35866 48164 36544 48192
rect 8938 48084 8944 48136
rect 8996 48124 9002 48136
rect 9401 48127 9459 48133
rect 9401 48124 9413 48127
rect 8996 48096 9413 48124
rect 8996 48084 9002 48096
rect 9401 48093 9413 48096
rect 9447 48093 9459 48127
rect 9401 48087 9459 48093
rect 9668 48127 9726 48133
rect 9668 48093 9680 48127
rect 9714 48124 9726 48127
rect 10410 48124 10416 48136
rect 9714 48096 10416 48124
rect 9714 48093 9726 48096
rect 9668 48087 9726 48093
rect 5252 48059 5310 48065
rect 5252 48025 5264 48059
rect 5298 48056 5310 48059
rect 5902 48056 5908 48068
rect 5298 48028 5908 48056
rect 5298 48025 5310 48028
rect 5252 48019 5310 48025
rect 5902 48016 5908 48028
rect 5960 48016 5966 48068
rect 9416 48056 9444 48087
rect 10410 48084 10416 48096
rect 10468 48084 10474 48136
rect 11514 48124 11520 48136
rect 11475 48096 11520 48124
rect 11514 48084 11520 48096
rect 11572 48084 11578 48136
rect 14918 48133 14924 48136
rect 14645 48127 14703 48133
rect 14645 48093 14657 48127
rect 14691 48093 14703 48127
rect 14912 48124 14924 48133
rect 14879 48096 14924 48124
rect 14645 48087 14703 48093
rect 14912 48087 14924 48096
rect 11532 48056 11560 48084
rect 9416 48028 11560 48056
rect 11784 48059 11842 48065
rect 11784 48025 11796 48059
rect 11830 48056 11842 48059
rect 12894 48056 12900 48068
rect 11830 48028 12900 48056
rect 11830 48025 11842 48028
rect 11784 48019 11842 48025
rect 12894 48016 12900 48028
rect 12952 48016 12958 48068
rect 14660 48056 14688 48087
rect 14918 48084 14924 48087
rect 14976 48084 14982 48136
rect 17304 48127 17362 48133
rect 17304 48093 17316 48127
rect 17350 48124 17362 48127
rect 18322 48124 18328 48136
rect 17350 48096 18328 48124
rect 17350 48093 17362 48096
rect 17304 48087 17362 48093
rect 18322 48084 18328 48096
rect 18380 48084 18386 48136
rect 21174 48084 21180 48136
rect 21232 48124 21238 48136
rect 21269 48127 21327 48133
rect 21269 48124 21281 48127
rect 21232 48096 21281 48124
rect 21232 48084 21238 48096
rect 21269 48093 21281 48096
rect 21315 48124 21327 48127
rect 25685 48127 25743 48133
rect 25685 48124 25697 48127
rect 21315 48096 25697 48124
rect 21315 48093 21327 48096
rect 21269 48087 21327 48093
rect 25685 48093 25697 48096
rect 25731 48124 25743 48127
rect 25774 48124 25780 48136
rect 25731 48096 25780 48124
rect 25731 48093 25743 48096
rect 25685 48087 25743 48093
rect 25774 48084 25780 48096
rect 25832 48084 25838 48136
rect 30098 48084 30104 48136
rect 30156 48124 30162 48136
rect 30377 48127 30435 48133
rect 30377 48124 30389 48127
rect 30156 48096 30389 48124
rect 30156 48084 30162 48096
rect 30377 48093 30389 48096
rect 30423 48093 30435 48127
rect 30377 48087 30435 48093
rect 30644 48127 30702 48133
rect 30644 48093 30656 48127
rect 30690 48124 30702 48127
rect 31570 48124 31576 48136
rect 30690 48096 31576 48124
rect 30690 48093 30702 48096
rect 30644 48087 30702 48093
rect 31570 48084 31576 48096
rect 31628 48084 31634 48136
rect 32214 48124 32220 48136
rect 32175 48096 32220 48124
rect 32214 48084 32220 48096
rect 32272 48084 32278 48136
rect 32484 48127 32542 48133
rect 32484 48093 32496 48127
rect 32530 48124 32542 48127
rect 33502 48124 33508 48136
rect 32530 48096 33508 48124
rect 32530 48093 32542 48096
rect 32484 48087 32542 48093
rect 33502 48084 33508 48096
rect 33560 48084 33566 48136
rect 34330 48084 34336 48136
rect 34388 48124 34394 48136
rect 34701 48127 34759 48133
rect 34701 48124 34713 48127
rect 34388 48096 34713 48124
rect 34388 48084 34394 48096
rect 34701 48093 34713 48096
rect 34747 48124 34759 48127
rect 35866 48124 35894 48164
rect 36538 48152 36544 48164
rect 36596 48152 36602 48204
rect 42426 48192 42432 48204
rect 42387 48164 42432 48192
rect 42426 48152 42432 48164
rect 42484 48152 42490 48204
rect 45002 48152 45008 48204
rect 45060 48192 45066 48204
rect 45097 48195 45155 48201
rect 45097 48192 45109 48195
rect 45060 48164 45109 48192
rect 45060 48152 45066 48164
rect 45097 48161 45109 48164
rect 45143 48161 45155 48195
rect 48222 48192 48228 48204
rect 48183 48164 48228 48192
rect 45097 48155 45155 48161
rect 48222 48152 48228 48164
rect 48280 48152 48286 48204
rect 50172 48201 50200 48232
rect 56594 48220 56600 48272
rect 56652 48260 56658 48272
rect 56689 48263 56747 48269
rect 56689 48260 56701 48263
rect 56652 48232 56701 48260
rect 56652 48220 56658 48232
rect 56689 48229 56701 48232
rect 56735 48229 56747 48263
rect 56689 48223 56747 48229
rect 50157 48195 50215 48201
rect 50157 48161 50169 48195
rect 50203 48161 50215 48195
rect 50157 48155 50215 48161
rect 34747 48096 35894 48124
rect 39853 48127 39911 48133
rect 34747 48093 34759 48096
rect 34701 48087 34759 48093
rect 39853 48093 39865 48127
rect 39899 48124 39911 48127
rect 40402 48124 40408 48136
rect 39899 48096 40408 48124
rect 39899 48093 39911 48096
rect 39853 48087 39911 48093
rect 40402 48084 40408 48096
rect 40460 48084 40466 48136
rect 42696 48127 42754 48133
rect 42696 48093 42708 48127
rect 42742 48124 42754 48127
rect 42978 48124 42984 48136
rect 42742 48096 42984 48124
rect 42742 48093 42754 48096
rect 42696 48087 42754 48093
rect 42978 48084 42984 48096
rect 43036 48084 43042 48136
rect 48492 48127 48550 48133
rect 48492 48093 48504 48127
rect 48538 48124 48550 48127
rect 49786 48124 49792 48136
rect 48538 48096 49792 48124
rect 48538 48093 48550 48096
rect 48492 48087 48550 48093
rect 49786 48084 49792 48096
rect 49844 48084 49850 48136
rect 51997 48127 52055 48133
rect 51997 48093 52009 48127
rect 52043 48124 52055 48127
rect 52730 48124 52736 48136
rect 52043 48096 52736 48124
rect 52043 48093 52055 48096
rect 51997 48087 52055 48093
rect 52730 48084 52736 48096
rect 52788 48084 52794 48136
rect 55306 48124 55312 48136
rect 55267 48096 55312 48124
rect 55306 48084 55312 48096
rect 55364 48084 55370 48136
rect 55576 48127 55634 48133
rect 55576 48093 55588 48127
rect 55622 48124 55634 48127
rect 56686 48124 56692 48136
rect 55622 48096 56692 48124
rect 55622 48093 55634 48096
rect 55576 48087 55634 48093
rect 56686 48084 56692 48096
rect 56744 48084 56750 48136
rect 14826 48056 14832 48068
rect 14660 48028 14832 48056
rect 14826 48016 14832 48028
rect 14884 48016 14890 48068
rect 19696 48059 19754 48065
rect 19696 48025 19708 48059
rect 19742 48056 19754 48059
rect 20898 48056 20904 48068
rect 19742 48028 20904 48056
rect 19742 48025 19754 48028
rect 19696 48019 19754 48025
rect 20898 48016 20904 48028
rect 20956 48016 20962 48068
rect 34968 48059 35026 48065
rect 34968 48025 34980 48059
rect 35014 48056 35026 48059
rect 35986 48056 35992 48068
rect 35014 48028 35992 48056
rect 35014 48025 35026 48028
rect 34968 48019 35026 48025
rect 35986 48016 35992 48028
rect 36044 48016 36050 48068
rect 36786 48059 36844 48065
rect 36786 48056 36798 48059
rect 36096 48028 36798 48056
rect 6362 47988 6368 48000
rect 6323 47960 6368 47988
rect 6362 47948 6368 47960
rect 6420 47948 6426 48000
rect 18414 47988 18420 48000
rect 18375 47960 18420 47988
rect 18414 47948 18420 47960
rect 18472 47948 18478 48000
rect 31754 47988 31760 48000
rect 31715 47960 31760 47988
rect 31754 47948 31760 47960
rect 31812 47948 31818 48000
rect 36096 47997 36124 48028
rect 36786 48025 36798 48028
rect 36832 48025 36844 48059
rect 36786 48019 36844 48025
rect 40120 48059 40178 48065
rect 40120 48025 40132 48059
rect 40166 48056 40178 48059
rect 41138 48056 41144 48068
rect 40166 48028 41144 48056
rect 40166 48025 40178 48028
rect 40120 48019 40178 48025
rect 41138 48016 41144 48028
rect 41196 48016 41202 48068
rect 45364 48059 45422 48065
rect 45364 48025 45376 48059
rect 45410 48056 45422 48059
rect 46382 48056 46388 48068
rect 45410 48028 46388 48056
rect 45410 48025 45422 48028
rect 45364 48019 45422 48025
rect 46382 48016 46388 48028
rect 46440 48016 46446 48068
rect 49694 48016 49700 48068
rect 49752 48056 49758 48068
rect 50402 48059 50460 48065
rect 50402 48056 50414 48059
rect 49752 48028 50414 48056
rect 49752 48016 49758 48028
rect 50402 48025 50414 48028
rect 50448 48025 50460 48059
rect 50402 48019 50460 48025
rect 52264 48059 52322 48065
rect 52264 48025 52276 48059
rect 52310 48056 52322 48059
rect 54110 48056 54116 48068
rect 52310 48028 54116 48056
rect 52310 48025 52322 48028
rect 52264 48019 52322 48025
rect 54110 48016 54116 48028
rect 54168 48016 54174 48068
rect 36081 47991 36139 47997
rect 36081 47957 36093 47991
rect 36127 47957 36139 47991
rect 37918 47988 37924 48000
rect 37879 47960 37924 47988
rect 36081 47951 36139 47957
rect 37918 47948 37924 47960
rect 37976 47948 37982 48000
rect 41233 47991 41291 47997
rect 41233 47957 41245 47991
rect 41279 47988 41291 47991
rect 41782 47988 41788 48000
rect 41279 47960 41788 47988
rect 41279 47957 41291 47960
rect 41233 47951 41291 47957
rect 41782 47948 41788 47960
rect 41840 47948 41846 48000
rect 46477 47991 46535 47997
rect 46477 47957 46489 47991
rect 46523 47988 46535 47991
rect 47854 47988 47860 48000
rect 46523 47960 47860 47988
rect 46523 47957 46535 47960
rect 46477 47951 46535 47957
rect 47854 47948 47860 47960
rect 47912 47948 47918 48000
rect 49602 47988 49608 48000
rect 49563 47960 49608 47988
rect 49602 47948 49608 47960
rect 49660 47948 49666 48000
rect 50890 47948 50896 48000
rect 50948 47988 50954 48000
rect 51537 47991 51595 47997
rect 51537 47988 51549 47991
rect 50948 47960 51549 47988
rect 50948 47948 50954 47960
rect 51537 47957 51549 47960
rect 51583 47957 51595 47991
rect 51537 47951 51595 47957
rect 1104 47898 59340 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 59340 47898
rect 1104 47824 59340 47846
rect 15470 47784 15476 47796
rect 15431 47756 15476 47784
rect 15470 47744 15476 47756
rect 15528 47744 15534 47796
rect 20898 47784 20904 47796
rect 20859 47756 20904 47784
rect 20898 47744 20904 47756
rect 20956 47744 20962 47796
rect 24394 47784 24400 47796
rect 24355 47756 24400 47784
rect 24394 47744 24400 47756
rect 24452 47744 24458 47796
rect 26418 47784 26424 47796
rect 26379 47756 26424 47784
rect 26418 47744 26424 47756
rect 26476 47744 26482 47796
rect 35618 47784 35624 47796
rect 35579 47756 35624 47784
rect 35618 47744 35624 47756
rect 35676 47744 35682 47796
rect 44450 47784 44456 47796
rect 44411 47756 44456 47784
rect 44450 47744 44456 47756
rect 44508 47744 44514 47796
rect 50062 47784 50068 47796
rect 50023 47756 50068 47784
rect 50062 47744 50068 47756
rect 50120 47744 50126 47796
rect 54110 47784 54116 47796
rect 54071 47756 54116 47784
rect 54110 47744 54116 47756
rect 54168 47744 54174 47796
rect 4982 47716 4988 47728
rect 3528 47688 4988 47716
rect 3528 47657 3556 47688
rect 4982 47676 4988 47688
rect 5040 47676 5046 47728
rect 11882 47716 11888 47728
rect 11843 47688 11888 47716
rect 11882 47676 11888 47688
rect 11940 47676 11946 47728
rect 17212 47719 17270 47725
rect 17212 47685 17224 47719
rect 17258 47716 17270 47719
rect 18414 47716 18420 47728
rect 17258 47688 18420 47716
rect 17258 47685 17270 47688
rect 17212 47679 17270 47685
rect 18414 47676 18420 47688
rect 18472 47676 18478 47728
rect 23284 47719 23342 47725
rect 23284 47685 23296 47719
rect 23330 47716 23342 47719
rect 26234 47716 26240 47728
rect 23330 47688 26240 47716
rect 23330 47685 23342 47688
rect 23284 47679 23342 47685
rect 26234 47676 26240 47688
rect 26292 47676 26298 47728
rect 28896 47719 28954 47725
rect 28896 47685 28908 47719
rect 28942 47716 28954 47719
rect 28994 47716 29000 47728
rect 28942 47688 29000 47716
rect 28942 47685 28954 47688
rect 28896 47679 28954 47685
rect 28994 47676 29000 47688
rect 29052 47676 29058 47728
rect 31754 47676 31760 47728
rect 31812 47716 31818 47728
rect 32646 47719 32704 47725
rect 32646 47716 32658 47719
rect 31812 47688 32658 47716
rect 31812 47676 31818 47688
rect 32646 47685 32658 47688
rect 32692 47685 32704 47719
rect 32646 47679 32704 47685
rect 39669 47719 39727 47725
rect 39669 47685 39681 47719
rect 39715 47716 39727 47719
rect 40310 47716 40316 47728
rect 39715 47688 40316 47716
rect 39715 47685 39727 47688
rect 39669 47679 39727 47685
rect 40310 47676 40316 47688
rect 40368 47676 40374 47728
rect 43340 47719 43398 47725
rect 43340 47685 43352 47719
rect 43386 47716 43398 47719
rect 46750 47716 46756 47728
rect 43386 47688 46756 47716
rect 43386 47685 43398 47688
rect 43340 47679 43398 47685
rect 46750 47676 46756 47688
rect 46808 47676 46814 47728
rect 48777 47719 48835 47725
rect 48777 47685 48789 47719
rect 48823 47716 48835 47719
rect 53190 47716 53196 47728
rect 48823 47688 53196 47716
rect 48823 47685 48835 47688
rect 48777 47679 48835 47685
rect 53190 47676 53196 47688
rect 53248 47676 53254 47728
rect 3513 47651 3571 47657
rect 3513 47617 3525 47651
rect 3559 47617 3571 47651
rect 3513 47611 3571 47617
rect 3780 47651 3838 47657
rect 3780 47617 3792 47651
rect 3826 47648 3838 47651
rect 5166 47648 5172 47660
rect 3826 47620 5172 47648
rect 3826 47617 3838 47620
rect 3780 47611 3838 47617
rect 5166 47608 5172 47620
rect 5224 47608 5230 47660
rect 6632 47651 6690 47657
rect 6632 47617 6644 47651
rect 6678 47648 6690 47651
rect 7742 47648 7748 47660
rect 6678 47620 7748 47648
rect 6678 47617 6690 47620
rect 6632 47611 6690 47617
rect 7742 47608 7748 47620
rect 7800 47608 7806 47660
rect 14182 47608 14188 47660
rect 14240 47648 14246 47660
rect 14349 47651 14407 47657
rect 14349 47648 14361 47651
rect 14240 47620 14361 47648
rect 14240 47608 14246 47620
rect 14349 47617 14361 47620
rect 14395 47617 14407 47651
rect 14349 47611 14407 47617
rect 16945 47651 17003 47657
rect 16945 47617 16957 47651
rect 16991 47648 17003 47651
rect 17034 47648 17040 47660
rect 16991 47620 17040 47648
rect 16991 47617 17003 47620
rect 16945 47611 17003 47617
rect 17034 47608 17040 47620
rect 17092 47608 17098 47660
rect 19426 47608 19432 47660
rect 19484 47648 19490 47660
rect 19521 47651 19579 47657
rect 19521 47648 19533 47651
rect 19484 47620 19533 47648
rect 19484 47608 19490 47620
rect 19521 47617 19533 47620
rect 19567 47617 19579 47651
rect 19521 47611 19579 47617
rect 19788 47651 19846 47657
rect 19788 47617 19800 47651
rect 19834 47648 19846 47651
rect 20898 47648 20904 47660
rect 19834 47620 20904 47648
rect 19834 47617 19846 47620
rect 19788 47611 19846 47617
rect 20898 47608 20904 47620
rect 20956 47608 20962 47660
rect 22462 47608 22468 47660
rect 22520 47648 22526 47660
rect 23017 47651 23075 47657
rect 23017 47648 23029 47651
rect 22520 47620 23029 47648
rect 22520 47608 22526 47620
rect 23017 47617 23029 47620
rect 23063 47648 23075 47651
rect 24854 47648 24860 47660
rect 23063 47620 24860 47648
rect 23063 47617 23075 47620
rect 23017 47611 23075 47617
rect 24854 47608 24860 47620
rect 24912 47648 24918 47660
rect 25041 47651 25099 47657
rect 25041 47648 25053 47651
rect 24912 47620 25053 47648
rect 24912 47608 24918 47620
rect 25041 47617 25053 47620
rect 25087 47617 25099 47651
rect 25041 47611 25099 47617
rect 25308 47651 25366 47657
rect 25308 47617 25320 47651
rect 25354 47648 25366 47651
rect 26786 47648 26792 47660
rect 25354 47620 26792 47648
rect 25354 47617 25366 47620
rect 25308 47611 25366 47617
rect 26786 47608 26792 47620
rect 26844 47608 26850 47660
rect 32214 47608 32220 47660
rect 32272 47648 32278 47660
rect 32401 47651 32459 47657
rect 32401 47648 32413 47651
rect 32272 47620 32413 47648
rect 32272 47608 32278 47620
rect 32401 47617 32413 47620
rect 32447 47648 32459 47651
rect 34241 47651 34299 47657
rect 34241 47648 34253 47651
rect 32447 47620 34253 47648
rect 32447 47617 32459 47620
rect 32401 47611 32459 47617
rect 34241 47617 34253 47620
rect 34287 47648 34299 47651
rect 34330 47648 34336 47660
rect 34287 47620 34336 47648
rect 34287 47617 34299 47620
rect 34241 47611 34299 47617
rect 34330 47608 34336 47620
rect 34388 47608 34394 47660
rect 34514 47657 34520 47660
rect 34508 47611 34520 47657
rect 34572 47648 34578 47660
rect 34572 47620 34608 47648
rect 34514 47608 34520 47611
rect 34572 47608 34578 47620
rect 36538 47608 36544 47660
rect 36596 47648 36602 47660
rect 37277 47651 37335 47657
rect 37277 47648 37289 47651
rect 36596 47620 37289 47648
rect 36596 47608 36602 47620
rect 37277 47617 37289 47620
rect 37323 47617 37335 47651
rect 37277 47611 37335 47617
rect 37366 47608 37372 47660
rect 37424 47648 37430 47660
rect 37533 47651 37591 47657
rect 37533 47648 37545 47651
rect 37424 47620 37545 47648
rect 37424 47608 37430 47620
rect 37533 47617 37545 47620
rect 37579 47617 37591 47651
rect 37533 47611 37591 47617
rect 42426 47608 42432 47660
rect 42484 47648 42490 47660
rect 43073 47651 43131 47657
rect 43073 47648 43085 47651
rect 42484 47620 43085 47648
rect 42484 47608 42490 47620
rect 43073 47617 43085 47620
rect 43119 47648 43131 47651
rect 44913 47651 44971 47657
rect 44913 47648 44925 47651
rect 43119 47620 44925 47648
rect 43119 47617 43131 47620
rect 43073 47611 43131 47617
rect 44913 47617 44925 47620
rect 44959 47617 44971 47651
rect 44913 47611 44971 47617
rect 45180 47651 45238 47657
rect 45180 47617 45192 47651
rect 45226 47648 45238 47651
rect 45646 47648 45652 47660
rect 45226 47620 45652 47648
rect 45226 47617 45238 47620
rect 45180 47611 45238 47617
rect 45646 47608 45652 47620
rect 45704 47608 45710 47660
rect 52546 47608 52552 47660
rect 52604 47648 52610 47660
rect 52989 47651 53047 47657
rect 52989 47648 53001 47651
rect 52604 47620 53001 47648
rect 52604 47608 52610 47620
rect 52989 47617 53001 47620
rect 53035 47617 53047 47651
rect 52989 47611 53047 47617
rect 4982 47540 4988 47592
rect 5040 47580 5046 47592
rect 5442 47580 5448 47592
rect 5040 47552 5448 47580
rect 5040 47540 5046 47552
rect 5442 47540 5448 47552
rect 5500 47580 5506 47592
rect 6365 47583 6423 47589
rect 6365 47580 6377 47583
rect 5500 47552 6377 47580
rect 5500 47540 5506 47552
rect 6365 47549 6377 47552
rect 6411 47549 6423 47583
rect 13630 47580 13636 47592
rect 13591 47552 13636 47580
rect 6365 47543 6423 47549
rect 13630 47540 13636 47552
rect 13688 47540 13694 47592
rect 14093 47583 14151 47589
rect 14093 47549 14105 47583
rect 14139 47549 14151 47583
rect 14093 47543 14151 47549
rect 4893 47447 4951 47453
rect 4893 47413 4905 47447
rect 4939 47444 4951 47447
rect 5718 47444 5724 47456
rect 4939 47416 5724 47444
rect 4939 47413 4951 47416
rect 4893 47407 4951 47413
rect 5718 47404 5724 47416
rect 5776 47404 5782 47456
rect 7282 47404 7288 47456
rect 7340 47444 7346 47456
rect 7745 47447 7803 47453
rect 7745 47444 7757 47447
rect 7340 47416 7757 47444
rect 7340 47404 7346 47416
rect 7745 47413 7757 47416
rect 7791 47413 7803 47447
rect 14108 47444 14136 47543
rect 27614 47540 27620 47592
rect 27672 47580 27678 47592
rect 28629 47583 28687 47589
rect 28629 47580 28641 47583
rect 27672 47552 28641 47580
rect 27672 47540 27678 47552
rect 28629 47549 28641 47552
rect 28675 47549 28687 47583
rect 41322 47580 41328 47592
rect 41283 47552 41328 47580
rect 28629 47543 28687 47549
rect 41322 47540 41328 47552
rect 41380 47540 41386 47592
rect 52730 47580 52736 47592
rect 52691 47552 52736 47580
rect 52730 47540 52736 47552
rect 52788 47540 52794 47592
rect 14826 47444 14832 47456
rect 14108 47416 14832 47444
rect 7745 47407 7803 47413
rect 14826 47404 14832 47416
rect 14884 47404 14890 47456
rect 18322 47444 18328 47456
rect 18283 47416 18328 47444
rect 18322 47404 18328 47416
rect 18380 47404 18386 47456
rect 30006 47444 30012 47456
rect 29967 47416 30012 47444
rect 30006 47404 30012 47416
rect 30064 47404 30070 47456
rect 33778 47444 33784 47456
rect 33739 47416 33784 47444
rect 33778 47404 33784 47416
rect 33836 47404 33842 47456
rect 38654 47444 38660 47456
rect 38615 47416 38660 47444
rect 38654 47404 38660 47416
rect 38712 47404 38718 47456
rect 44542 47404 44548 47456
rect 44600 47444 44606 47456
rect 46293 47447 46351 47453
rect 46293 47444 46305 47447
rect 44600 47416 46305 47444
rect 44600 47404 44606 47416
rect 46293 47413 46305 47416
rect 46339 47413 46351 47447
rect 46293 47407 46351 47413
rect 1104 47354 59340 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 59340 47354
rect 1104 47280 59340 47302
rect 5166 47240 5172 47252
rect 5127 47212 5172 47240
rect 5166 47200 5172 47212
rect 5224 47200 5230 47252
rect 5810 47200 5816 47252
rect 5868 47240 5874 47252
rect 7009 47243 7067 47249
rect 7009 47240 7021 47243
rect 5868 47212 7021 47240
rect 5868 47200 5874 47212
rect 7009 47209 7021 47212
rect 7055 47209 7067 47243
rect 20898 47240 20904 47252
rect 20859 47212 20904 47240
rect 7009 47203 7067 47209
rect 20898 47200 20904 47212
rect 20956 47200 20962 47252
rect 26786 47240 26792 47252
rect 26747 47212 26792 47240
rect 26786 47200 26792 47212
rect 26844 47200 26850 47252
rect 35986 47200 35992 47252
rect 36044 47240 36050 47252
rect 36081 47243 36139 47249
rect 36081 47240 36093 47243
rect 36044 47212 36093 47240
rect 36044 47200 36050 47212
rect 36081 47209 36093 47212
rect 36127 47209 36139 47243
rect 46382 47240 46388 47252
rect 46343 47212 46388 47240
rect 36081 47203 36139 47209
rect 46382 47200 46388 47212
rect 46440 47200 46446 47252
rect 49605 47243 49663 47249
rect 49605 47209 49617 47243
rect 49651 47240 49663 47243
rect 49694 47240 49700 47252
rect 49651 47212 49700 47240
rect 49651 47209 49663 47212
rect 49605 47203 49663 47209
rect 49694 47200 49700 47212
rect 49752 47200 49758 47252
rect 53926 47240 53932 47252
rect 53887 47212 53932 47240
rect 53926 47200 53932 47212
rect 53984 47200 53990 47252
rect 28997 47175 29055 47181
rect 28997 47141 29009 47175
rect 29043 47172 29055 47175
rect 29178 47172 29184 47184
rect 29043 47144 29184 47172
rect 29043 47141 29055 47144
rect 28997 47135 29055 47141
rect 29178 47132 29184 47144
rect 29236 47132 29242 47184
rect 5442 47064 5448 47116
rect 5500 47104 5506 47116
rect 5629 47107 5687 47113
rect 5629 47104 5641 47107
rect 5500 47076 5641 47104
rect 5500 47064 5506 47076
rect 5629 47073 5641 47076
rect 5675 47073 5687 47107
rect 5629 47067 5687 47073
rect 19426 47064 19432 47116
rect 19484 47104 19490 47116
rect 19521 47107 19579 47113
rect 19521 47104 19533 47107
rect 19484 47076 19533 47104
rect 19484 47064 19490 47076
rect 19521 47073 19533 47076
rect 19567 47073 19579 47107
rect 22462 47104 22468 47116
rect 22423 47076 22468 47104
rect 19521 47067 19579 47073
rect 22462 47064 22468 47076
rect 22520 47064 22526 47116
rect 24854 47064 24860 47116
rect 24912 47104 24918 47116
rect 25409 47107 25467 47113
rect 25409 47104 25421 47107
rect 24912 47076 25421 47104
rect 24912 47064 24918 47076
rect 25409 47073 25421 47076
rect 25455 47073 25467 47107
rect 27614 47104 27620 47116
rect 27575 47076 27620 47104
rect 25409 47067 25467 47073
rect 3789 47039 3847 47045
rect 3789 47005 3801 47039
rect 3835 47036 3847 47039
rect 4338 47036 4344 47048
rect 3835 47008 4344 47036
rect 3835 47005 3847 47008
rect 3789 46999 3847 47005
rect 4338 46996 4344 47008
rect 4396 46996 4402 47048
rect 5718 46996 5724 47048
rect 5776 47036 5782 47048
rect 5885 47039 5943 47045
rect 5885 47036 5897 47039
rect 5776 47008 5897 47036
rect 5776 46996 5782 47008
rect 5885 47005 5897 47008
rect 5931 47005 5943 47039
rect 5885 46999 5943 47005
rect 10597 47039 10655 47045
rect 10597 47005 10609 47039
rect 10643 47036 10655 47039
rect 11422 47036 11428 47048
rect 10643 47008 11428 47036
rect 10643 47005 10655 47008
rect 10597 46999 10655 47005
rect 11422 46996 11428 47008
rect 11480 46996 11486 47048
rect 14826 47036 14832 47048
rect 14787 47008 14832 47036
rect 14826 46996 14832 47008
rect 14884 46996 14890 47048
rect 16853 47039 16911 47045
rect 16853 47005 16865 47039
rect 16899 47036 16911 47039
rect 16942 47036 16948 47048
rect 16899 47008 16948 47036
rect 16899 47005 16911 47008
rect 16853 46999 16911 47005
rect 16942 46996 16948 47008
rect 17000 46996 17006 47048
rect 17120 47039 17178 47045
rect 17120 47005 17132 47039
rect 17166 47036 17178 47039
rect 18322 47036 18328 47048
rect 17166 47008 18328 47036
rect 17166 47005 17178 47008
rect 17120 46999 17178 47005
rect 18322 46996 18328 47008
rect 18380 46996 18386 47048
rect 22732 47039 22790 47045
rect 22732 47005 22744 47039
rect 22778 47036 22790 47039
rect 23842 47036 23848 47048
rect 22778 47008 23848 47036
rect 22778 47005 22790 47008
rect 22732 46999 22790 47005
rect 23842 46996 23848 47008
rect 23900 46996 23906 47048
rect 25424 47036 25452 47067
rect 27614 47064 27620 47076
rect 27672 47064 27678 47116
rect 48222 47104 48228 47116
rect 48183 47076 48228 47104
rect 48222 47064 48228 47076
rect 48280 47064 48286 47116
rect 27632 47036 27660 47064
rect 25424 47008 27660 47036
rect 27884 47039 27942 47045
rect 27884 47005 27896 47039
rect 27930 47036 27942 47039
rect 30006 47036 30012 47048
rect 27930 47008 30012 47036
rect 27930 47005 27942 47008
rect 27884 46999 27942 47005
rect 30006 46996 30012 47008
rect 30064 46996 30070 47048
rect 30098 46996 30104 47048
rect 30156 47036 30162 47048
rect 31113 47039 31171 47045
rect 31113 47036 31125 47039
rect 30156 47008 31125 47036
rect 30156 46996 30162 47008
rect 31113 47005 31125 47008
rect 31159 47005 31171 47039
rect 31113 46999 31171 47005
rect 31380 47039 31438 47045
rect 31380 47005 31392 47039
rect 31426 47036 31438 47039
rect 33778 47036 33784 47048
rect 31426 47008 33784 47036
rect 31426 47005 31438 47008
rect 31380 46999 31438 47005
rect 33778 46996 33784 47008
rect 33836 46996 33842 47048
rect 34422 46996 34428 47048
rect 34480 47036 34486 47048
rect 34701 47039 34759 47045
rect 34701 47036 34713 47039
rect 34480 47008 34713 47036
rect 34480 46996 34486 47008
rect 34701 47005 34713 47008
rect 34747 47005 34759 47039
rect 34701 46999 34759 47005
rect 36541 47039 36599 47045
rect 36541 47005 36553 47039
rect 36587 47005 36599 47039
rect 36541 46999 36599 47005
rect 36808 47039 36866 47045
rect 36808 47005 36820 47039
rect 36854 47036 36866 47039
rect 37918 47036 37924 47048
rect 36854 47008 37924 47036
rect 36854 47005 36866 47008
rect 36808 46999 36866 47005
rect 4056 46971 4114 46977
rect 4056 46937 4068 46971
rect 4102 46968 4114 46971
rect 5534 46968 5540 46980
rect 4102 46940 5540 46968
rect 4102 46937 4114 46940
rect 4056 46931 4114 46937
rect 5534 46928 5540 46940
rect 5592 46928 5598 46980
rect 10864 46971 10922 46977
rect 10864 46937 10876 46971
rect 10910 46968 10922 46971
rect 12158 46968 12164 46980
rect 10910 46940 12164 46968
rect 10910 46937 10922 46940
rect 10864 46931 10922 46937
rect 12158 46928 12164 46940
rect 12216 46928 12222 46980
rect 15096 46971 15154 46977
rect 15096 46937 15108 46971
rect 15142 46968 15154 46971
rect 17954 46968 17960 46980
rect 15142 46940 17960 46968
rect 15142 46937 15154 46940
rect 15096 46931 15154 46937
rect 17954 46928 17960 46940
rect 18012 46928 18018 46980
rect 19788 46971 19846 46977
rect 19788 46937 19800 46971
rect 19834 46968 19846 46971
rect 20990 46968 20996 46980
rect 19834 46940 20996 46968
rect 19834 46937 19846 46940
rect 19788 46931 19846 46937
rect 20990 46928 20996 46940
rect 21048 46928 21054 46980
rect 25676 46971 25734 46977
rect 25676 46937 25688 46971
rect 25722 46968 25734 46971
rect 26418 46968 26424 46980
rect 25722 46940 26424 46968
rect 25722 46937 25734 46940
rect 25676 46931 25734 46937
rect 26418 46928 26424 46940
rect 26476 46928 26482 46980
rect 34968 46971 35026 46977
rect 34968 46937 34980 46971
rect 35014 46968 35026 46971
rect 35342 46968 35348 46980
rect 35014 46940 35348 46968
rect 35014 46937 35026 46940
rect 34968 46931 35026 46937
rect 35342 46928 35348 46940
rect 35400 46928 35406 46980
rect 36556 46968 36584 46999
rect 37918 46996 37924 47008
rect 37976 46996 37982 47048
rect 39853 47039 39911 47045
rect 39853 47005 39865 47039
rect 39899 47036 39911 47039
rect 40402 47036 40408 47048
rect 39899 47008 40408 47036
rect 39899 47005 39911 47008
rect 39853 46999 39911 47005
rect 40402 46996 40408 47008
rect 40460 47036 40466 47048
rect 41322 47036 41328 47048
rect 40460 47008 41328 47036
rect 40460 46996 40466 47008
rect 41322 46996 41328 47008
rect 41380 47036 41386 47048
rect 41693 47039 41751 47045
rect 41693 47036 41705 47039
rect 41380 47008 41705 47036
rect 41380 46996 41386 47008
rect 41693 47005 41705 47008
rect 41739 47005 41751 47039
rect 41693 46999 41751 47005
rect 41782 46996 41788 47048
rect 41840 47036 41846 47048
rect 41949 47039 42007 47045
rect 41949 47036 41961 47039
rect 41840 47008 41961 47036
rect 41840 46996 41846 47008
rect 41949 47005 41961 47008
rect 41995 47005 42007 47039
rect 41949 46999 42007 47005
rect 45005 47039 45063 47045
rect 45005 47005 45017 47039
rect 45051 47036 45063 47039
rect 46934 47036 46940 47048
rect 45051 47008 46940 47036
rect 45051 47005 45063 47008
rect 45005 46999 45063 47005
rect 46934 46996 46940 47008
rect 46992 46996 46998 47048
rect 48492 47039 48550 47045
rect 48492 47005 48504 47039
rect 48538 47036 48550 47039
rect 49602 47036 49608 47048
rect 48538 47008 49608 47036
rect 48538 47005 48550 47008
rect 48492 46999 48550 47005
rect 49602 46996 49608 47008
rect 49660 46996 49666 47048
rect 50614 47036 50620 47048
rect 50527 47008 50620 47036
rect 50614 46996 50620 47008
rect 50672 46996 50678 47048
rect 50890 47045 50896 47048
rect 50884 47036 50896 47045
rect 50851 47008 50896 47036
rect 50884 46999 50896 47008
rect 50890 46996 50896 46999
rect 50948 46996 50954 47048
rect 52549 47039 52607 47045
rect 52549 47005 52561 47039
rect 52595 47005 52607 47039
rect 52549 46999 52607 47005
rect 52816 47039 52874 47045
rect 52816 47005 52828 47039
rect 52862 47036 52874 47039
rect 53834 47036 53840 47048
rect 52862 47008 53840 47036
rect 52862 47005 52874 47008
rect 52816 46999 52874 47005
rect 37458 46968 37464 46980
rect 36556 46940 37464 46968
rect 37458 46928 37464 46940
rect 37516 46928 37522 46980
rect 40126 46977 40132 46980
rect 40120 46931 40132 46977
rect 40184 46968 40190 46980
rect 45272 46971 45330 46977
rect 40184 46940 40220 46968
rect 40126 46928 40132 46931
rect 40184 46928 40190 46940
rect 45272 46937 45284 46971
rect 45318 46968 45330 46971
rect 46198 46968 46204 46980
rect 45318 46940 46204 46968
rect 45318 46937 45330 46940
rect 45272 46931 45330 46937
rect 46198 46928 46204 46940
rect 46256 46928 46262 46980
rect 50632 46968 50660 46996
rect 52454 46968 52460 46980
rect 50632 46940 52460 46968
rect 52454 46928 52460 46940
rect 52512 46968 52518 46980
rect 52564 46968 52592 46999
rect 53834 46996 53840 47008
rect 53892 46996 53898 47048
rect 52730 46968 52736 46980
rect 52512 46940 52736 46968
rect 52512 46928 52518 46940
rect 52730 46928 52736 46940
rect 52788 46968 52794 46980
rect 53650 46968 53656 46980
rect 52788 46940 53656 46968
rect 52788 46928 52794 46940
rect 53650 46928 53656 46940
rect 53708 46968 53714 46980
rect 55306 46968 55312 46980
rect 53708 46940 55312 46968
rect 53708 46928 53714 46940
rect 55306 46928 55312 46940
rect 55364 46928 55370 46980
rect 11974 46900 11980 46912
rect 11935 46872 11980 46900
rect 11974 46860 11980 46872
rect 12032 46860 12038 46912
rect 16206 46900 16212 46912
rect 16167 46872 16212 46900
rect 16206 46860 16212 46872
rect 16264 46860 16270 46912
rect 18230 46900 18236 46912
rect 18191 46872 18236 46900
rect 18230 46860 18236 46872
rect 18288 46860 18294 46912
rect 23842 46900 23848 46912
rect 23803 46872 23848 46900
rect 23842 46860 23848 46872
rect 23900 46860 23906 46912
rect 32490 46900 32496 46912
rect 32451 46872 32496 46900
rect 32490 46860 32496 46872
rect 32548 46860 32554 46912
rect 37274 46860 37280 46912
rect 37332 46900 37338 46912
rect 37921 46903 37979 46909
rect 37921 46900 37933 46903
rect 37332 46872 37933 46900
rect 37332 46860 37338 46872
rect 37921 46869 37933 46872
rect 37967 46869 37979 46903
rect 41230 46900 41236 46912
rect 41191 46872 41236 46900
rect 37921 46863 37979 46869
rect 41230 46860 41236 46872
rect 41288 46860 41294 46912
rect 43070 46900 43076 46912
rect 43031 46872 43076 46900
rect 43070 46860 43076 46872
rect 43128 46860 43134 46912
rect 51994 46900 52000 46912
rect 51955 46872 52000 46900
rect 51994 46860 52000 46872
rect 52052 46860 52058 46912
rect 1104 46810 59340 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 59340 46810
rect 1104 46736 59340 46758
rect 3789 46699 3847 46705
rect 3789 46665 3801 46699
rect 3835 46665 3847 46699
rect 3789 46659 3847 46665
rect 3804 46628 3832 46659
rect 5534 46656 5540 46708
rect 5592 46696 5598 46708
rect 5629 46699 5687 46705
rect 5629 46696 5641 46699
rect 5592 46668 5641 46696
rect 5592 46656 5598 46668
rect 5629 46665 5641 46668
rect 5675 46665 5687 46699
rect 7742 46696 7748 46708
rect 7703 46668 7748 46696
rect 5629 46659 5687 46665
rect 7742 46656 7748 46668
rect 7800 46656 7806 46708
rect 12894 46696 12900 46708
rect 12855 46668 12900 46696
rect 12894 46656 12900 46668
rect 12952 46656 12958 46708
rect 20990 46696 20996 46708
rect 20951 46668 20996 46696
rect 20990 46656 20996 46668
rect 21048 46656 21054 46708
rect 24026 46696 24032 46708
rect 23987 46668 24032 46696
rect 24026 46656 24032 46668
rect 24084 46656 24090 46708
rect 26418 46696 26424 46708
rect 26379 46668 26424 46696
rect 26418 46656 26424 46668
rect 26476 46656 26482 46708
rect 35342 46696 35348 46708
rect 35303 46668 35348 46696
rect 35342 46656 35348 46668
rect 35400 46656 35406 46708
rect 45646 46696 45652 46708
rect 45607 46668 45652 46696
rect 45646 46656 45652 46668
rect 45704 46656 45710 46708
rect 50614 46696 50620 46708
rect 50356 46668 50620 46696
rect 4494 46631 4552 46637
rect 4494 46628 4506 46631
rect 3804 46600 4506 46628
rect 4494 46597 4506 46600
rect 4540 46597 4552 46631
rect 4494 46591 4552 46597
rect 4614 46588 4620 46640
rect 4672 46588 4678 46640
rect 6362 46588 6368 46640
rect 6420 46628 6426 46640
rect 6610 46631 6668 46637
rect 6610 46628 6622 46631
rect 6420 46600 6622 46628
rect 6420 46588 6426 46600
rect 6610 46597 6622 46600
rect 6656 46597 6668 46631
rect 6610 46591 6668 46597
rect 11784 46631 11842 46637
rect 11784 46597 11796 46631
rect 11830 46628 11842 46631
rect 11974 46628 11980 46640
rect 11830 46600 11980 46628
rect 11830 46597 11842 46600
rect 11784 46591 11842 46597
rect 11974 46588 11980 46600
rect 12032 46588 12038 46640
rect 15004 46631 15062 46637
rect 15004 46597 15016 46631
rect 15050 46628 15062 46631
rect 16206 46628 16212 46640
rect 15050 46600 16212 46628
rect 15050 46597 15062 46600
rect 15004 46591 15062 46597
rect 16206 46588 16212 46600
rect 16264 46588 16270 46640
rect 17028 46631 17086 46637
rect 17028 46597 17040 46631
rect 17074 46628 17086 46631
rect 18230 46628 18236 46640
rect 17074 46600 18236 46628
rect 17074 46597 17086 46600
rect 17028 46591 17086 46597
rect 18230 46588 18236 46600
rect 18288 46588 18294 46640
rect 22916 46631 22974 46637
rect 22916 46597 22928 46631
rect 22962 46628 22974 46631
rect 23842 46628 23848 46640
rect 22962 46600 23848 46628
rect 22962 46597 22974 46600
rect 22916 46591 22974 46597
rect 23842 46588 23848 46600
rect 23900 46588 23906 46640
rect 32392 46631 32450 46637
rect 32392 46597 32404 46631
rect 32438 46628 32450 46631
rect 32490 46628 32496 46640
rect 32438 46600 32496 46628
rect 32438 46597 32450 46600
rect 32392 46591 32450 46597
rect 32490 46588 32496 46600
rect 32548 46588 32554 46640
rect 34238 46637 34244 46640
rect 34232 46628 34244 46637
rect 34199 46600 34244 46628
rect 34232 46591 34244 46600
rect 34238 46588 34244 46591
rect 34296 46588 34302 46640
rect 34422 46588 34428 46640
rect 34480 46588 34486 46640
rect 37544 46631 37602 46637
rect 37544 46597 37556 46631
rect 37590 46628 37602 46631
rect 38654 46628 38660 46640
rect 37590 46600 38660 46628
rect 37590 46597 37602 46600
rect 37544 46591 37602 46597
rect 38654 46588 38660 46600
rect 38712 46588 38718 46640
rect 39384 46631 39442 46637
rect 39384 46597 39396 46631
rect 39430 46628 39442 46631
rect 41230 46628 41236 46640
rect 39430 46600 41236 46628
rect 39430 46597 39442 46600
rect 39384 46591 39442 46597
rect 41230 46588 41236 46600
rect 41288 46588 41294 46640
rect 47854 46637 47860 46640
rect 47848 46628 47860 46637
rect 47815 46600 47860 46628
rect 47848 46591 47860 46600
rect 47854 46588 47860 46591
rect 47912 46588 47918 46640
rect 2676 46563 2734 46569
rect 2676 46529 2688 46563
rect 2722 46560 2734 46563
rect 3234 46560 3240 46572
rect 2722 46532 3240 46560
rect 2722 46529 2734 46532
rect 2676 46523 2734 46529
rect 3234 46520 3240 46532
rect 3292 46520 3298 46572
rect 4249 46563 4307 46569
rect 4249 46529 4261 46563
rect 4295 46560 4307 46563
rect 4338 46560 4344 46572
rect 4295 46532 4344 46560
rect 4295 46529 4307 46532
rect 4249 46523 4307 46529
rect 4338 46520 4344 46532
rect 4396 46560 4402 46572
rect 4632 46560 4660 46588
rect 4396 46532 5488 46560
rect 4396 46520 4402 46532
rect 5460 46504 5488 46532
rect 7834 46520 7840 46572
rect 7892 46560 7898 46572
rect 8461 46563 8519 46569
rect 8461 46560 8473 46563
rect 7892 46532 8473 46560
rect 7892 46520 7898 46532
rect 8461 46529 8473 46532
rect 8507 46529 8519 46563
rect 8461 46523 8519 46529
rect 13630 46520 13636 46572
rect 13688 46560 13694 46572
rect 14737 46563 14795 46569
rect 14737 46560 14749 46563
rect 13688 46532 14749 46560
rect 13688 46520 13694 46532
rect 14737 46529 14749 46532
rect 14783 46529 14795 46563
rect 14737 46523 14795 46529
rect 16761 46563 16819 46569
rect 16761 46529 16773 46563
rect 16807 46560 16819 46563
rect 19426 46560 19432 46572
rect 16807 46532 19432 46560
rect 16807 46529 16819 46532
rect 16761 46523 16819 46529
rect 19426 46520 19432 46532
rect 19484 46560 19490 46572
rect 19613 46563 19671 46569
rect 19613 46560 19625 46563
rect 19484 46532 19625 46560
rect 19484 46520 19490 46532
rect 19613 46529 19625 46532
rect 19659 46529 19671 46563
rect 19613 46523 19671 46529
rect 19880 46563 19938 46569
rect 19880 46529 19892 46563
rect 19926 46560 19938 46563
rect 21082 46560 21088 46572
rect 19926 46532 21088 46560
rect 19926 46529 19938 46532
rect 19880 46523 19938 46529
rect 21082 46520 21088 46532
rect 21140 46520 21146 46572
rect 22554 46520 22560 46572
rect 22612 46560 22618 46572
rect 22649 46563 22707 46569
rect 22649 46560 22661 46563
rect 22612 46532 22661 46560
rect 22612 46520 22618 46532
rect 22649 46529 22661 46532
rect 22695 46529 22707 46563
rect 22649 46523 22707 46529
rect 24854 46520 24860 46572
rect 24912 46560 24918 46572
rect 25041 46563 25099 46569
rect 25041 46560 25053 46563
rect 24912 46532 25053 46560
rect 24912 46520 24918 46532
rect 25041 46529 25053 46532
rect 25087 46529 25099 46563
rect 25041 46523 25099 46529
rect 25308 46563 25366 46569
rect 25308 46529 25320 46563
rect 25354 46560 25366 46563
rect 26234 46560 26240 46572
rect 25354 46532 26240 46560
rect 25354 46529 25366 46532
rect 25308 46523 25366 46529
rect 26234 46520 26240 46532
rect 26292 46520 26298 46572
rect 29086 46569 29092 46572
rect 29080 46523 29092 46569
rect 29144 46560 29150 46572
rect 32125 46563 32183 46569
rect 29144 46532 29180 46560
rect 29086 46520 29092 46523
rect 29144 46520 29150 46532
rect 32125 46529 32137 46563
rect 32171 46560 32183 46563
rect 33965 46563 34023 46569
rect 33965 46560 33977 46563
rect 32171 46532 33977 46560
rect 32171 46529 32183 46532
rect 32125 46523 32183 46529
rect 33965 46529 33977 46532
rect 34011 46560 34023 46563
rect 34440 46560 34468 46588
rect 34011 46532 34468 46560
rect 37277 46563 37335 46569
rect 34011 46529 34023 46532
rect 33965 46523 34023 46529
rect 37277 46529 37289 46563
rect 37323 46560 37335 46563
rect 39117 46563 39175 46569
rect 39117 46560 39129 46563
rect 37323 46532 39129 46560
rect 37323 46529 37335 46532
rect 37277 46523 37335 46529
rect 39117 46529 39129 46532
rect 39163 46560 39175 46563
rect 40402 46560 40408 46572
rect 39163 46532 40408 46560
rect 39163 46529 39175 46532
rect 39117 46523 39175 46529
rect 1854 46452 1860 46504
rect 1912 46492 1918 46504
rect 2409 46495 2467 46501
rect 2409 46492 2421 46495
rect 1912 46464 2421 46492
rect 1912 46452 1918 46464
rect 2409 46461 2421 46464
rect 2455 46461 2467 46495
rect 2409 46455 2467 46461
rect 5442 46452 5448 46504
rect 5500 46492 5506 46504
rect 6365 46495 6423 46501
rect 6365 46492 6377 46495
rect 5500 46464 6377 46492
rect 5500 46452 5506 46464
rect 6365 46461 6377 46464
rect 6411 46461 6423 46495
rect 6365 46455 6423 46461
rect 8205 46495 8263 46501
rect 8205 46461 8217 46495
rect 8251 46461 8263 46495
rect 11514 46492 11520 46504
rect 11475 46464 11520 46492
rect 8205 46455 8263 46461
rect 8220 46356 8248 46455
rect 11514 46452 11520 46464
rect 11572 46452 11578 46504
rect 28813 46495 28871 46501
rect 28813 46461 28825 46495
rect 28859 46461 28871 46495
rect 28813 46455 28871 46461
rect 8938 46356 8944 46368
rect 8220 46328 8944 46356
rect 8938 46316 8944 46328
rect 8996 46316 9002 46368
rect 9582 46356 9588 46368
rect 9543 46328 9588 46356
rect 9582 46316 9588 46328
rect 9640 46316 9646 46368
rect 16114 46356 16120 46368
rect 16075 46328 16120 46356
rect 16114 46316 16120 46328
rect 16172 46316 16178 46368
rect 18138 46356 18144 46368
rect 18099 46328 18144 46356
rect 18138 46316 18144 46328
rect 18196 46316 18202 46368
rect 28828 46356 28856 46455
rect 30006 46356 30012 46368
rect 28828 46328 30012 46356
rect 30006 46316 30012 46328
rect 30064 46316 30070 46368
rect 30190 46356 30196 46368
rect 30151 46328 30196 46356
rect 30190 46316 30196 46328
rect 30248 46316 30254 46368
rect 33502 46356 33508 46368
rect 33463 46328 33508 46356
rect 33502 46316 33508 46328
rect 33560 46316 33566 46368
rect 37292 46356 37320 46523
rect 40402 46520 40408 46532
rect 40460 46520 40466 46572
rect 42426 46560 42432 46572
rect 42387 46532 42432 46560
rect 42426 46520 42432 46532
rect 42484 46520 42490 46572
rect 42696 46563 42754 46569
rect 42696 46529 42708 46563
rect 42742 46560 42754 46563
rect 43806 46560 43812 46572
rect 42742 46532 43812 46560
rect 42742 46529 42754 46532
rect 42696 46523 42754 46529
rect 43806 46520 43812 46532
rect 43864 46520 43870 46572
rect 44174 46520 44180 46572
rect 44232 46560 44238 46572
rect 44525 46563 44583 46569
rect 44525 46560 44537 46563
rect 44232 46532 44537 46560
rect 44232 46520 44238 46532
rect 44525 46529 44537 46532
rect 44571 46529 44583 46563
rect 44525 46523 44583 46529
rect 46934 46520 46940 46572
rect 46992 46560 46998 46572
rect 47581 46563 47639 46569
rect 47581 46560 47593 46563
rect 46992 46532 47593 46560
rect 46992 46520 46998 46532
rect 47581 46529 47593 46532
rect 47627 46560 47639 46563
rect 48222 46560 48228 46572
rect 47627 46532 48228 46560
rect 47627 46529 47639 46532
rect 47581 46523 47639 46529
rect 48222 46520 48228 46532
rect 48280 46520 48286 46572
rect 50157 46563 50215 46569
rect 50157 46529 50169 46563
rect 50203 46560 50215 46563
rect 50356 46560 50384 46668
rect 50614 46656 50620 46668
rect 50672 46656 50678 46708
rect 50424 46631 50482 46637
rect 50424 46597 50436 46631
rect 50470 46628 50482 46631
rect 51994 46628 52000 46640
rect 50470 46600 52000 46628
rect 50470 46597 50482 46600
rect 50424 46591 50482 46597
rect 51994 46588 52000 46600
rect 52052 46588 52058 46640
rect 53650 46560 53656 46572
rect 50203 46532 50384 46560
rect 53611 46532 53656 46560
rect 50203 46529 50215 46532
rect 50157 46523 50215 46529
rect 53650 46520 53656 46532
rect 53708 46520 53714 46572
rect 53920 46563 53978 46569
rect 53920 46529 53932 46563
rect 53966 46560 53978 46563
rect 55490 46560 55496 46572
rect 53966 46532 55496 46560
rect 53966 46529 53978 46532
rect 53920 46523 53978 46529
rect 55490 46520 55496 46532
rect 55548 46520 55554 46572
rect 55852 46563 55910 46569
rect 55852 46529 55864 46563
rect 55898 46560 55910 46563
rect 56686 46560 56692 46572
rect 55898 46532 56692 46560
rect 55898 46529 55910 46532
rect 55852 46523 55910 46529
rect 56686 46520 56692 46532
rect 56744 46520 56750 46572
rect 44266 46492 44272 46504
rect 44227 46464 44272 46492
rect 44266 46452 44272 46464
rect 44324 46452 44330 46504
rect 55306 46452 55312 46504
rect 55364 46492 55370 46504
rect 55585 46495 55643 46501
rect 55585 46492 55597 46495
rect 55364 46464 55597 46492
rect 55364 46452 55370 46464
rect 55585 46461 55597 46464
rect 55631 46461 55643 46495
rect 55585 46455 55643 46461
rect 38657 46427 38715 46433
rect 38657 46393 38669 46427
rect 38703 46424 38715 46427
rect 38746 46424 38752 46436
rect 38703 46396 38752 46424
rect 38703 46393 38715 46396
rect 38657 46387 38715 46393
rect 38746 46384 38752 46396
rect 38804 46384 38810 46436
rect 37458 46356 37464 46368
rect 37292 46328 37464 46356
rect 37458 46316 37464 46328
rect 37516 46316 37522 46368
rect 40497 46359 40555 46365
rect 40497 46325 40509 46359
rect 40543 46356 40555 46359
rect 40678 46356 40684 46368
rect 40543 46328 40684 46356
rect 40543 46325 40555 46328
rect 40497 46319 40555 46325
rect 40678 46316 40684 46328
rect 40736 46316 40742 46368
rect 42794 46316 42800 46368
rect 42852 46356 42858 46368
rect 43809 46359 43867 46365
rect 43809 46356 43821 46359
rect 42852 46328 43821 46356
rect 42852 46316 42858 46328
rect 43809 46325 43821 46328
rect 43855 46325 43867 46359
rect 48958 46356 48964 46368
rect 48919 46328 48964 46356
rect 43809 46319 43867 46325
rect 48958 46316 48964 46328
rect 49016 46316 49022 46368
rect 51534 46356 51540 46368
rect 51495 46328 51540 46356
rect 51534 46316 51540 46328
rect 51592 46316 51598 46368
rect 55030 46356 55036 46368
rect 54991 46328 55036 46356
rect 55030 46316 55036 46328
rect 55088 46316 55094 46368
rect 56965 46359 57023 46365
rect 56965 46325 56977 46359
rect 57011 46356 57023 46359
rect 57238 46356 57244 46368
rect 57011 46328 57244 46356
rect 57011 46325 57023 46328
rect 56965 46319 57023 46325
rect 57238 46316 57244 46328
rect 57296 46316 57302 46368
rect 1104 46266 59340 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 59340 46266
rect 1104 46192 59340 46214
rect 3234 46152 3240 46164
rect 3195 46124 3240 46152
rect 3234 46112 3240 46124
rect 3292 46112 3298 46164
rect 5442 46112 5448 46164
rect 5500 46112 5506 46164
rect 5902 46152 5908 46164
rect 5863 46124 5908 46152
rect 5902 46112 5908 46124
rect 5960 46112 5966 46164
rect 7834 46152 7840 46164
rect 7795 46124 7840 46152
rect 7834 46112 7840 46124
rect 7892 46112 7898 46164
rect 12158 46152 12164 46164
rect 12119 46124 12164 46152
rect 12158 46112 12164 46124
rect 12216 46112 12222 46164
rect 16942 46152 16948 46164
rect 16684 46124 16948 46152
rect 5460 46084 5488 46112
rect 5460 46056 6500 46084
rect 1854 46016 1860 46028
rect 1815 45988 1860 46016
rect 1854 45976 1860 45988
rect 1912 45976 1918 46028
rect 4522 46016 4528 46028
rect 4483 45988 4528 46016
rect 4522 45976 4528 45988
rect 4580 45976 4586 46028
rect 6472 46025 6500 46056
rect 16684 46025 16712 46124
rect 16942 46112 16948 46124
rect 17000 46112 17006 46164
rect 21082 46152 21088 46164
rect 21043 46124 21088 46152
rect 21082 46112 21088 46124
rect 21140 46112 21146 46164
rect 23750 46112 23756 46164
rect 23808 46152 23814 46164
rect 23845 46155 23903 46161
rect 23845 46152 23857 46155
rect 23808 46124 23857 46152
rect 23808 46112 23814 46124
rect 23845 46121 23857 46124
rect 23891 46121 23903 46155
rect 23845 46115 23903 46121
rect 26234 46112 26240 46164
rect 26292 46152 26298 46164
rect 28994 46152 29000 46164
rect 26292 46124 26337 46152
rect 28955 46124 29000 46152
rect 26292 46112 26298 46124
rect 28994 46112 29000 46124
rect 29052 46112 29058 46164
rect 33505 46155 33563 46161
rect 33505 46121 33517 46155
rect 33551 46152 33563 46155
rect 34514 46152 34520 46164
rect 33551 46124 34520 46152
rect 33551 46121 33563 46124
rect 33505 46115 33563 46121
rect 34514 46112 34520 46124
rect 34572 46112 34578 46164
rect 37001 46155 37059 46161
rect 37001 46121 37013 46155
rect 37047 46152 37059 46155
rect 37366 46152 37372 46164
rect 37047 46124 37372 46152
rect 37047 46121 37059 46124
rect 37001 46115 37059 46121
rect 37366 46112 37372 46124
rect 37424 46112 37430 46164
rect 38841 46155 38899 46161
rect 38841 46121 38853 46155
rect 38887 46152 38899 46155
rect 40126 46152 40132 46164
rect 38887 46124 40132 46152
rect 38887 46121 38899 46124
rect 38841 46115 38899 46121
rect 40126 46112 40132 46124
rect 40184 46112 40190 46164
rect 43806 46152 43812 46164
rect 43767 46124 43812 46152
rect 43806 46112 43812 46124
rect 43864 46112 43870 46164
rect 46198 46112 46204 46164
rect 46256 46152 46262 46164
rect 46385 46155 46443 46161
rect 46385 46152 46397 46155
rect 46256 46124 46397 46152
rect 46256 46112 46262 46124
rect 46385 46121 46397 46124
rect 46431 46121 46443 46155
rect 46385 46115 46443 46121
rect 51905 46155 51963 46161
rect 51905 46121 51917 46155
rect 51951 46152 51963 46155
rect 52546 46152 52552 46164
rect 51951 46124 52552 46152
rect 51951 46121 51963 46124
rect 51905 46115 51963 46121
rect 52546 46112 52552 46124
rect 52604 46112 52610 46164
rect 56686 46152 56692 46164
rect 56647 46124 56692 46152
rect 56686 46112 56692 46124
rect 56744 46112 56750 46164
rect 6457 46019 6515 46025
rect 6457 45985 6469 46019
rect 6503 45985 6515 46019
rect 16669 46019 16727 46025
rect 16669 46016 16681 46019
rect 6457 45979 6515 45985
rect 16546 45988 16681 46016
rect 4792 45951 4850 45957
rect 4792 45917 4804 45951
rect 4838 45948 4850 45951
rect 5810 45948 5816 45960
rect 4838 45920 5816 45948
rect 4838 45917 4850 45920
rect 4792 45911 4850 45917
rect 5810 45908 5816 45920
rect 5868 45908 5874 45960
rect 6724 45951 6782 45957
rect 6724 45917 6736 45951
rect 6770 45948 6782 45951
rect 7282 45948 7288 45960
rect 6770 45920 7288 45948
rect 6770 45917 6782 45920
rect 6724 45911 6782 45917
rect 7282 45908 7288 45920
rect 7340 45908 7346 45960
rect 8938 45948 8944 45960
rect 8851 45920 8944 45948
rect 8938 45908 8944 45920
rect 8996 45948 9002 45960
rect 10781 45951 10839 45957
rect 10781 45948 10793 45951
rect 8996 45920 10793 45948
rect 8996 45908 9002 45920
rect 10781 45917 10793 45920
rect 10827 45948 10839 45951
rect 11514 45948 11520 45960
rect 10827 45920 11520 45948
rect 10827 45917 10839 45920
rect 10781 45911 10839 45917
rect 11514 45908 11520 45920
rect 11572 45908 11578 45960
rect 14369 45951 14427 45957
rect 14369 45917 14381 45951
rect 14415 45917 14427 45951
rect 14369 45911 14427 45917
rect 14636 45951 14694 45957
rect 14636 45917 14648 45951
rect 14682 45948 14694 45951
rect 16114 45948 16120 45960
rect 14682 45920 16120 45948
rect 14682 45917 14694 45920
rect 14636 45911 14694 45917
rect 2124 45883 2182 45889
rect 2124 45849 2136 45883
rect 2170 45880 2182 45883
rect 4614 45880 4620 45892
rect 2170 45852 4620 45880
rect 2170 45849 2182 45852
rect 2124 45843 2182 45849
rect 4614 45840 4620 45852
rect 4672 45840 4678 45892
rect 8570 45840 8576 45892
rect 8628 45880 8634 45892
rect 9186 45883 9244 45889
rect 9186 45880 9198 45883
rect 8628 45852 9198 45880
rect 8628 45840 8634 45852
rect 9186 45849 9198 45852
rect 9232 45849 9244 45883
rect 9186 45843 9244 45849
rect 11048 45883 11106 45889
rect 11048 45849 11060 45883
rect 11094 45880 11106 45883
rect 12894 45880 12900 45892
rect 11094 45852 12900 45880
rect 11094 45849 11106 45852
rect 11048 45843 11106 45849
rect 12894 45840 12900 45852
rect 12952 45840 12958 45892
rect 14384 45880 14412 45911
rect 16114 45908 16120 45920
rect 16172 45908 16178 45960
rect 14826 45880 14832 45892
rect 14384 45852 14832 45880
rect 14826 45840 14832 45852
rect 14884 45880 14890 45892
rect 16546 45880 16574 45988
rect 16669 45985 16681 45988
rect 16715 45985 16727 46019
rect 16669 45979 16727 45985
rect 19426 45976 19432 46028
rect 19484 46016 19490 46028
rect 19705 46019 19763 46025
rect 19705 46016 19717 46019
rect 19484 45988 19717 46016
rect 19484 45976 19490 45988
rect 19705 45985 19717 45988
rect 19751 45985 19763 46019
rect 24854 46016 24860 46028
rect 24815 45988 24860 46016
rect 19705 45979 19763 45985
rect 24854 45976 24860 45988
rect 24912 45976 24918 46028
rect 27614 46016 27620 46028
rect 27575 45988 27620 46016
rect 27614 45976 27620 45988
rect 27672 45976 27678 46028
rect 30006 45976 30012 46028
rect 30064 46016 30070 46028
rect 30285 46019 30343 46025
rect 30285 46016 30297 46019
rect 30064 45988 30297 46016
rect 30064 45976 30070 45988
rect 30285 45985 30297 45988
rect 30331 45985 30343 46019
rect 30285 45979 30343 45985
rect 16936 45951 16994 45957
rect 16936 45917 16948 45951
rect 16982 45948 16994 45951
rect 18138 45948 18144 45960
rect 16982 45920 18144 45948
rect 16982 45917 16994 45920
rect 16936 45911 16994 45917
rect 18138 45908 18144 45920
rect 18196 45908 18202 45960
rect 22465 45951 22523 45957
rect 22465 45917 22477 45951
rect 22511 45948 22523 45951
rect 22554 45948 22560 45960
rect 22511 45920 22560 45948
rect 22511 45917 22523 45920
rect 22465 45911 22523 45917
rect 22554 45908 22560 45920
rect 22612 45908 22618 45960
rect 22732 45951 22790 45957
rect 22732 45917 22744 45951
rect 22778 45948 22790 45951
rect 23106 45948 23112 45960
rect 22778 45920 23112 45948
rect 22778 45917 22790 45920
rect 22732 45911 22790 45917
rect 23106 45908 23112 45920
rect 23164 45908 23170 45960
rect 27884 45951 27942 45957
rect 27884 45917 27896 45951
rect 27930 45948 27942 45951
rect 30190 45948 30196 45960
rect 27930 45920 30196 45948
rect 27930 45917 27942 45920
rect 27884 45911 27942 45917
rect 30190 45908 30196 45920
rect 30248 45908 30254 45960
rect 30300 45948 30328 45979
rect 34422 45976 34428 46028
rect 34480 46016 34486 46028
rect 35621 46019 35679 46025
rect 35621 46016 35633 46019
rect 34480 45988 35633 46016
rect 34480 45976 34486 45988
rect 35621 45985 35633 45988
rect 35667 45985 35679 46019
rect 37458 46016 37464 46028
rect 37419 45988 37464 46016
rect 35621 45979 35679 45985
rect 37458 45976 37464 45988
rect 37516 45976 37522 46028
rect 44266 45976 44272 46028
rect 44324 46016 44330 46028
rect 45005 46019 45063 46025
rect 45005 46016 45017 46019
rect 44324 45988 45017 46016
rect 44324 45976 44330 45988
rect 45005 45985 45017 45988
rect 45051 45985 45063 46019
rect 45005 45979 45063 45985
rect 32125 45951 32183 45957
rect 32125 45948 32137 45951
rect 30300 45920 32137 45948
rect 32125 45917 32137 45920
rect 32171 45917 32183 45951
rect 32125 45911 32183 45917
rect 32392 45951 32450 45957
rect 32392 45917 32404 45951
rect 32438 45948 32450 45951
rect 33502 45948 33508 45960
rect 32438 45920 33508 45948
rect 32438 45917 32450 45920
rect 32392 45911 32450 45917
rect 33502 45908 33508 45920
rect 33560 45908 33566 45960
rect 35888 45951 35946 45957
rect 35888 45917 35900 45951
rect 35934 45948 35946 45951
rect 37274 45948 37280 45960
rect 35934 45920 37280 45948
rect 35934 45917 35946 45920
rect 35888 45911 35946 45917
rect 37274 45908 37280 45920
rect 37332 45908 37338 45960
rect 37728 45951 37786 45957
rect 37728 45917 37740 45951
rect 37774 45948 37786 45951
rect 38010 45948 38016 45960
rect 37774 45920 38016 45948
rect 37774 45917 37786 45920
rect 37728 45911 37786 45917
rect 38010 45908 38016 45920
rect 38068 45908 38074 45960
rect 40586 45948 40592 45960
rect 40499 45920 40592 45948
rect 14884 45852 16574 45880
rect 19972 45883 20030 45889
rect 14884 45840 14890 45852
rect 19972 45849 19984 45883
rect 20018 45880 20030 45883
rect 21266 45880 21272 45892
rect 20018 45852 21272 45880
rect 20018 45849 20030 45852
rect 19972 45843 20030 45849
rect 21266 45840 21272 45852
rect 21324 45840 21330 45892
rect 24946 45840 24952 45892
rect 25004 45880 25010 45892
rect 25102 45883 25160 45889
rect 25102 45880 25114 45883
rect 25004 45852 25114 45880
rect 25004 45840 25010 45852
rect 25102 45849 25114 45852
rect 25148 45849 25160 45883
rect 25102 45843 25160 45849
rect 30552 45883 30610 45889
rect 30552 45849 30564 45883
rect 30598 45880 30610 45883
rect 31202 45880 31208 45892
rect 30598 45852 31208 45880
rect 30598 45849 30610 45852
rect 30552 45843 30610 45849
rect 31202 45840 31208 45852
rect 31260 45840 31266 45892
rect 40512 45880 40540 45920
rect 40586 45908 40592 45920
rect 40644 45908 40650 45960
rect 40678 45908 40684 45960
rect 40736 45948 40742 45960
rect 40845 45951 40903 45957
rect 40845 45948 40857 45951
rect 40736 45920 40857 45948
rect 40736 45908 40742 45920
rect 40845 45917 40857 45920
rect 40891 45917 40903 45951
rect 40845 45911 40903 45917
rect 41322 45908 41328 45960
rect 41380 45948 41386 45960
rect 42426 45948 42432 45960
rect 41380 45920 42432 45948
rect 41380 45908 41386 45920
rect 42426 45908 42432 45920
rect 42484 45908 42490 45960
rect 42696 45951 42754 45957
rect 42696 45917 42708 45951
rect 42742 45948 42754 45951
rect 43070 45948 43076 45960
rect 42742 45920 43076 45948
rect 42742 45917 42754 45920
rect 42696 45911 42754 45917
rect 43070 45908 43076 45920
rect 43128 45908 43134 45960
rect 45020 45948 45048 45979
rect 50062 45976 50068 46028
rect 50120 46016 50126 46028
rect 50525 46019 50583 46025
rect 50525 46016 50537 46019
rect 50120 45988 50537 46016
rect 50120 45976 50126 45988
rect 50525 45985 50537 45988
rect 50571 45985 50583 46019
rect 55306 46016 55312 46028
rect 55267 45988 55312 46016
rect 50525 45979 50583 45985
rect 55306 45976 55312 45988
rect 55364 45976 55370 46028
rect 45738 45948 45744 45960
rect 45020 45920 45744 45948
rect 45738 45908 45744 45920
rect 45796 45908 45802 45960
rect 46845 45951 46903 45957
rect 46845 45917 46857 45951
rect 46891 45948 46903 45951
rect 46934 45948 46940 45960
rect 46891 45920 46940 45948
rect 46891 45917 46903 45920
rect 46845 45911 46903 45917
rect 46934 45908 46940 45920
rect 46992 45908 46998 45960
rect 47112 45951 47170 45957
rect 47112 45917 47124 45951
rect 47158 45948 47170 45951
rect 48958 45948 48964 45960
rect 47158 45920 48964 45948
rect 47158 45917 47170 45920
rect 47112 45911 47170 45917
rect 48958 45908 48964 45920
rect 49016 45908 49022 45960
rect 50792 45951 50850 45957
rect 50792 45917 50804 45951
rect 50838 45948 50850 45951
rect 51534 45948 51540 45960
rect 50838 45920 51540 45948
rect 50838 45917 50850 45920
rect 50792 45911 50850 45917
rect 51534 45908 51540 45920
rect 51592 45908 51598 45960
rect 52365 45951 52423 45957
rect 52365 45917 52377 45951
rect 52411 45948 52423 45951
rect 52454 45948 52460 45960
rect 52411 45920 52460 45948
rect 52411 45917 52423 45920
rect 52365 45911 52423 45917
rect 52454 45908 52460 45920
rect 52512 45908 52518 45960
rect 41340 45880 41368 45908
rect 40512 45852 41368 45880
rect 45272 45883 45330 45889
rect 45272 45849 45284 45883
rect 45318 45880 45330 45883
rect 45646 45880 45652 45892
rect 45318 45852 45652 45880
rect 45318 45849 45330 45852
rect 45272 45843 45330 45849
rect 45646 45840 45652 45852
rect 45704 45840 45710 45892
rect 52632 45883 52690 45889
rect 52632 45849 52644 45883
rect 52678 45880 52690 45883
rect 53374 45880 53380 45892
rect 52678 45852 53380 45880
rect 52678 45849 52690 45852
rect 52632 45843 52690 45849
rect 53374 45840 53380 45852
rect 53432 45840 53438 45892
rect 55576 45883 55634 45889
rect 55576 45849 55588 45883
rect 55622 45880 55634 45883
rect 56686 45880 56692 45892
rect 55622 45852 56692 45880
rect 55622 45849 55634 45852
rect 55576 45843 55634 45849
rect 56686 45840 56692 45852
rect 56744 45840 56750 45892
rect 10318 45812 10324 45824
rect 10279 45784 10324 45812
rect 10318 45772 10324 45784
rect 10376 45772 10382 45824
rect 15746 45812 15752 45824
rect 15707 45784 15752 45812
rect 15746 45772 15752 45784
rect 15804 45772 15810 45824
rect 18046 45812 18052 45824
rect 18007 45784 18052 45812
rect 18046 45772 18052 45784
rect 18104 45772 18110 45824
rect 30282 45772 30288 45824
rect 30340 45812 30346 45824
rect 31665 45815 31723 45821
rect 31665 45812 31677 45815
rect 30340 45784 31677 45812
rect 30340 45772 30346 45784
rect 31665 45781 31677 45784
rect 31711 45781 31723 45815
rect 41966 45812 41972 45824
rect 41927 45784 41972 45812
rect 31665 45775 31723 45781
rect 41966 45772 41972 45784
rect 42024 45772 42030 45824
rect 48222 45812 48228 45824
rect 48183 45784 48228 45812
rect 48222 45772 48228 45784
rect 48280 45772 48286 45824
rect 53742 45812 53748 45824
rect 53703 45784 53748 45812
rect 53742 45772 53748 45784
rect 53800 45772 53806 45824
rect 1104 45722 59340 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 59340 45722
rect 1104 45648 59340 45670
rect 4614 45568 4620 45620
rect 4672 45608 4678 45620
rect 5077 45611 5135 45617
rect 5077 45608 5089 45611
rect 4672 45580 5089 45608
rect 4672 45568 4678 45580
rect 5077 45577 5089 45580
rect 5123 45577 5135 45611
rect 8570 45608 8576 45620
rect 8531 45580 8576 45608
rect 5077 45571 5135 45577
rect 8570 45568 8576 45580
rect 8628 45568 8634 45620
rect 12894 45608 12900 45620
rect 12855 45580 12900 45608
rect 12894 45568 12900 45580
rect 12952 45568 12958 45620
rect 21266 45608 21272 45620
rect 21227 45580 21272 45608
rect 21266 45568 21272 45580
rect 21324 45568 21330 45620
rect 45646 45608 45652 45620
rect 45607 45580 45652 45608
rect 45646 45568 45652 45580
rect 45704 45568 45710 45620
rect 55490 45568 55496 45620
rect 55548 45608 55554 45620
rect 55953 45611 56011 45617
rect 55953 45608 55965 45611
rect 55548 45580 55965 45608
rect 55548 45568 55554 45580
rect 55953 45577 55965 45580
rect 55999 45577 56011 45611
rect 55953 45571 56011 45577
rect 9300 45543 9358 45549
rect 9300 45509 9312 45543
rect 9346 45540 9358 45543
rect 10318 45540 10324 45552
rect 9346 45512 10324 45540
rect 9346 45509 9358 45512
rect 9300 45503 9358 45509
rect 10318 45500 10324 45512
rect 10376 45500 10382 45552
rect 13630 45540 13636 45552
rect 11532 45512 13636 45540
rect 11532 45484 11560 45512
rect 13630 45500 13636 45512
rect 13688 45540 13694 45552
rect 14360 45543 14418 45549
rect 13688 45512 14136 45540
rect 13688 45500 13694 45512
rect 2124 45475 2182 45481
rect 2124 45441 2136 45475
rect 2170 45472 2182 45475
rect 3142 45472 3148 45484
rect 2170 45444 3148 45472
rect 2170 45441 2182 45444
rect 2124 45435 2182 45441
rect 3142 45432 3148 45444
rect 3200 45432 3206 45484
rect 3953 45475 4011 45481
rect 3953 45472 3965 45475
rect 3252 45444 3965 45472
rect 1670 45364 1676 45416
rect 1728 45404 1734 45416
rect 1857 45407 1915 45413
rect 1857 45404 1869 45407
rect 1728 45376 1869 45404
rect 1728 45364 1734 45376
rect 1857 45373 1869 45376
rect 1903 45373 1915 45407
rect 1857 45367 1915 45373
rect 3252 45345 3280 45444
rect 3953 45441 3965 45444
rect 3999 45441 4011 45475
rect 3953 45435 4011 45441
rect 7460 45475 7518 45481
rect 7460 45441 7472 45475
rect 7506 45472 7518 45475
rect 9582 45472 9588 45484
rect 7506 45444 9588 45472
rect 7506 45441 7518 45444
rect 7460 45435 7518 45441
rect 9582 45432 9588 45444
rect 9640 45432 9646 45484
rect 11514 45472 11520 45484
rect 11475 45444 11520 45472
rect 11514 45432 11520 45444
rect 11572 45432 11578 45484
rect 11784 45475 11842 45481
rect 11784 45441 11796 45475
rect 11830 45472 11842 45475
rect 12894 45472 12900 45484
rect 11830 45444 12900 45472
rect 11830 45441 11842 45444
rect 11784 45435 11842 45441
rect 12894 45432 12900 45444
rect 12952 45432 12958 45484
rect 14108 45481 14136 45512
rect 14360 45509 14372 45543
rect 14406 45540 14418 45543
rect 15746 45540 15752 45552
rect 14406 45512 15752 45540
rect 14406 45509 14418 45512
rect 14360 45503 14418 45509
rect 15746 45500 15752 45512
rect 15804 45500 15810 45552
rect 16936 45543 16994 45549
rect 16936 45509 16948 45543
rect 16982 45540 16994 45543
rect 18046 45540 18052 45552
rect 16982 45512 18052 45540
rect 16982 45509 16994 45512
rect 16936 45503 16994 45509
rect 18046 45500 18052 45512
rect 18104 45500 18110 45552
rect 25038 45540 25044 45552
rect 21836 45512 25044 45540
rect 14093 45475 14151 45481
rect 14093 45441 14105 45475
rect 14139 45441 14151 45475
rect 19889 45475 19947 45481
rect 19889 45472 19901 45475
rect 14093 45435 14151 45441
rect 16684 45444 19901 45472
rect 16684 45416 16712 45444
rect 19889 45441 19901 45444
rect 19935 45472 19947 45475
rect 19978 45472 19984 45484
rect 19935 45444 19984 45472
rect 19935 45441 19947 45444
rect 19889 45435 19947 45441
rect 19978 45432 19984 45444
rect 20036 45432 20042 45484
rect 20156 45475 20214 45481
rect 20156 45441 20168 45475
rect 20202 45472 20214 45475
rect 21358 45472 21364 45484
rect 20202 45444 21364 45472
rect 20202 45441 20214 45444
rect 20156 45435 20214 45441
rect 21358 45432 21364 45444
rect 21416 45432 21422 45484
rect 21836 45416 21864 45512
rect 22088 45475 22146 45481
rect 22088 45441 22100 45475
rect 22134 45472 22146 45475
rect 23198 45472 23204 45484
rect 22134 45444 23204 45472
rect 22134 45441 22146 45444
rect 22088 45435 22146 45441
rect 23198 45432 23204 45444
rect 23256 45432 23262 45484
rect 24320 45481 24348 45512
rect 25038 45500 25044 45512
rect 25096 45500 25102 45552
rect 40586 45540 40592 45552
rect 33520 45512 35388 45540
rect 24305 45475 24363 45481
rect 24305 45441 24317 45475
rect 24351 45441 24363 45475
rect 24305 45435 24363 45441
rect 24572 45475 24630 45481
rect 24572 45441 24584 45475
rect 24618 45472 24630 45475
rect 25774 45472 25780 45484
rect 24618 45444 25780 45472
rect 24618 45441 24630 45444
rect 24572 45435 24630 45441
rect 25774 45432 25780 45444
rect 25832 45432 25838 45484
rect 28620 45475 28678 45481
rect 28620 45441 28632 45475
rect 28666 45472 28678 45475
rect 30098 45472 30104 45484
rect 28666 45444 30104 45472
rect 28666 45441 28678 45444
rect 28620 45435 28678 45441
rect 30098 45432 30104 45444
rect 30156 45432 30162 45484
rect 30460 45475 30518 45481
rect 30460 45441 30472 45475
rect 30506 45472 30518 45475
rect 31478 45472 31484 45484
rect 30506 45444 31484 45472
rect 30506 45441 30518 45444
rect 30460 45435 30518 45441
rect 31478 45432 31484 45444
rect 31536 45432 31542 45484
rect 3697 45407 3755 45413
rect 3697 45373 3709 45407
rect 3743 45373 3755 45407
rect 7190 45404 7196 45416
rect 7151 45376 7196 45404
rect 3697 45367 3755 45373
rect 3237 45339 3295 45345
rect 3237 45305 3249 45339
rect 3283 45305 3295 45339
rect 3237 45299 3295 45305
rect 3712 45268 3740 45367
rect 7190 45364 7196 45376
rect 7248 45364 7254 45416
rect 9030 45404 9036 45416
rect 8991 45376 9036 45404
rect 9030 45364 9036 45376
rect 9088 45364 9094 45416
rect 16666 45404 16672 45416
rect 16627 45376 16672 45404
rect 16666 45364 16672 45376
rect 16724 45364 16730 45416
rect 21818 45404 21824 45416
rect 21779 45376 21824 45404
rect 21818 45364 21824 45376
rect 21876 45364 21882 45416
rect 27706 45364 27712 45416
rect 27764 45404 27770 45416
rect 28353 45407 28411 45413
rect 28353 45404 28365 45407
rect 27764 45376 28365 45404
rect 27764 45364 27770 45376
rect 28353 45373 28365 45376
rect 28399 45373 28411 45407
rect 28353 45367 28411 45373
rect 30193 45407 30251 45413
rect 30193 45373 30205 45407
rect 30239 45373 30251 45407
rect 30193 45367 30251 45373
rect 17954 45296 17960 45348
rect 18012 45336 18018 45348
rect 18049 45339 18107 45345
rect 18049 45336 18061 45339
rect 18012 45308 18061 45336
rect 18012 45296 18018 45308
rect 18049 45305 18061 45308
rect 18095 45305 18107 45339
rect 18049 45299 18107 45305
rect 6362 45268 6368 45280
rect 3712 45240 6368 45268
rect 6362 45228 6368 45240
rect 6420 45268 6426 45280
rect 7190 45268 7196 45280
rect 6420 45240 7196 45268
rect 6420 45228 6426 45240
rect 7190 45228 7196 45240
rect 7248 45228 7254 45280
rect 10410 45268 10416 45280
rect 10371 45240 10416 45268
rect 10410 45228 10416 45240
rect 10468 45228 10474 45280
rect 15470 45268 15476 45280
rect 15431 45240 15476 45268
rect 15470 45228 15476 45240
rect 15528 45228 15534 45280
rect 20254 45228 20260 45280
rect 20312 45268 20318 45280
rect 23201 45271 23259 45277
rect 23201 45268 23213 45271
rect 20312 45240 23213 45268
rect 20312 45228 20318 45240
rect 23201 45237 23213 45240
rect 23247 45237 23259 45271
rect 25682 45268 25688 45280
rect 25643 45240 25688 45268
rect 23201 45231 23259 45237
rect 25682 45228 25688 45240
rect 25740 45228 25746 45280
rect 29730 45268 29736 45280
rect 29691 45240 29736 45268
rect 29730 45228 29736 45240
rect 29788 45228 29794 45280
rect 30208 45268 30236 45367
rect 31662 45364 31668 45416
rect 31720 45404 31726 45416
rect 33520 45413 33548 45512
rect 33772 45475 33830 45481
rect 33772 45441 33784 45475
rect 33818 45472 33830 45475
rect 34790 45472 34796 45484
rect 33818 45444 34796 45472
rect 33818 45441 33830 45444
rect 33772 45435 33830 45441
rect 34790 45432 34796 45444
rect 34848 45432 34854 45484
rect 35360 45481 35388 45512
rect 39868 45512 40592 45540
rect 35345 45475 35403 45481
rect 35345 45441 35357 45475
rect 35391 45441 35403 45475
rect 35345 45435 35403 45441
rect 35612 45475 35670 45481
rect 35612 45441 35624 45475
rect 35658 45472 35670 45475
rect 36538 45472 36544 45484
rect 35658 45444 36544 45472
rect 35658 45441 35670 45444
rect 35612 45435 35670 45441
rect 36538 45432 36544 45444
rect 36596 45432 36602 45484
rect 38280 45475 38338 45481
rect 38280 45441 38292 45475
rect 38326 45472 38338 45475
rect 39206 45472 39212 45484
rect 38326 45444 39212 45472
rect 38326 45441 38338 45444
rect 38280 45435 38338 45441
rect 39206 45432 39212 45444
rect 39264 45432 39270 45484
rect 39868 45481 39896 45512
rect 40586 45500 40592 45512
rect 40644 45500 40650 45552
rect 42696 45543 42754 45549
rect 42696 45509 42708 45543
rect 42742 45540 42754 45543
rect 42794 45540 42800 45552
rect 42742 45512 42800 45540
rect 42742 45509 42754 45512
rect 42696 45503 42754 45509
rect 42794 45500 42800 45512
rect 42852 45500 42858 45552
rect 44542 45549 44548 45552
rect 44536 45540 44548 45549
rect 44503 45512 44548 45540
rect 44536 45503 44548 45512
rect 44542 45500 44548 45503
rect 44600 45500 44606 45552
rect 47848 45543 47906 45549
rect 47848 45509 47860 45543
rect 47894 45540 47906 45543
rect 48222 45540 48228 45552
rect 47894 45512 48228 45540
rect 47894 45509 47906 45512
rect 47848 45503 47906 45509
rect 48222 45500 48228 45512
rect 48280 45500 48286 45552
rect 39853 45475 39911 45481
rect 39853 45441 39865 45475
rect 39899 45441 39911 45475
rect 39853 45435 39911 45441
rect 40120 45475 40178 45481
rect 40120 45441 40132 45475
rect 40166 45472 40178 45475
rect 41966 45472 41972 45484
rect 40166 45444 41972 45472
rect 40166 45441 40178 45444
rect 40120 45435 40178 45441
rect 41966 45432 41972 45444
rect 42024 45432 42030 45484
rect 42426 45472 42432 45484
rect 42387 45444 42432 45472
rect 42426 45432 42432 45444
rect 42484 45432 42490 45484
rect 42518 45432 42524 45484
rect 42576 45472 42582 45484
rect 44269 45475 44327 45481
rect 44269 45472 44281 45475
rect 42576 45444 44281 45472
rect 42576 45432 42582 45444
rect 44269 45441 44281 45444
rect 44315 45441 44327 45475
rect 44269 45435 44327 45441
rect 46934 45432 46940 45484
rect 46992 45472 46998 45484
rect 47578 45472 47584 45484
rect 46992 45444 47584 45472
rect 46992 45432 46998 45444
rect 47578 45432 47584 45444
rect 47636 45432 47642 45484
rect 50516 45475 50574 45481
rect 50516 45441 50528 45475
rect 50562 45472 50574 45475
rect 51534 45472 51540 45484
rect 50562 45444 51540 45472
rect 50562 45441 50574 45444
rect 50516 45435 50574 45441
rect 51534 45432 51540 45444
rect 51592 45432 51598 45484
rect 53000 45475 53058 45481
rect 53000 45441 53012 45475
rect 53046 45472 53058 45475
rect 54018 45472 54024 45484
rect 53046 45444 54024 45472
rect 53046 45441 53058 45444
rect 53000 45435 53058 45441
rect 54018 45432 54024 45444
rect 54076 45432 54082 45484
rect 54829 45475 54887 45481
rect 54829 45472 54841 45475
rect 54128 45444 54841 45472
rect 33505 45407 33563 45413
rect 33505 45404 33517 45407
rect 31720 45376 33517 45404
rect 31720 45364 31726 45376
rect 33505 45373 33517 45376
rect 33551 45373 33563 45407
rect 33505 45367 33563 45373
rect 37918 45364 37924 45416
rect 37976 45404 37982 45416
rect 38013 45407 38071 45413
rect 38013 45404 38025 45407
rect 37976 45376 38025 45404
rect 37976 45364 37982 45376
rect 38013 45373 38025 45376
rect 38059 45373 38071 45407
rect 38013 45367 38071 45373
rect 49418 45364 49424 45416
rect 49476 45404 49482 45416
rect 50249 45407 50307 45413
rect 50249 45404 50261 45407
rect 49476 45376 50261 45404
rect 49476 45364 49482 45376
rect 50249 45373 50261 45376
rect 50295 45373 50307 45407
rect 52730 45404 52736 45416
rect 52691 45376 52736 45404
rect 50249 45367 50307 45373
rect 52730 45364 52736 45376
rect 52788 45364 52794 45416
rect 41138 45296 41144 45348
rect 41196 45336 41202 45348
rect 41233 45339 41291 45345
rect 41233 45336 41245 45339
rect 41196 45308 41245 45336
rect 41196 45296 41202 45308
rect 41233 45305 41245 45308
rect 41279 45305 41291 45339
rect 41233 45299 41291 45305
rect 43809 45339 43867 45345
rect 43809 45305 43821 45339
rect 43855 45336 43867 45339
rect 44174 45336 44180 45348
rect 43855 45308 44180 45336
rect 43855 45305 43867 45308
rect 43809 45299 43867 45305
rect 44174 45296 44180 45308
rect 44232 45296 44238 45348
rect 54128 45345 54156 45444
rect 54829 45441 54841 45444
rect 54875 45441 54887 45475
rect 54829 45435 54887 45441
rect 54573 45407 54631 45413
rect 54573 45373 54585 45407
rect 54619 45373 54631 45407
rect 54573 45367 54631 45373
rect 54113 45339 54171 45345
rect 54113 45305 54125 45339
rect 54159 45305 54171 45339
rect 54113 45299 54171 45305
rect 30374 45268 30380 45280
rect 30208 45240 30380 45268
rect 30374 45228 30380 45240
rect 30432 45228 30438 45280
rect 31570 45268 31576 45280
rect 31531 45240 31576 45268
rect 31570 45228 31576 45240
rect 31628 45228 31634 45280
rect 33778 45228 33784 45280
rect 33836 45268 33842 45280
rect 34885 45271 34943 45277
rect 34885 45268 34897 45271
rect 33836 45240 34897 45268
rect 33836 45228 33842 45240
rect 34885 45237 34897 45240
rect 34931 45237 34943 45271
rect 34885 45231 34943 45237
rect 35342 45228 35348 45280
rect 35400 45268 35406 45280
rect 36725 45271 36783 45277
rect 36725 45268 36737 45271
rect 35400 45240 36737 45268
rect 35400 45228 35406 45240
rect 36725 45237 36737 45240
rect 36771 45237 36783 45271
rect 39390 45268 39396 45280
rect 39351 45240 39396 45268
rect 36725 45231 36783 45237
rect 39390 45228 39396 45240
rect 39448 45228 39454 45280
rect 48958 45268 48964 45280
rect 48919 45240 48964 45268
rect 48958 45228 48964 45240
rect 49016 45228 49022 45280
rect 51629 45271 51687 45277
rect 51629 45237 51641 45271
rect 51675 45268 51687 45271
rect 52086 45268 52092 45280
rect 51675 45240 52092 45268
rect 51675 45237 51687 45240
rect 51629 45231 51687 45237
rect 52086 45228 52092 45240
rect 52144 45228 52150 45280
rect 54588 45268 54616 45367
rect 56502 45268 56508 45280
rect 54588 45240 56508 45268
rect 56502 45228 56508 45240
rect 56560 45228 56566 45280
rect 1104 45178 59340 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 59340 45178
rect 1104 45104 59340 45126
rect 3142 45064 3148 45076
rect 3103 45036 3148 45064
rect 3142 45024 3148 45036
rect 3200 45024 3206 45076
rect 21358 45064 21364 45076
rect 21319 45036 21364 45064
rect 21358 45024 21364 45036
rect 21416 45024 21422 45076
rect 23198 45064 23204 45076
rect 23159 45036 23204 45064
rect 23198 45024 23204 45036
rect 23256 45024 23262 45076
rect 28997 45067 29055 45073
rect 28997 45033 29009 45067
rect 29043 45064 29055 45067
rect 29086 45064 29092 45076
rect 29043 45036 29092 45064
rect 29043 45033 29055 45036
rect 28997 45027 29055 45033
rect 29086 45024 29092 45036
rect 29144 45024 29150 45076
rect 31202 45024 31208 45076
rect 31260 45064 31266 45076
rect 31665 45067 31723 45073
rect 31665 45064 31677 45067
rect 31260 45036 31677 45064
rect 31260 45024 31266 45036
rect 31665 45033 31677 45036
rect 31711 45033 31723 45067
rect 51534 45064 51540 45076
rect 51495 45036 51540 45064
rect 31665 45027 31723 45033
rect 51534 45024 51540 45036
rect 51592 45024 51598 45076
rect 53374 45064 53380 45076
rect 53335 45036 53380 45064
rect 53374 45024 53380 45036
rect 53432 45024 53438 45076
rect 56686 45064 56692 45076
rect 56647 45036 56692 45064
rect 56686 45024 56692 45036
rect 56744 45024 56750 45076
rect 16666 44888 16672 44940
rect 16724 44928 16730 44940
rect 16853 44931 16911 44937
rect 16853 44928 16865 44931
rect 16724 44900 16865 44928
rect 16724 44888 16730 44900
rect 16853 44897 16865 44900
rect 16899 44897 16911 44931
rect 19978 44928 19984 44940
rect 19939 44900 19984 44928
rect 16853 44891 16911 44897
rect 19978 44888 19984 44900
rect 20036 44888 20042 44940
rect 45738 44928 45744 44940
rect 45699 44900 45744 44928
rect 45738 44888 45744 44900
rect 45796 44888 45802 44940
rect 47578 44928 47584 44940
rect 47539 44900 47584 44928
rect 47578 44888 47584 44900
rect 47636 44888 47642 44940
rect 56502 44888 56508 44940
rect 56560 44928 56566 44940
rect 57149 44931 57207 44937
rect 57149 44928 57161 44931
rect 56560 44900 57161 44928
rect 56560 44888 56566 44900
rect 57149 44897 57161 44900
rect 57195 44897 57207 44931
rect 57149 44891 57207 44897
rect 1670 44820 1676 44872
rect 1728 44860 1734 44872
rect 1765 44863 1823 44869
rect 1765 44860 1777 44863
rect 1728 44832 1777 44860
rect 1728 44820 1734 44832
rect 1765 44829 1777 44832
rect 1811 44829 1823 44863
rect 6362 44860 6368 44872
rect 6323 44832 6368 44860
rect 1765 44823 1823 44829
rect 6362 44820 6368 44832
rect 6420 44820 6426 44872
rect 8941 44863 8999 44869
rect 8941 44829 8953 44863
rect 8987 44860 8999 44863
rect 9030 44860 9036 44872
rect 8987 44832 9036 44860
rect 8987 44829 8999 44832
rect 8941 44823 8999 44829
rect 9030 44820 9036 44832
rect 9088 44860 9094 44872
rect 9490 44860 9496 44872
rect 9088 44832 9496 44860
rect 9088 44820 9094 44832
rect 9490 44820 9496 44832
rect 9548 44820 9554 44872
rect 10778 44860 10784 44872
rect 10739 44832 10784 44860
rect 10778 44820 10784 44832
rect 10836 44820 10842 44872
rect 14090 44860 14096 44872
rect 14051 44832 14096 44860
rect 14090 44820 14096 44832
rect 14148 44820 14154 44872
rect 14360 44863 14418 44869
rect 14360 44829 14372 44863
rect 14406 44860 14418 44863
rect 15470 44860 15476 44872
rect 14406 44832 15476 44860
rect 14406 44829 14418 44832
rect 14360 44823 14418 44829
rect 15470 44820 15476 44832
rect 15528 44820 15534 44872
rect 20254 44869 20260 44872
rect 20248 44860 20260 44869
rect 20215 44832 20260 44860
rect 20248 44823 20260 44832
rect 20254 44820 20260 44823
rect 20312 44820 20318 44872
rect 21542 44820 21548 44872
rect 21600 44860 21606 44872
rect 21821 44863 21879 44869
rect 21821 44860 21833 44863
rect 21600 44832 21833 44860
rect 21600 44820 21606 44832
rect 21821 44829 21833 44832
rect 21867 44829 21879 44863
rect 23014 44860 23020 44872
rect 21821 44823 21879 44829
rect 22020 44832 23020 44860
rect 2032 44795 2090 44801
rect 2032 44761 2044 44795
rect 2078 44792 2090 44795
rect 3050 44792 3056 44804
rect 2078 44764 3056 44792
rect 2078 44761 2090 44764
rect 2032 44755 2090 44761
rect 3050 44752 3056 44764
rect 3108 44752 3114 44804
rect 6632 44795 6690 44801
rect 6632 44761 6644 44795
rect 6678 44792 6690 44795
rect 7650 44792 7656 44804
rect 6678 44764 7656 44792
rect 6678 44761 6690 44764
rect 6632 44755 6690 44761
rect 7650 44752 7656 44764
rect 7708 44752 7714 44804
rect 9208 44795 9266 44801
rect 9208 44761 9220 44795
rect 9254 44792 9266 44795
rect 9582 44792 9588 44804
rect 9254 44764 9588 44792
rect 9254 44761 9266 44764
rect 9208 44755 9266 44761
rect 9582 44752 9588 44764
rect 9640 44752 9646 44804
rect 11026 44795 11084 44801
rect 11026 44792 11038 44795
rect 10336 44764 11038 44792
rect 7742 44724 7748 44736
rect 7703 44696 7748 44724
rect 7742 44684 7748 44696
rect 7800 44684 7806 44736
rect 10336 44733 10364 44764
rect 11026 44761 11038 44764
rect 11072 44761 11084 44795
rect 11026 44755 11084 44761
rect 17120 44795 17178 44801
rect 17120 44761 17132 44795
rect 17166 44792 17178 44795
rect 22020 44792 22048 44832
rect 23014 44820 23020 44832
rect 23072 44820 23078 44872
rect 25777 44863 25835 44869
rect 25777 44829 25789 44863
rect 25823 44860 25835 44863
rect 27617 44863 27675 44869
rect 27617 44860 27629 44863
rect 25823 44832 27629 44860
rect 25823 44829 25835 44832
rect 25777 44823 25835 44829
rect 27617 44829 27629 44832
rect 27663 44860 27675 44863
rect 27706 44860 27712 44872
rect 27663 44832 27712 44860
rect 27663 44829 27675 44832
rect 27617 44823 27675 44829
rect 27706 44820 27712 44832
rect 27764 44820 27770 44872
rect 27884 44863 27942 44869
rect 27884 44829 27896 44863
rect 27930 44860 27942 44863
rect 29730 44860 29736 44872
rect 27930 44832 29736 44860
rect 27930 44829 27942 44832
rect 27884 44823 27942 44829
rect 29730 44820 29736 44832
rect 29788 44820 29794 44872
rect 30285 44863 30343 44869
rect 30285 44829 30297 44863
rect 30331 44860 30343 44863
rect 30374 44860 30380 44872
rect 30331 44832 30380 44860
rect 30331 44829 30343 44832
rect 30285 44823 30343 44829
rect 30374 44820 30380 44832
rect 30432 44860 30438 44872
rect 31662 44860 31668 44872
rect 30432 44832 31668 44860
rect 30432 44820 30438 44832
rect 31662 44820 31668 44832
rect 31720 44860 31726 44872
rect 32125 44863 32183 44869
rect 32125 44860 32137 44863
rect 31720 44832 32137 44860
rect 31720 44820 31726 44832
rect 32125 44829 32137 44832
rect 32171 44829 32183 44863
rect 32125 44823 32183 44829
rect 36081 44863 36139 44869
rect 36081 44829 36093 44863
rect 36127 44860 36139 44863
rect 37918 44860 37924 44872
rect 36127 44832 37924 44860
rect 36127 44829 36139 44832
rect 36081 44823 36139 44829
rect 37918 44820 37924 44832
rect 37976 44820 37982 44872
rect 40402 44820 40408 44872
rect 40460 44860 40466 44872
rect 40589 44863 40647 44869
rect 40589 44860 40601 44863
rect 40460 44832 40601 44860
rect 40460 44820 40466 44832
rect 40589 44829 40601 44832
rect 40635 44860 40647 44863
rect 42426 44860 42432 44872
rect 40635 44832 42432 44860
rect 40635 44829 40647 44832
rect 40589 44823 40647 44829
rect 42426 44820 42432 44832
rect 42484 44820 42490 44872
rect 47848 44863 47906 44869
rect 47848 44829 47860 44863
rect 47894 44860 47906 44863
rect 48958 44860 48964 44872
rect 47894 44832 48964 44860
rect 47894 44829 47906 44832
rect 47848 44823 47906 44829
rect 48958 44820 48964 44832
rect 49016 44820 49022 44872
rect 50157 44863 50215 44869
rect 50157 44829 50169 44863
rect 50203 44860 50215 44863
rect 51997 44863 52055 44869
rect 51997 44860 52009 44863
rect 50203 44832 52009 44860
rect 50203 44829 50215 44832
rect 50157 44823 50215 44829
rect 51997 44829 52009 44832
rect 52043 44860 52055 44863
rect 52730 44860 52736 44872
rect 52043 44832 52736 44860
rect 52043 44829 52055 44832
rect 51997 44823 52055 44829
rect 52730 44820 52736 44832
rect 52788 44820 52794 44872
rect 54570 44820 54576 44872
rect 54628 44860 54634 44872
rect 55309 44863 55367 44869
rect 55309 44860 55321 44863
rect 54628 44832 55321 44860
rect 54628 44820 54634 44832
rect 55309 44829 55321 44832
rect 55355 44829 55367 44863
rect 55309 44823 55367 44829
rect 57238 44820 57244 44872
rect 57296 44860 57302 44872
rect 57405 44863 57463 44869
rect 57405 44860 57417 44863
rect 57296 44832 57417 44860
rect 57296 44820 57302 44832
rect 57405 44829 57417 44832
rect 57451 44829 57463 44863
rect 57405 44823 57463 44829
rect 17166 44764 22048 44792
rect 22088 44795 22146 44801
rect 17166 44761 17178 44764
rect 17120 44755 17178 44761
rect 22088 44761 22100 44795
rect 22134 44792 22146 44795
rect 23106 44792 23112 44804
rect 22134 44764 23112 44792
rect 22134 44761 22146 44764
rect 22088 44755 22146 44761
rect 23106 44752 23112 44764
rect 23164 44752 23170 44804
rect 26044 44795 26102 44801
rect 26044 44761 26056 44795
rect 26090 44792 26102 44795
rect 27522 44792 27528 44804
rect 26090 44764 27528 44792
rect 26090 44761 26102 44764
rect 26044 44755 26102 44761
rect 27522 44752 27528 44764
rect 27580 44752 27586 44804
rect 30552 44795 30610 44801
rect 30552 44761 30564 44795
rect 30598 44792 30610 44795
rect 32030 44792 32036 44804
rect 30598 44764 32036 44792
rect 30598 44761 30610 44764
rect 30552 44755 30610 44761
rect 32030 44752 32036 44764
rect 32088 44752 32094 44804
rect 32392 44795 32450 44801
rect 32392 44761 32404 44795
rect 32438 44792 32450 44795
rect 34054 44792 34060 44804
rect 32438 44764 34060 44792
rect 32438 44761 32450 44764
rect 32392 44755 32450 44761
rect 34054 44752 34060 44764
rect 34112 44752 34118 44804
rect 36348 44795 36406 44801
rect 36348 44761 36360 44795
rect 36394 44792 36406 44795
rect 38010 44792 38016 44804
rect 36394 44764 38016 44792
rect 36394 44761 36406 44764
rect 36348 44755 36406 44761
rect 38010 44752 38016 44764
rect 38068 44752 38074 44804
rect 38188 44795 38246 44801
rect 38188 44761 38200 44795
rect 38234 44792 38246 44795
rect 39114 44792 39120 44804
rect 38234 44764 39120 44792
rect 38234 44761 38246 44764
rect 38188 44755 38246 44761
rect 39114 44752 39120 44764
rect 39172 44752 39178 44804
rect 40856 44795 40914 44801
rect 40856 44761 40868 44795
rect 40902 44792 40914 44795
rect 41874 44792 41880 44804
rect 40902 44764 41880 44792
rect 40902 44761 40914 44764
rect 40856 44755 40914 44761
rect 41874 44752 41880 44764
rect 41932 44752 41938 44804
rect 42702 44801 42708 44804
rect 42696 44755 42708 44801
rect 42760 44792 42766 44804
rect 46008 44795 46066 44801
rect 42760 44764 42796 44792
rect 42702 44752 42708 44755
rect 42760 44752 42766 44764
rect 46008 44761 46020 44795
rect 46054 44792 46066 44795
rect 48866 44792 48872 44804
rect 46054 44764 48872 44792
rect 46054 44761 46066 44764
rect 46008 44755 46066 44761
rect 48866 44752 48872 44764
rect 48924 44752 48930 44804
rect 50424 44795 50482 44801
rect 50424 44761 50436 44795
rect 50470 44792 50482 44795
rect 51350 44792 51356 44804
rect 50470 44764 51356 44792
rect 50470 44761 50482 44764
rect 50424 44755 50482 44761
rect 51350 44752 51356 44764
rect 51408 44752 51414 44804
rect 52264 44795 52322 44801
rect 52264 44761 52276 44795
rect 52310 44792 52322 44795
rect 53374 44792 53380 44804
rect 52310 44764 53380 44792
rect 52310 44761 52322 44764
rect 52264 44755 52322 44761
rect 53374 44752 53380 44764
rect 53432 44752 53438 44804
rect 55576 44795 55634 44801
rect 55576 44761 55588 44795
rect 55622 44792 55634 44795
rect 55950 44792 55956 44804
rect 55622 44764 55956 44792
rect 55622 44761 55634 44764
rect 55576 44755 55634 44761
rect 55950 44752 55956 44764
rect 56008 44752 56014 44804
rect 10321 44727 10379 44733
rect 10321 44693 10333 44727
rect 10367 44693 10379 44727
rect 12158 44724 12164 44736
rect 12119 44696 12164 44724
rect 10321 44687 10379 44693
rect 12158 44684 12164 44696
rect 12216 44684 12222 44736
rect 15470 44724 15476 44736
rect 15431 44696 15476 44724
rect 15470 44684 15476 44696
rect 15528 44684 15534 44736
rect 18230 44724 18236 44736
rect 18191 44696 18236 44724
rect 18230 44684 18236 44696
rect 18288 44684 18294 44736
rect 27154 44724 27160 44736
rect 27115 44696 27160 44724
rect 27154 44684 27160 44696
rect 27212 44684 27218 44736
rect 31938 44684 31944 44736
rect 31996 44724 32002 44736
rect 33505 44727 33563 44733
rect 33505 44724 33517 44727
rect 31996 44696 33517 44724
rect 31996 44684 32002 44696
rect 33505 44693 33517 44696
rect 33551 44693 33563 44727
rect 33505 44687 33563 44693
rect 36722 44684 36728 44736
rect 36780 44724 36786 44736
rect 37461 44727 37519 44733
rect 37461 44724 37473 44727
rect 36780 44696 37473 44724
rect 36780 44684 36786 44696
rect 37461 44693 37473 44696
rect 37507 44693 37519 44727
rect 39298 44724 39304 44736
rect 39259 44696 39304 44724
rect 37461 44687 37519 44693
rect 39298 44684 39304 44696
rect 39356 44684 39362 44736
rect 41046 44684 41052 44736
rect 41104 44724 41110 44736
rect 41969 44727 42027 44733
rect 41969 44724 41981 44727
rect 41104 44696 41981 44724
rect 41104 44684 41110 44696
rect 41969 44693 41981 44696
rect 42015 44693 42027 44727
rect 43806 44724 43812 44736
rect 43767 44696 43812 44724
rect 41969 44687 42027 44693
rect 43806 44684 43812 44696
rect 43864 44684 43870 44736
rect 47118 44724 47124 44736
rect 47079 44696 47124 44724
rect 47118 44684 47124 44696
rect 47176 44684 47182 44736
rect 48958 44724 48964 44736
rect 48919 44696 48964 44724
rect 48958 44684 48964 44696
rect 49016 44684 49022 44736
rect 58526 44724 58532 44736
rect 58487 44696 58532 44724
rect 58526 44684 58532 44696
rect 58584 44684 58590 44736
rect 1104 44634 59340 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 59340 44634
rect 1104 44560 59340 44582
rect 3050 44520 3056 44532
rect 3011 44492 3056 44520
rect 3050 44480 3056 44492
rect 3108 44480 3114 44532
rect 7650 44480 7656 44532
rect 7708 44520 7714 44532
rect 7745 44523 7803 44529
rect 7745 44520 7757 44523
rect 7708 44492 7757 44520
rect 7708 44480 7714 44492
rect 7745 44489 7757 44492
rect 7791 44489 7803 44523
rect 9582 44520 9588 44532
rect 9543 44492 9588 44520
rect 7745 44483 7803 44489
rect 9582 44480 9588 44492
rect 9640 44480 9646 44532
rect 12894 44520 12900 44532
rect 12855 44492 12900 44520
rect 12894 44480 12900 44492
rect 12952 44480 12958 44532
rect 23106 44480 23112 44532
rect 23164 44520 23170 44532
rect 23201 44523 23259 44529
rect 23201 44520 23213 44523
rect 23164 44492 23213 44520
rect 23164 44480 23170 44492
rect 23201 44489 23213 44492
rect 23247 44489 23259 44523
rect 23201 44483 23259 44489
rect 31478 44480 31484 44532
rect 31536 44520 31542 44532
rect 31573 44523 31631 44529
rect 31573 44520 31585 44523
rect 31536 44492 31585 44520
rect 31536 44480 31542 44492
rect 31573 44489 31585 44492
rect 31619 44489 31631 44523
rect 31573 44483 31631 44489
rect 54018 44480 54024 44532
rect 54076 44520 54082 44532
rect 54113 44523 54171 44529
rect 54113 44520 54125 44523
rect 54076 44492 54125 44520
rect 54076 44480 54082 44492
rect 54113 44489 54125 44492
rect 54159 44489 54171 44523
rect 55950 44520 55956 44532
rect 55911 44492 55956 44520
rect 54113 44483 54171 44489
rect 55950 44480 55956 44492
rect 56008 44480 56014 44532
rect 1688 44424 5488 44452
rect 1688 44396 1716 44424
rect 1670 44384 1676 44396
rect 1583 44356 1676 44384
rect 1670 44344 1676 44356
rect 1728 44344 1734 44396
rect 1940 44387 1998 44393
rect 1940 44353 1952 44387
rect 1986 44384 1998 44387
rect 3050 44384 3056 44396
rect 1986 44356 3056 44384
rect 1986 44353 1998 44356
rect 1940 44347 1998 44353
rect 3050 44344 3056 44356
rect 3108 44344 3114 44396
rect 4356 44393 4384 44424
rect 4341 44387 4399 44393
rect 4341 44353 4353 44387
rect 4387 44353 4399 44387
rect 4341 44347 4399 44353
rect 4608 44387 4666 44393
rect 4608 44353 4620 44387
rect 4654 44384 4666 44387
rect 5350 44384 5356 44396
rect 4654 44356 5356 44384
rect 4654 44353 4666 44356
rect 4608 44347 4666 44353
rect 5350 44344 5356 44356
rect 5408 44344 5414 44396
rect 5460 44316 5488 44424
rect 7190 44412 7196 44464
rect 7248 44452 7254 44464
rect 8472 44455 8530 44461
rect 7248 44424 8248 44452
rect 7248 44412 7254 44424
rect 6632 44387 6690 44393
rect 6632 44353 6644 44387
rect 6678 44384 6690 44387
rect 7466 44384 7472 44396
rect 6678 44356 7472 44384
rect 6678 44353 6690 44356
rect 6632 44347 6690 44353
rect 7466 44344 7472 44356
rect 7524 44344 7530 44396
rect 8220 44393 8248 44424
rect 8472 44421 8484 44455
rect 8518 44452 8530 44455
rect 10410 44452 10416 44464
rect 8518 44424 10416 44452
rect 8518 44421 8530 44424
rect 8472 44415 8530 44421
rect 10410 44412 10416 44424
rect 10468 44412 10474 44464
rect 11784 44455 11842 44461
rect 11784 44421 11796 44455
rect 11830 44452 11842 44455
rect 12158 44452 12164 44464
rect 11830 44424 12164 44452
rect 11830 44421 11842 44424
rect 11784 44415 11842 44421
rect 12158 44412 12164 44424
rect 12216 44412 12222 44464
rect 13900 44455 13958 44461
rect 13900 44421 13912 44455
rect 13946 44452 13958 44455
rect 15470 44452 15476 44464
rect 13946 44424 15476 44452
rect 13946 44421 13958 44424
rect 13900 44415 13958 44421
rect 15470 44412 15476 44424
rect 15528 44412 15534 44464
rect 17212 44455 17270 44461
rect 17212 44421 17224 44455
rect 17258 44452 17270 44455
rect 18230 44452 18236 44464
rect 17258 44424 18236 44452
rect 17258 44421 17270 44424
rect 17212 44415 17270 44421
rect 18230 44412 18236 44424
rect 18288 44412 18294 44464
rect 28620 44455 28678 44461
rect 28620 44421 28632 44455
rect 28666 44452 28678 44455
rect 30282 44452 30288 44464
rect 28666 44424 30288 44452
rect 28666 44421 28678 44424
rect 28620 44415 28678 44421
rect 30282 44412 30288 44424
rect 30340 44412 30346 44464
rect 30374 44412 30380 44464
rect 30432 44412 30438 44464
rect 33778 44461 33784 44464
rect 33772 44452 33784 44461
rect 33739 44424 33784 44452
rect 33772 44415 33784 44424
rect 33778 44412 33784 44415
rect 33836 44412 33842 44464
rect 40764 44455 40822 44461
rect 40764 44421 40776 44455
rect 40810 44452 40822 44455
rect 43806 44452 43812 44464
rect 40810 44424 43812 44452
rect 40810 44421 40822 44424
rect 40764 44415 40822 44421
rect 43806 44412 43812 44424
rect 43864 44412 43870 44464
rect 45738 44412 45744 44464
rect 45796 44452 45802 44464
rect 47848 44455 47906 44461
rect 45796 44424 47624 44452
rect 45796 44412 45802 44424
rect 8205 44387 8263 44393
rect 8205 44353 8217 44387
rect 8251 44384 8263 44387
rect 10778 44384 10784 44396
rect 8251 44356 10784 44384
rect 8251 44353 8263 44356
rect 8205 44347 8263 44353
rect 10778 44344 10784 44356
rect 10836 44344 10842 44396
rect 13630 44384 13636 44396
rect 13591 44356 13636 44384
rect 13630 44344 13636 44356
rect 13688 44344 13694 44396
rect 16666 44344 16672 44396
rect 16724 44384 16730 44396
rect 16945 44387 17003 44393
rect 16945 44384 16957 44387
rect 16724 44356 16957 44384
rect 16724 44344 16730 44356
rect 16945 44353 16957 44356
rect 16991 44353 17003 44387
rect 21818 44384 21824 44396
rect 21779 44356 21824 44384
rect 16945 44347 17003 44353
rect 21818 44344 21824 44356
rect 21876 44344 21882 44396
rect 22088 44387 22146 44393
rect 22088 44353 22100 44387
rect 22134 44384 22146 44387
rect 23842 44384 23848 44396
rect 22134 44356 23848 44384
rect 22134 44353 22146 44356
rect 22088 44347 22146 44353
rect 23842 44344 23848 44356
rect 23900 44344 23906 44396
rect 25038 44384 25044 44396
rect 24999 44356 25044 44384
rect 25038 44344 25044 44356
rect 25096 44344 25102 44396
rect 25308 44387 25366 44393
rect 25308 44353 25320 44387
rect 25354 44384 25366 44387
rect 27062 44384 27068 44396
rect 25354 44356 27068 44384
rect 25354 44353 25366 44356
rect 25308 44347 25366 44353
rect 27062 44344 27068 44356
rect 27120 44344 27126 44396
rect 30193 44387 30251 44393
rect 30193 44353 30205 44387
rect 30239 44384 30251 44387
rect 30392 44384 30420 44412
rect 30239 44356 30420 44384
rect 30460 44387 30518 44393
rect 30239 44353 30251 44356
rect 30193 44347 30251 44353
rect 30460 44353 30472 44387
rect 30506 44384 30518 44387
rect 32214 44384 32220 44396
rect 30506 44356 32220 44384
rect 30506 44353 30518 44356
rect 30460 44347 30518 44353
rect 32214 44344 32220 44356
rect 32272 44344 32278 44396
rect 35345 44387 35403 44393
rect 35345 44384 35357 44387
rect 33520 44356 35357 44384
rect 6362 44316 6368 44328
rect 5460 44288 6368 44316
rect 6362 44276 6368 44288
rect 6420 44276 6426 44328
rect 9490 44276 9496 44328
rect 9548 44316 9554 44328
rect 11422 44316 11428 44328
rect 9548 44288 11428 44316
rect 9548 44276 9554 44288
rect 11422 44276 11428 44288
rect 11480 44316 11486 44328
rect 11517 44319 11575 44325
rect 11517 44316 11529 44319
rect 11480 44288 11529 44316
rect 11480 44276 11486 44288
rect 11517 44285 11529 44288
rect 11563 44285 11575 44319
rect 11517 44279 11575 44285
rect 27706 44276 27712 44328
rect 27764 44316 27770 44328
rect 28353 44319 28411 44325
rect 28353 44316 28365 44319
rect 27764 44288 28365 44316
rect 27764 44276 27770 44288
rect 28353 44285 28365 44288
rect 28399 44285 28411 44319
rect 28353 44279 28411 44285
rect 32766 44276 32772 44328
rect 32824 44316 32830 44328
rect 33520 44325 33548 44356
rect 35345 44353 35357 44356
rect 35391 44384 35403 44387
rect 35434 44384 35440 44396
rect 35391 44356 35440 44384
rect 35391 44353 35403 44356
rect 35345 44347 35403 44353
rect 35434 44344 35440 44356
rect 35492 44344 35498 44396
rect 35612 44387 35670 44393
rect 35612 44353 35624 44387
rect 35658 44384 35670 44387
rect 36630 44384 36636 44396
rect 35658 44356 36636 44384
rect 35658 44353 35670 44356
rect 35612 44347 35670 44353
rect 36630 44344 36636 44356
rect 36688 44344 36694 44396
rect 38924 44387 38982 44393
rect 38924 44353 38936 44387
rect 38970 44384 38982 44387
rect 41782 44384 41788 44396
rect 38970 44356 41788 44384
rect 38970 44353 38982 44356
rect 38924 44347 38982 44353
rect 41782 44344 41788 44356
rect 41840 44344 41846 44396
rect 42426 44344 42432 44396
rect 42484 44384 42490 44396
rect 43073 44387 43131 44393
rect 43073 44384 43085 44387
rect 42484 44356 43085 44384
rect 42484 44344 42490 44356
rect 43073 44353 43085 44356
rect 43119 44353 43131 44387
rect 43073 44347 43131 44353
rect 43340 44387 43398 44393
rect 43340 44353 43352 44387
rect 43386 44384 43398 44387
rect 44450 44384 44456 44396
rect 43386 44356 44456 44384
rect 43386 44353 43398 44356
rect 43340 44347 43398 44353
rect 44450 44344 44456 44356
rect 44508 44344 44514 44396
rect 45640 44387 45698 44393
rect 45640 44353 45652 44387
rect 45686 44384 45698 44387
rect 46658 44384 46664 44396
rect 45686 44356 46664 44384
rect 45686 44353 45698 44356
rect 45640 44347 45698 44353
rect 46658 44344 46664 44356
rect 46716 44344 46722 44396
rect 47596 44393 47624 44424
rect 47848 44421 47860 44455
rect 47894 44452 47906 44455
rect 48958 44452 48964 44464
rect 47894 44424 48964 44452
rect 47894 44421 47906 44424
rect 47848 44415 47906 44421
rect 48958 44412 48964 44424
rect 49016 44412 49022 44464
rect 53000 44455 53058 44461
rect 53000 44421 53012 44455
rect 53046 44452 53058 44455
rect 53742 44452 53748 44464
rect 53046 44424 53748 44452
rect 53046 44421 53058 44424
rect 53000 44415 53058 44421
rect 53742 44412 53748 44424
rect 53800 44412 53806 44464
rect 54840 44455 54898 44461
rect 54840 44421 54852 44455
rect 54886 44452 54898 44455
rect 55030 44452 55036 44464
rect 54886 44424 55036 44452
rect 54886 44421 54898 44424
rect 54840 44415 54898 44421
rect 55030 44412 55036 44424
rect 55088 44412 55094 44464
rect 47581 44387 47639 44393
rect 47581 44353 47593 44387
rect 47627 44384 47639 44387
rect 48314 44384 48320 44396
rect 47627 44356 48320 44384
rect 47627 44353 47639 44356
rect 47581 44347 47639 44353
rect 48314 44344 48320 44356
rect 48372 44344 48378 44396
rect 49677 44387 49735 44393
rect 49677 44384 49689 44387
rect 48976 44356 49689 44384
rect 33505 44319 33563 44325
rect 33505 44316 33517 44319
rect 32824 44288 33517 44316
rect 32824 44276 32830 44288
rect 33505 44285 33517 44288
rect 33551 44285 33563 44319
rect 33505 44279 33563 44285
rect 37918 44276 37924 44328
rect 37976 44316 37982 44328
rect 38657 44319 38715 44325
rect 38657 44316 38669 44319
rect 37976 44288 38669 44316
rect 37976 44276 37982 44288
rect 38657 44285 38669 44288
rect 38703 44285 38715 44319
rect 38657 44279 38715 44285
rect 40402 44276 40408 44328
rect 40460 44316 40466 44328
rect 40497 44319 40555 44325
rect 40497 44316 40509 44319
rect 40460 44288 40509 44316
rect 40460 44276 40466 44288
rect 40497 44285 40509 44288
rect 40543 44285 40555 44319
rect 40497 44279 40555 44285
rect 45278 44276 45284 44328
rect 45336 44316 45342 44328
rect 45373 44319 45431 44325
rect 45373 44316 45385 44319
rect 45336 44288 45385 44316
rect 45336 44276 45342 44288
rect 45373 44285 45385 44288
rect 45419 44285 45431 44319
rect 45373 44279 45431 44285
rect 48976 44257 49004 44356
rect 49677 44353 49689 44356
rect 49723 44353 49735 44387
rect 52730 44384 52736 44396
rect 52643 44356 52736 44384
rect 49677 44347 49735 44353
rect 52730 44344 52736 44356
rect 52788 44384 52794 44396
rect 53282 44384 53288 44396
rect 52788 44356 53288 44384
rect 52788 44344 52794 44356
rect 53282 44344 53288 44356
rect 53340 44384 53346 44396
rect 54570 44384 54576 44396
rect 53340 44356 54576 44384
rect 53340 44344 53346 44356
rect 54570 44344 54576 44356
rect 54628 44344 54634 44396
rect 49418 44316 49424 44328
rect 49379 44288 49424 44316
rect 49418 44276 49424 44288
rect 49476 44276 49482 44328
rect 48961 44251 49019 44257
rect 48961 44217 48973 44251
rect 49007 44217 49019 44251
rect 48961 44211 49019 44217
rect 5718 44180 5724 44192
rect 5679 44152 5724 44180
rect 5718 44140 5724 44152
rect 5776 44140 5782 44192
rect 14366 44140 14372 44192
rect 14424 44180 14430 44192
rect 15013 44183 15071 44189
rect 15013 44180 15025 44183
rect 14424 44152 15025 44180
rect 14424 44140 14430 44152
rect 15013 44149 15025 44152
rect 15059 44149 15071 44183
rect 18322 44180 18328 44192
rect 18283 44152 18328 44180
rect 15013 44143 15071 44149
rect 18322 44140 18328 44152
rect 18380 44140 18386 44192
rect 26418 44180 26424 44192
rect 26379 44152 26424 44180
rect 26418 44140 26424 44152
rect 26476 44140 26482 44192
rect 29730 44180 29736 44192
rect 29691 44152 29736 44180
rect 29730 44140 29736 44152
rect 29788 44140 29794 44192
rect 33318 44140 33324 44192
rect 33376 44180 33382 44192
rect 34885 44183 34943 44189
rect 34885 44180 34897 44183
rect 33376 44152 34897 44180
rect 33376 44140 33382 44152
rect 34885 44149 34897 44152
rect 34931 44149 34943 44183
rect 34885 44143 34943 44149
rect 36354 44140 36360 44192
rect 36412 44180 36418 44192
rect 36725 44183 36783 44189
rect 36725 44180 36737 44183
rect 36412 44152 36737 44180
rect 36412 44140 36418 44152
rect 36725 44149 36737 44152
rect 36771 44149 36783 44183
rect 40034 44180 40040 44192
rect 39995 44152 40040 44180
rect 36725 44143 36783 44149
rect 40034 44140 40040 44152
rect 40092 44140 40098 44192
rect 40770 44140 40776 44192
rect 40828 44180 40834 44192
rect 41877 44183 41935 44189
rect 41877 44180 41889 44183
rect 40828 44152 41889 44180
rect 40828 44140 40834 44152
rect 41877 44149 41889 44152
rect 41923 44149 41935 44183
rect 41877 44143 41935 44149
rect 42794 44140 42800 44192
rect 42852 44180 42858 44192
rect 44453 44183 44511 44189
rect 44453 44180 44465 44183
rect 42852 44152 44465 44180
rect 42852 44140 42858 44152
rect 44453 44149 44465 44152
rect 44499 44149 44511 44183
rect 44453 44143 44511 44149
rect 46753 44183 46811 44189
rect 46753 44149 46765 44183
rect 46799 44180 46811 44183
rect 47854 44180 47860 44192
rect 46799 44152 47860 44180
rect 46799 44149 46811 44152
rect 46753 44143 46811 44149
rect 47854 44140 47860 44152
rect 47912 44140 47918 44192
rect 49694 44140 49700 44192
rect 49752 44180 49758 44192
rect 50801 44183 50859 44189
rect 50801 44180 50813 44183
rect 49752 44152 50813 44180
rect 49752 44140 49758 44152
rect 50801 44149 50813 44152
rect 50847 44149 50859 44183
rect 50801 44143 50859 44149
rect 1104 44090 59340 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 59340 44090
rect 1104 44016 59340 44038
rect 6362 43936 6368 43988
rect 6420 43976 6426 43988
rect 6822 43976 6828 43988
rect 6420 43948 6828 43976
rect 6420 43936 6426 43948
rect 6822 43936 6828 43948
rect 6880 43976 6886 43988
rect 6917 43979 6975 43985
rect 6917 43976 6929 43979
rect 6880 43948 6929 43976
rect 6880 43936 6886 43948
rect 6917 43945 6929 43948
rect 6963 43945 6975 43979
rect 23842 43976 23848 43988
rect 23803 43948 23848 43976
rect 6917 43939 6975 43945
rect 23842 43936 23848 43948
rect 23900 43936 23906 43988
rect 27062 43976 27068 43988
rect 27023 43948 27068 43976
rect 27062 43936 27068 43948
rect 27120 43936 27126 43988
rect 27522 43936 27528 43988
rect 27580 43976 27586 43988
rect 28905 43979 28963 43985
rect 28905 43976 28917 43979
rect 27580 43948 28917 43976
rect 27580 43936 27586 43948
rect 28905 43945 28917 43948
rect 28951 43945 28963 43979
rect 32214 43976 32220 43988
rect 32175 43948 32220 43976
rect 28905 43939 28963 43945
rect 32214 43936 32220 43948
rect 32272 43936 32278 43988
rect 35434 43936 35440 43988
rect 35492 43976 35498 43988
rect 36357 43979 36415 43985
rect 36357 43976 36369 43979
rect 35492 43948 36369 43976
rect 35492 43936 35498 43948
rect 36357 43945 36369 43948
rect 36403 43945 36415 43979
rect 36357 43939 36415 43945
rect 39206 43936 39212 43988
rect 39264 43976 39270 43988
rect 39301 43979 39359 43985
rect 39301 43976 39313 43979
rect 39264 43948 39313 43976
rect 39264 43936 39270 43948
rect 39301 43945 39313 43948
rect 39347 43945 39359 43979
rect 39301 43939 39359 43945
rect 42613 43979 42671 43985
rect 42613 43945 42625 43979
rect 42659 43976 42671 43979
rect 42702 43976 42708 43988
rect 42659 43948 42708 43976
rect 42659 43945 42671 43948
rect 42613 43939 42671 43945
rect 42702 43936 42708 43948
rect 42760 43936 42766 43988
rect 45646 43976 45652 43988
rect 43088 43948 45652 43976
rect 1670 43800 1676 43852
rect 1728 43840 1734 43852
rect 1857 43843 1915 43849
rect 1857 43840 1869 43843
rect 1728 43812 1869 43840
rect 1728 43800 1734 43812
rect 1857 43809 1869 43812
rect 1903 43809 1915 43843
rect 14090 43840 14096 43852
rect 14051 43812 14096 43840
rect 1857 43803 1915 43809
rect 14090 43800 14096 43812
rect 14148 43800 14154 43852
rect 16666 43800 16672 43852
rect 16724 43840 16730 43852
rect 17126 43840 17132 43852
rect 16724 43812 17132 43840
rect 16724 43800 16730 43812
rect 17126 43800 17132 43812
rect 17184 43800 17190 43852
rect 25038 43800 25044 43852
rect 25096 43840 25102 43852
rect 25590 43840 25596 43852
rect 25096 43812 25596 43840
rect 25096 43800 25102 43812
rect 25590 43800 25596 43812
rect 25648 43840 25654 43852
rect 25685 43843 25743 43849
rect 25685 43840 25697 43843
rect 25648 43812 25697 43840
rect 25648 43800 25654 43812
rect 25685 43809 25697 43812
rect 25731 43809 25743 43843
rect 25685 43803 25743 43809
rect 30374 43800 30380 43852
rect 30432 43840 30438 43852
rect 43088 43849 43116 43948
rect 45646 43936 45652 43948
rect 45704 43936 45710 43988
rect 46658 43976 46664 43988
rect 46619 43948 46664 43976
rect 46658 43936 46664 43948
rect 46716 43936 46722 43988
rect 53374 43976 53380 43988
rect 53335 43948 53380 43976
rect 53374 43936 53380 43948
rect 53432 43936 53438 43988
rect 44450 43908 44456 43920
rect 44411 43880 44456 43908
rect 44450 43868 44456 43880
rect 44508 43868 44514 43920
rect 30837 43843 30895 43849
rect 30837 43840 30849 43843
rect 30432 43812 30849 43840
rect 30432 43800 30438 43812
rect 30837 43809 30849 43812
rect 30883 43809 30895 43843
rect 30837 43803 30895 43809
rect 43073 43843 43131 43849
rect 43073 43809 43085 43843
rect 43119 43809 43131 43843
rect 56502 43840 56508 43852
rect 56463 43812 56508 43840
rect 43073 43803 43131 43809
rect 2124 43775 2182 43781
rect 2124 43741 2136 43775
rect 2170 43772 2182 43775
rect 7742 43772 7748 43784
rect 2170 43744 7748 43772
rect 2170 43741 2182 43744
rect 2124 43735 2182 43741
rect 7742 43732 7748 43744
rect 7800 43732 7806 43784
rect 9582 43772 9588 43784
rect 9543 43744 9588 43772
rect 9582 43732 9588 43744
rect 9640 43732 9646 43784
rect 11422 43732 11428 43784
rect 11480 43772 11486 43784
rect 14366 43781 14372 43784
rect 12161 43775 12219 43781
rect 12161 43772 12173 43775
rect 11480 43744 12173 43772
rect 11480 43732 11486 43744
rect 12161 43741 12173 43744
rect 12207 43741 12219 43775
rect 14360 43772 14372 43781
rect 14327 43744 14372 43772
rect 12161 43735 12219 43741
rect 14360 43735 14372 43744
rect 14366 43732 14372 43735
rect 14424 43732 14430 43784
rect 17396 43775 17454 43781
rect 17396 43741 17408 43775
rect 17442 43772 17454 43775
rect 18322 43772 18328 43784
rect 17442 43744 18328 43772
rect 17442 43741 17454 43744
rect 17396 43735 17454 43741
rect 18322 43732 18328 43744
rect 18380 43732 18386 43784
rect 21542 43732 21548 43784
rect 21600 43772 21606 43784
rect 22465 43775 22523 43781
rect 22465 43772 22477 43775
rect 21600 43744 22477 43772
rect 21600 43732 21606 43744
rect 22465 43741 22477 43744
rect 22511 43741 22523 43775
rect 22465 43735 22523 43741
rect 25952 43775 26010 43781
rect 25952 43741 25964 43775
rect 25998 43772 26010 43775
rect 27154 43772 27160 43784
rect 25998 43744 27160 43772
rect 25998 43741 26010 43744
rect 25952 43735 26010 43741
rect 27154 43732 27160 43744
rect 27212 43732 27218 43784
rect 27525 43775 27583 43781
rect 27525 43741 27537 43775
rect 27571 43772 27583 43775
rect 27792 43775 27850 43781
rect 27571 43744 27752 43772
rect 27571 43741 27583 43744
rect 27525 43735 27583 43741
rect 27724 43716 27752 43744
rect 27792 43741 27804 43775
rect 27838 43772 27850 43775
rect 29178 43772 29184 43784
rect 27838 43744 29184 43772
rect 27838 43741 27850 43744
rect 27792 43735 27850 43741
rect 29178 43732 29184 43744
rect 29236 43732 29242 43784
rect 5626 43704 5632 43716
rect 5587 43676 5632 43704
rect 5626 43664 5632 43676
rect 5684 43704 5690 43716
rect 9674 43704 9680 43716
rect 5684 43676 9680 43704
rect 5684 43664 5690 43676
rect 9674 43664 9680 43676
rect 9732 43664 9738 43716
rect 9852 43707 9910 43713
rect 9852 43673 9864 43707
rect 9898 43704 9910 43707
rect 10870 43704 10876 43716
rect 9898 43676 10876 43704
rect 9898 43673 9910 43676
rect 9852 43667 9910 43673
rect 10870 43664 10876 43676
rect 10928 43664 10934 43716
rect 12428 43707 12486 43713
rect 12428 43673 12440 43707
rect 12474 43704 12486 43707
rect 14826 43704 14832 43716
rect 12474 43676 14832 43704
rect 12474 43673 12486 43676
rect 12428 43667 12486 43673
rect 14826 43664 14832 43676
rect 14884 43664 14890 43716
rect 20257 43707 20315 43713
rect 20257 43673 20269 43707
rect 20303 43704 20315 43707
rect 20530 43704 20536 43716
rect 20303 43676 20536 43704
rect 20303 43673 20315 43676
rect 20257 43667 20315 43673
rect 20530 43664 20536 43676
rect 20588 43664 20594 43716
rect 22732 43707 22790 43713
rect 22732 43673 22744 43707
rect 22778 43704 22790 43707
rect 23198 43704 23204 43716
rect 22778 43676 23204 43704
rect 22778 43673 22790 43676
rect 22732 43667 22790 43673
rect 23198 43664 23204 43676
rect 23256 43664 23262 43716
rect 27706 43664 27712 43716
rect 27764 43664 27770 43716
rect 30852 43704 30880 43803
rect 56502 43800 56508 43812
rect 56560 43800 56566 43852
rect 31104 43775 31162 43781
rect 31104 43741 31116 43775
rect 31150 43772 31162 43775
rect 31938 43772 31944 43784
rect 31150 43744 31944 43772
rect 31150 43741 31162 43744
rect 31104 43735 31162 43741
rect 31938 43732 31944 43744
rect 31996 43732 32002 43784
rect 32766 43772 32772 43784
rect 32679 43744 32772 43772
rect 32766 43732 32772 43744
rect 32824 43732 32830 43784
rect 33036 43775 33094 43781
rect 33036 43741 33048 43775
rect 33082 43772 33094 43775
rect 33318 43772 33324 43784
rect 33082 43744 33324 43772
rect 33082 43741 33094 43744
rect 33036 43735 33094 43741
rect 33318 43732 33324 43744
rect 33376 43732 33382 43784
rect 37366 43732 37372 43784
rect 37424 43772 37430 43784
rect 37918 43772 37924 43784
rect 37424 43744 37924 43772
rect 37424 43732 37430 43744
rect 37918 43732 37924 43744
rect 37976 43732 37982 43784
rect 38188 43775 38246 43781
rect 38188 43741 38200 43775
rect 38234 43772 38246 43775
rect 39298 43772 39304 43784
rect 38234 43744 39304 43772
rect 38234 43741 38246 43744
rect 38188 43735 38246 43741
rect 39298 43732 39304 43744
rect 39356 43732 39362 43784
rect 40494 43732 40500 43784
rect 40552 43772 40558 43784
rect 41233 43775 41291 43781
rect 41233 43772 41245 43775
rect 40552 43744 41245 43772
rect 40552 43732 40558 43744
rect 41233 43741 41245 43744
rect 41279 43741 41291 43775
rect 41233 43735 41291 43741
rect 41500 43775 41558 43781
rect 41500 43741 41512 43775
rect 41546 43772 41558 43775
rect 42794 43772 42800 43784
rect 41546 43744 42800 43772
rect 41546 43741 41558 43744
rect 41500 43735 41558 43741
rect 42794 43732 42800 43744
rect 42852 43732 42858 43784
rect 44450 43732 44456 43784
rect 44508 43772 44514 43784
rect 45278 43772 45284 43784
rect 44508 43744 45284 43772
rect 44508 43732 44514 43744
rect 45278 43732 45284 43744
rect 45336 43732 45342 43784
rect 47118 43772 47124 43784
rect 45388 43744 47124 43772
rect 32784 43704 32812 43732
rect 30852 43676 32812 43704
rect 32950 43664 32956 43716
rect 33008 43704 33014 43716
rect 35069 43707 35127 43713
rect 35069 43704 35081 43707
rect 33008 43676 35081 43704
rect 33008 43664 33014 43676
rect 35069 43673 35081 43676
rect 35115 43704 35127 43707
rect 39206 43704 39212 43716
rect 35115 43676 39212 43704
rect 35115 43673 35127 43676
rect 35069 43667 35127 43673
rect 39206 43664 39212 43676
rect 39264 43664 39270 43716
rect 43340 43707 43398 43713
rect 43340 43673 43352 43707
rect 43386 43704 43398 43707
rect 45388 43704 45416 43744
rect 47118 43732 47124 43744
rect 47176 43732 47182 43784
rect 50157 43775 50215 43781
rect 50157 43741 50169 43775
rect 50203 43772 50215 43775
rect 51997 43775 52055 43781
rect 50203 43744 51672 43772
rect 50203 43741 50215 43744
rect 50157 43735 50215 43741
rect 51644 43716 51672 43744
rect 51997 43741 52009 43775
rect 52043 43741 52055 43775
rect 51997 43735 52055 43741
rect 43386 43676 45416 43704
rect 45548 43707 45606 43713
rect 43386 43673 43398 43676
rect 43340 43667 43398 43673
rect 45548 43673 45560 43707
rect 45594 43704 45606 43707
rect 46474 43704 46480 43716
rect 45594 43676 46480 43704
rect 45594 43673 45606 43676
rect 45548 43667 45606 43673
rect 46474 43664 46480 43676
rect 46532 43664 46538 43716
rect 47857 43707 47915 43713
rect 47857 43673 47869 43707
rect 47903 43704 47915 43707
rect 47946 43704 47952 43716
rect 47903 43676 47952 43704
rect 47903 43673 47915 43676
rect 47857 43667 47915 43673
rect 47946 43664 47952 43676
rect 48004 43664 48010 43716
rect 49602 43664 49608 43716
rect 49660 43704 49666 43716
rect 50402 43707 50460 43713
rect 50402 43704 50414 43707
rect 49660 43676 50414 43704
rect 49660 43664 49666 43676
rect 50402 43673 50414 43676
rect 50448 43673 50460 43707
rect 50402 43667 50460 43673
rect 51626 43664 51632 43716
rect 51684 43704 51690 43716
rect 52012 43704 52040 43735
rect 52086 43732 52092 43784
rect 52144 43772 52150 43784
rect 52253 43775 52311 43781
rect 52253 43772 52265 43775
rect 52144 43744 52265 43772
rect 52144 43732 52150 43744
rect 52253 43741 52265 43744
rect 52299 43741 52311 43775
rect 52253 43735 52311 43741
rect 56772 43775 56830 43781
rect 56772 43741 56784 43775
rect 56818 43772 56830 43775
rect 58526 43772 58532 43784
rect 56818 43744 58532 43772
rect 56818 43741 56830 43744
rect 56772 43735 56830 43741
rect 58526 43732 58532 43744
rect 58584 43732 58590 43784
rect 53282 43704 53288 43716
rect 51684 43676 53288 43704
rect 51684 43664 51690 43676
rect 53282 43664 53288 43676
rect 53340 43664 53346 43716
rect 3234 43636 3240 43648
rect 3195 43608 3240 43636
rect 3234 43596 3240 43608
rect 3292 43596 3298 43648
rect 10965 43639 11023 43645
rect 10965 43605 10977 43639
rect 11011 43636 11023 43639
rect 11514 43636 11520 43648
rect 11011 43608 11520 43636
rect 11011 43605 11023 43608
rect 10965 43599 11023 43605
rect 11514 43596 11520 43608
rect 11572 43596 11578 43648
rect 13538 43636 13544 43648
rect 13499 43608 13544 43636
rect 13538 43596 13544 43608
rect 13596 43596 13602 43648
rect 15470 43636 15476 43648
rect 15431 43608 15476 43636
rect 15470 43596 15476 43608
rect 15528 43596 15534 43648
rect 18506 43636 18512 43648
rect 18467 43608 18512 43636
rect 18506 43596 18512 43608
rect 18564 43596 18570 43648
rect 21542 43636 21548 43648
rect 21503 43608 21548 43636
rect 21542 43596 21548 43608
rect 21600 43596 21606 43648
rect 34146 43636 34152 43648
rect 34107 43608 34152 43636
rect 34146 43596 34152 43608
rect 34204 43596 34210 43648
rect 48314 43596 48320 43648
rect 48372 43636 48378 43648
rect 49145 43639 49203 43645
rect 49145 43636 49157 43639
rect 48372 43608 49157 43636
rect 48372 43596 48378 43608
rect 49145 43605 49157 43608
rect 49191 43636 49203 43639
rect 49418 43636 49424 43648
rect 49191 43608 49424 43636
rect 49191 43605 49203 43608
rect 49145 43599 49203 43605
rect 49418 43596 49424 43608
rect 49476 43596 49482 43648
rect 51534 43636 51540 43648
rect 51495 43608 51540 43636
rect 51534 43596 51540 43608
rect 51592 43596 51598 43648
rect 57882 43636 57888 43648
rect 57843 43608 57888 43636
rect 57882 43596 57888 43608
rect 57940 43596 57946 43648
rect 1104 43546 59340 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 59340 43546
rect 1104 43472 59340 43494
rect 3050 43432 3056 43444
rect 3011 43404 3056 43432
rect 3050 43392 3056 43404
rect 3108 43392 3114 43444
rect 5350 43432 5356 43444
rect 5311 43404 5356 43432
rect 5350 43392 5356 43404
rect 5408 43392 5414 43444
rect 7466 43392 7472 43444
rect 7524 43432 7530 43444
rect 7745 43435 7803 43441
rect 7745 43432 7757 43435
rect 7524 43404 7757 43432
rect 7524 43392 7530 43404
rect 7745 43401 7757 43404
rect 7791 43401 7803 43435
rect 14826 43432 14832 43444
rect 14787 43404 14832 43432
rect 7745 43395 7803 43401
rect 14826 43392 14832 43404
rect 14884 43392 14890 43444
rect 20530 43392 20536 43444
rect 20588 43432 20594 43444
rect 23198 43432 23204 43444
rect 20588 43404 22775 43432
rect 23159 43404 23204 43432
rect 20588 43392 20594 43404
rect 1940 43367 1998 43373
rect 1940 43333 1952 43367
rect 1986 43364 1998 43367
rect 3234 43364 3240 43376
rect 1986 43336 3240 43364
rect 1986 43333 1998 43336
rect 1940 43327 1998 43333
rect 3234 43324 3240 43336
rect 3292 43324 3298 43376
rect 5718 43324 5724 43376
rect 5776 43364 5782 43376
rect 6610 43367 6668 43373
rect 6610 43364 6622 43367
rect 5776 43336 6622 43364
rect 5776 43324 5782 43336
rect 6610 43333 6622 43336
rect 6656 43333 6668 43367
rect 6610 43327 6668 43333
rect 6822 43324 6828 43376
rect 6880 43324 6886 43376
rect 13716 43367 13774 43373
rect 13716 43333 13728 43367
rect 13762 43364 13774 43367
rect 15470 43364 15476 43376
rect 13762 43336 15476 43364
rect 13762 43333 13774 43336
rect 13716 43327 13774 43333
rect 15470 43324 15476 43336
rect 15528 43324 15534 43376
rect 17488 43367 17546 43373
rect 17488 43333 17500 43367
rect 17534 43364 17546 43367
rect 18506 43364 18512 43376
rect 17534 43336 18512 43364
rect 17534 43333 17546 43336
rect 17488 43327 17546 43333
rect 18506 43324 18512 43336
rect 18564 43324 18570 43376
rect 22646 43364 22652 43376
rect 21836 43336 22652 43364
rect 1670 43296 1676 43308
rect 1631 43268 1676 43296
rect 1670 43256 1676 43268
rect 1728 43256 1734 43308
rect 4240 43299 4298 43305
rect 4240 43265 4252 43299
rect 4286 43296 4298 43299
rect 5166 43296 5172 43308
rect 4286 43268 5172 43296
rect 4286 43265 4298 43268
rect 4240 43259 4298 43265
rect 5166 43256 5172 43268
rect 5224 43256 5230 43308
rect 6365 43299 6423 43305
rect 6365 43265 6377 43299
rect 6411 43296 6423 43299
rect 6840 43296 6868 43324
rect 21836 43308 21864 43336
rect 22646 43324 22652 43336
rect 22704 43324 22710 43376
rect 22747 43364 22775 43404
rect 23198 43392 23204 43404
rect 23256 43392 23262 43444
rect 25590 43392 25596 43444
rect 25648 43432 25654 43444
rect 25777 43435 25835 43441
rect 25777 43432 25789 43435
rect 25648 43404 25789 43432
rect 25648 43392 25654 43404
rect 25777 43401 25789 43404
rect 25823 43401 25835 43435
rect 25777 43395 25835 43401
rect 30098 43392 30104 43444
rect 30156 43432 30162 43444
rect 30469 43435 30527 43441
rect 30469 43432 30481 43435
rect 30156 43404 30481 43432
rect 30156 43392 30162 43404
rect 30469 43401 30481 43404
rect 30515 43401 30527 43435
rect 30469 43395 30527 43401
rect 34790 43392 34796 43444
rect 34848 43432 34854 43444
rect 34885 43435 34943 43441
rect 34885 43432 34897 43435
rect 34848 43404 34897 43432
rect 34848 43392 34854 43404
rect 34885 43401 34897 43404
rect 34931 43401 34943 43435
rect 34885 43395 34943 43401
rect 35342 43392 35348 43444
rect 35400 43392 35406 43444
rect 38010 43392 38016 43444
rect 38068 43432 38074 43444
rect 38749 43435 38807 43441
rect 38749 43432 38761 43435
rect 38068 43404 38761 43432
rect 38068 43392 38074 43404
rect 38749 43401 38761 43404
rect 38795 43401 38807 43435
rect 46474 43432 46480 43444
rect 46435 43404 46480 43432
rect 38749 43395 38807 43401
rect 46474 43392 46480 43404
rect 46532 43392 46538 43444
rect 49602 43432 49608 43444
rect 49563 43404 49608 43432
rect 49602 43392 49608 43404
rect 49660 43392 49666 43444
rect 54570 43432 54576 43444
rect 54531 43404 54576 43432
rect 54570 43392 54576 43404
rect 54628 43392 54634 43444
rect 24489 43367 24547 43373
rect 24489 43364 24501 43367
rect 22747 43336 24501 43364
rect 24489 43333 24501 43336
rect 24535 43364 24547 43367
rect 27338 43364 27344 43376
rect 24535 43336 27344 43364
rect 24535 43333 24547 43336
rect 24489 43327 24547 43333
rect 27338 43324 27344 43336
rect 27396 43324 27402 43376
rect 27706 43364 27712 43376
rect 27448 43336 27712 43364
rect 6411 43268 6868 43296
rect 9852 43299 9910 43305
rect 6411 43265 6423 43268
rect 6365 43259 6423 43265
rect 9852 43265 9864 43299
rect 9898 43296 9910 43299
rect 10962 43296 10968 43308
rect 9898 43268 10968 43296
rect 9898 43265 9910 43268
rect 9852 43259 9910 43265
rect 10962 43256 10968 43268
rect 11020 43256 11026 43308
rect 11876 43299 11934 43305
rect 11876 43265 11888 43299
rect 11922 43296 11934 43299
rect 13354 43296 13360 43308
rect 11922 43268 13360 43296
rect 11922 43265 11934 43268
rect 11876 43259 11934 43265
rect 13354 43256 13360 43268
rect 13412 43256 13418 43308
rect 13449 43299 13507 43305
rect 13449 43265 13461 43299
rect 13495 43296 13507 43299
rect 14090 43296 14096 43308
rect 13495 43268 14096 43296
rect 13495 43265 13507 43268
rect 13449 43259 13507 43265
rect 14090 43256 14096 43268
rect 14148 43256 14154 43308
rect 17126 43256 17132 43308
rect 17184 43296 17190 43308
rect 17221 43299 17279 43305
rect 17221 43296 17233 43299
rect 17184 43268 17233 43296
rect 17184 43256 17190 43268
rect 17221 43265 17233 43268
rect 17267 43296 17279 43299
rect 19242 43296 19248 43308
rect 17267 43268 19248 43296
rect 17267 43265 17279 43268
rect 17221 43259 17279 43265
rect 19242 43256 19248 43268
rect 19300 43256 19306 43308
rect 19334 43256 19340 43308
rect 19392 43296 19398 43308
rect 19501 43299 19559 43305
rect 19501 43296 19513 43299
rect 19392 43268 19513 43296
rect 19392 43256 19398 43268
rect 19501 43265 19513 43268
rect 19547 43265 19559 43299
rect 21818 43296 21824 43308
rect 21779 43268 21824 43296
rect 19501 43259 19559 43265
rect 21818 43256 21824 43268
rect 21876 43256 21882 43308
rect 22088 43299 22146 43305
rect 22088 43265 22100 43299
rect 22134 43296 22146 43299
rect 23658 43296 23664 43308
rect 22134 43268 23664 43296
rect 22134 43265 22146 43268
rect 22088 43259 22146 43265
rect 23658 43256 23664 43268
rect 23716 43256 23722 43308
rect 27249 43299 27307 43305
rect 27249 43265 27261 43299
rect 27295 43296 27307 43299
rect 27448 43296 27476 43336
rect 27706 43324 27712 43336
rect 27764 43364 27770 43376
rect 29356 43367 29414 43373
rect 27764 43336 29132 43364
rect 27764 43324 27770 43336
rect 27295 43268 27476 43296
rect 27516 43299 27574 43305
rect 27295 43265 27307 43268
rect 27249 43259 27307 43265
rect 27516 43265 27528 43299
rect 27562 43296 27574 43299
rect 28902 43296 28908 43308
rect 27562 43268 28908 43296
rect 27562 43265 27574 43268
rect 27516 43259 27574 43265
rect 28902 43256 28908 43268
rect 28960 43256 28966 43308
rect 29104 43305 29132 43336
rect 29356 43333 29368 43367
rect 29402 43364 29414 43367
rect 29730 43364 29736 43376
rect 29402 43336 29736 43364
rect 29402 43333 29414 43336
rect 29356 43327 29414 43333
rect 29730 43324 29736 43336
rect 29788 43324 29794 43376
rect 33772 43367 33830 43373
rect 33772 43333 33784 43367
rect 33818 43364 33830 43367
rect 35360 43364 35388 43392
rect 33818 43336 35388 43364
rect 35612 43367 35670 43373
rect 33818 43333 33830 43336
rect 33772 43327 33830 43333
rect 35612 43333 35624 43367
rect 35658 43364 35670 43367
rect 36722 43364 36728 43376
rect 35658 43336 36728 43364
rect 35658 43333 35670 43336
rect 35612 43327 35670 43333
rect 36722 43324 36728 43336
rect 36780 43324 36786 43376
rect 37636 43367 37694 43373
rect 37636 43333 37648 43367
rect 37682 43364 37694 43367
rect 39390 43364 39396 43376
rect 37682 43336 39396 43364
rect 37682 43333 37694 43336
rect 37636 43327 37694 43333
rect 39390 43324 39396 43336
rect 39448 43324 39454 43376
rect 42696 43367 42754 43373
rect 42696 43333 42708 43367
rect 42742 43364 42754 43367
rect 46198 43364 46204 43376
rect 42742 43336 46204 43364
rect 42742 43333 42754 43336
rect 42696 43327 42754 43333
rect 46198 43324 46204 43336
rect 46256 43324 46262 43376
rect 48492 43367 48550 43373
rect 48492 43333 48504 43367
rect 48538 43364 48550 43367
rect 49694 43364 49700 43376
rect 48538 43336 49700 43364
rect 48538 43333 48550 43336
rect 48492 43327 48550 43333
rect 49694 43324 49700 43336
rect 49752 43324 49758 43376
rect 50332 43367 50390 43373
rect 50332 43333 50344 43367
rect 50378 43364 50390 43367
rect 51534 43364 51540 43376
rect 50378 43336 51540 43364
rect 50378 43333 50390 43336
rect 50332 43327 50390 43333
rect 51534 43324 51540 43336
rect 51592 43324 51598 43376
rect 56502 43364 56508 43376
rect 55968 43336 56508 43364
rect 29089 43299 29147 43305
rect 29089 43265 29101 43299
rect 29135 43265 29147 43299
rect 29089 43259 29147 43265
rect 32766 43256 32772 43308
rect 32824 43296 32830 43308
rect 33505 43299 33563 43305
rect 33505 43296 33517 43299
rect 32824 43268 33517 43296
rect 32824 43256 32830 43268
rect 33505 43265 33517 43268
rect 33551 43265 33563 43299
rect 33505 43259 33563 43265
rect 35345 43299 35403 43305
rect 35345 43265 35357 43299
rect 35391 43296 35403 43299
rect 39206 43296 39212 43308
rect 35391 43268 37412 43296
rect 39167 43268 39212 43296
rect 35391 43265 35403 43268
rect 35345 43259 35403 43265
rect 37384 43240 37412 43268
rect 39206 43256 39212 43268
rect 39264 43296 39270 43308
rect 40310 43296 40316 43308
rect 39264 43268 40316 43296
rect 39264 43256 39270 43268
rect 40310 43256 40316 43268
rect 40368 43256 40374 43308
rect 45097 43299 45155 43305
rect 45097 43265 45109 43299
rect 45143 43296 45155 43299
rect 45186 43296 45192 43308
rect 45143 43268 45192 43296
rect 45143 43265 45155 43268
rect 45097 43259 45155 43265
rect 45186 43256 45192 43268
rect 45244 43256 45250 43308
rect 45364 43299 45422 43305
rect 45364 43265 45376 43299
rect 45410 43296 45422 43299
rect 46382 43296 46388 43308
rect 45410 43268 46388 43296
rect 45410 43265 45422 43268
rect 45364 43259 45422 43265
rect 46382 43256 46388 43268
rect 46440 43256 46446 43308
rect 48225 43299 48283 43305
rect 48225 43265 48237 43299
rect 48271 43296 48283 43299
rect 48314 43296 48320 43308
rect 48271 43268 48320 43296
rect 48271 43265 48283 43268
rect 48225 43259 48283 43265
rect 48314 43256 48320 43268
rect 48372 43256 48378 43308
rect 49418 43256 49424 43308
rect 49476 43296 49482 43308
rect 50065 43299 50123 43305
rect 50065 43296 50077 43299
rect 49476 43268 50077 43296
rect 49476 43256 49482 43268
rect 50065 43265 50077 43268
rect 50111 43265 50123 43299
rect 53098 43296 53104 43308
rect 53059 43268 53104 43296
rect 50065 43259 50123 43265
rect 53098 43256 53104 43268
rect 53156 43296 53162 43308
rect 55582 43296 55588 43308
rect 53156 43268 55588 43296
rect 53156 43256 53162 43268
rect 55582 43256 55588 43268
rect 55640 43256 55646 43308
rect 55968 43305 55996 43336
rect 56502 43324 56508 43336
rect 56560 43324 56566 43376
rect 55953 43299 56011 43305
rect 55953 43265 55965 43299
rect 55999 43265 56011 43299
rect 55953 43259 56011 43265
rect 56220 43299 56278 43305
rect 56220 43265 56232 43299
rect 56266 43296 56278 43299
rect 58158 43296 58164 43308
rect 56266 43268 58164 43296
rect 56266 43265 56278 43268
rect 56220 43259 56278 43265
rect 58158 43256 58164 43268
rect 58216 43256 58222 43308
rect 3786 43188 3792 43240
rect 3844 43228 3850 43240
rect 3973 43231 4031 43237
rect 3973 43228 3985 43231
rect 3844 43200 3985 43228
rect 3844 43188 3850 43200
rect 3973 43197 3985 43200
rect 4019 43197 4031 43231
rect 9582 43228 9588 43240
rect 9543 43200 9588 43228
rect 3973 43191 4031 43197
rect 9582 43188 9588 43200
rect 9640 43188 9646 43240
rect 11422 43188 11428 43240
rect 11480 43228 11486 43240
rect 11609 43231 11667 43237
rect 11609 43228 11621 43231
rect 11480 43200 11621 43228
rect 11480 43188 11486 43200
rect 11609 43197 11621 43200
rect 11655 43197 11667 43231
rect 37366 43228 37372 43240
rect 37327 43200 37372 43228
rect 11609 43191 11667 43197
rect 37366 43188 37372 43200
rect 37424 43188 37430 43240
rect 42426 43228 42432 43240
rect 42387 43200 42432 43228
rect 42426 43188 42432 43200
rect 42484 43188 42490 43240
rect 36630 43120 36636 43172
rect 36688 43160 36694 43172
rect 36725 43163 36783 43169
rect 36725 43160 36737 43163
rect 36688 43132 36737 43160
rect 36688 43120 36694 43132
rect 36725 43129 36737 43132
rect 36771 43129 36783 43163
rect 36725 43123 36783 43129
rect 9490 43052 9496 43104
rect 9548 43092 9554 43104
rect 10965 43095 11023 43101
rect 10965 43092 10977 43095
rect 9548 43064 10977 43092
rect 9548 43052 9554 43064
rect 10965 43061 10977 43064
rect 11011 43061 11023 43095
rect 10965 43055 11023 43061
rect 12618 43052 12624 43104
rect 12676 43092 12682 43104
rect 12989 43095 13047 43101
rect 12989 43092 13001 43095
rect 12676 43064 13001 43092
rect 12676 43052 12682 43064
rect 12989 43061 13001 43064
rect 13035 43061 13047 43095
rect 18598 43092 18604 43104
rect 18559 43064 18604 43092
rect 12989 43055 13047 43061
rect 18598 43052 18604 43064
rect 18656 43052 18662 43104
rect 18782 43052 18788 43104
rect 18840 43092 18846 43104
rect 20625 43095 20683 43101
rect 20625 43092 20637 43095
rect 18840 43064 20637 43092
rect 18840 43052 18846 43064
rect 20625 43061 20637 43064
rect 20671 43061 20683 43095
rect 20625 43055 20683 43061
rect 27430 43052 27436 43104
rect 27488 43092 27494 43104
rect 28629 43095 28687 43101
rect 28629 43092 28641 43095
rect 27488 43064 28641 43092
rect 27488 43052 27494 43064
rect 28629 43061 28641 43064
rect 28675 43061 28687 43095
rect 40494 43092 40500 43104
rect 40455 43064 40500 43092
rect 28629 43055 28687 43061
rect 40494 43052 40500 43064
rect 40552 43052 40558 43104
rect 43070 43052 43076 43104
rect 43128 43092 43134 43104
rect 43809 43095 43867 43101
rect 43809 43092 43821 43095
rect 43128 43064 43821 43092
rect 43128 43052 43134 43064
rect 43809 43061 43821 43064
rect 43855 43061 43867 43095
rect 51442 43092 51448 43104
rect 51403 43064 51448 43092
rect 43809 43055 43867 43061
rect 51442 43052 51448 43064
rect 51500 43052 51506 43104
rect 57330 43092 57336 43104
rect 57291 43064 57336 43092
rect 57330 43052 57336 43064
rect 57388 43052 57394 43104
rect 1104 43002 59340 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 59340 43002
rect 1104 42928 59340 42950
rect 5166 42888 5172 42900
rect 5127 42860 5172 42888
rect 5166 42848 5172 42860
rect 5224 42848 5230 42900
rect 11422 42848 11428 42900
rect 11480 42888 11486 42900
rect 11517 42891 11575 42897
rect 11517 42888 11529 42891
rect 11480 42860 11529 42888
rect 11480 42848 11486 42860
rect 11517 42857 11529 42860
rect 11563 42857 11575 42891
rect 23658 42888 23664 42900
rect 23619 42860 23664 42888
rect 11517 42851 11575 42857
rect 23658 42848 23664 42860
rect 23716 42848 23722 42900
rect 42518 42848 42524 42900
rect 42576 42888 42582 42900
rect 44450 42888 44456 42900
rect 42576 42860 44456 42888
rect 42576 42848 42582 42860
rect 44450 42848 44456 42860
rect 44508 42848 44514 42900
rect 46382 42888 46388 42900
rect 46343 42860 46388 42888
rect 46382 42848 46388 42860
rect 46440 42848 46446 42900
rect 48314 42888 48320 42900
rect 47596 42860 48320 42888
rect 19242 42780 19248 42832
rect 19300 42820 19306 42832
rect 19300 42792 19380 42820
rect 19300 42780 19306 42792
rect 6822 42712 6828 42764
rect 6880 42752 6886 42764
rect 7009 42755 7067 42761
rect 7009 42752 7021 42755
rect 6880 42724 7021 42752
rect 6880 42712 6886 42724
rect 7009 42721 7021 42724
rect 7055 42721 7067 42755
rect 7009 42715 7067 42721
rect 17126 42712 17132 42764
rect 17184 42752 17190 42764
rect 17313 42755 17371 42761
rect 17313 42752 17325 42755
rect 17184 42724 17325 42752
rect 17184 42712 17190 42724
rect 17313 42721 17325 42724
rect 17359 42721 17371 42755
rect 19352 42752 19380 42792
rect 19978 42752 19984 42764
rect 19352 42724 19984 42752
rect 17313 42715 17371 42721
rect 19978 42712 19984 42724
rect 20036 42752 20042 42764
rect 47596 42761 47624 42860
rect 48314 42848 48320 42860
rect 48372 42848 48378 42900
rect 58158 42888 58164 42900
rect 58119 42860 58164 42888
rect 58158 42848 58164 42860
rect 58216 42848 58222 42900
rect 20441 42755 20499 42761
rect 20441 42752 20453 42755
rect 20036 42724 20453 42752
rect 20036 42712 20042 42724
rect 20441 42721 20453 42724
rect 20487 42721 20499 42755
rect 20441 42715 20499 42721
rect 47581 42755 47639 42761
rect 47581 42721 47593 42755
rect 47627 42721 47639 42755
rect 47581 42715 47639 42721
rect 3789 42687 3847 42693
rect 3789 42653 3801 42687
rect 3835 42684 3847 42687
rect 6840 42684 6868 42712
rect 3835 42656 6868 42684
rect 3835 42653 3847 42656
rect 3789 42647 3847 42653
rect 9674 42644 9680 42696
rect 9732 42684 9738 42696
rect 10229 42687 10287 42693
rect 10229 42684 10241 42687
rect 9732 42656 10241 42684
rect 9732 42644 9738 42656
rect 10229 42653 10241 42656
rect 10275 42684 10287 42687
rect 11330 42684 11336 42696
rect 10275 42656 11336 42684
rect 10275 42653 10287 42656
rect 10229 42647 10287 42653
rect 11330 42644 11336 42656
rect 11388 42644 11394 42696
rect 15286 42644 15292 42696
rect 15344 42684 15350 42696
rect 15473 42687 15531 42693
rect 15473 42684 15485 42687
rect 15344 42656 15485 42684
rect 15344 42644 15350 42656
rect 15473 42653 15485 42656
rect 15519 42653 15531 42687
rect 15473 42647 15531 42653
rect 17580 42687 17638 42693
rect 17580 42653 17592 42687
rect 17626 42684 17638 42687
rect 18598 42684 18604 42696
rect 17626 42656 18604 42684
rect 17626 42653 17638 42656
rect 17580 42647 17638 42653
rect 18598 42644 18604 42656
rect 18656 42644 18662 42696
rect 20456 42684 20484 42715
rect 49418 42712 49424 42764
rect 49476 42752 49482 42764
rect 50157 42755 50215 42761
rect 50157 42752 50169 42755
rect 49476 42724 50169 42752
rect 49476 42712 49482 42724
rect 50157 42721 50169 42724
rect 50203 42721 50215 42755
rect 50157 42715 50215 42721
rect 53282 42712 53288 42764
rect 53340 42752 53346 42764
rect 53377 42755 53435 42761
rect 53377 42752 53389 42755
rect 53340 42724 53389 42752
rect 53340 42712 53346 42724
rect 53377 42721 53389 42724
rect 53423 42721 53435 42755
rect 53377 42715 53435 42721
rect 56502 42712 56508 42764
rect 56560 42752 56566 42764
rect 56781 42755 56839 42761
rect 56781 42752 56793 42755
rect 56560 42724 56793 42752
rect 56560 42712 56566 42724
rect 56781 42721 56793 42724
rect 56827 42721 56839 42755
rect 56781 42715 56839 42721
rect 21542 42684 21548 42696
rect 20456 42656 21548 42684
rect 21542 42644 21548 42656
rect 21600 42684 21606 42696
rect 22002 42684 22008 42696
rect 21600 42656 22008 42684
rect 21600 42644 21606 42656
rect 22002 42644 22008 42656
rect 22060 42684 22066 42696
rect 22281 42687 22339 42693
rect 22281 42684 22293 42687
rect 22060 42656 22293 42684
rect 22060 42644 22066 42656
rect 22281 42653 22293 42656
rect 22327 42653 22339 42687
rect 22281 42647 22339 42653
rect 24397 42687 24455 42693
rect 24397 42653 24409 42687
rect 24443 42653 24455 42687
rect 24397 42647 24455 42653
rect 24664 42687 24722 42693
rect 24664 42653 24676 42687
rect 24710 42684 24722 42687
rect 26418 42684 26424 42696
rect 24710 42656 26424 42684
rect 24710 42653 24722 42656
rect 24664 42647 24722 42653
rect 4056 42619 4114 42625
rect 4056 42585 4068 42619
rect 4102 42616 4114 42619
rect 5166 42616 5172 42628
rect 4102 42588 5172 42616
rect 4102 42585 4114 42588
rect 4056 42579 4114 42585
rect 5166 42576 5172 42588
rect 5224 42576 5230 42628
rect 7276 42619 7334 42625
rect 7276 42585 7288 42619
rect 7322 42616 7334 42619
rect 8294 42616 8300 42628
rect 7322 42588 8300 42616
rect 7322 42585 7334 42588
rect 7276 42579 7334 42585
rect 8294 42576 8300 42588
rect 8352 42576 8358 42628
rect 15740 42619 15798 42625
rect 15740 42585 15752 42619
rect 15786 42616 15798 42619
rect 16022 42616 16028 42628
rect 15786 42588 16028 42616
rect 15786 42585 15798 42588
rect 15740 42579 15798 42585
rect 16022 42576 16028 42588
rect 16080 42576 16086 42628
rect 20708 42619 20766 42625
rect 20708 42585 20720 42619
rect 20754 42616 20766 42619
rect 21266 42616 21272 42628
rect 20754 42588 21272 42616
rect 20754 42585 20766 42588
rect 20708 42579 20766 42585
rect 21266 42576 21272 42588
rect 21324 42576 21330 42628
rect 22526 42619 22584 42625
rect 22526 42616 22538 42619
rect 21836 42588 22538 42616
rect 7650 42508 7656 42560
rect 7708 42548 7714 42560
rect 8389 42551 8447 42557
rect 8389 42548 8401 42551
rect 7708 42520 8401 42548
rect 7708 42508 7714 42520
rect 8389 42517 8401 42520
rect 8435 42517 8447 42551
rect 16850 42548 16856 42560
rect 16811 42520 16856 42548
rect 8389 42511 8447 42517
rect 16850 42508 16856 42520
rect 16908 42508 16914 42560
rect 18690 42548 18696 42560
rect 18651 42520 18696 42548
rect 18690 42508 18696 42520
rect 18748 42508 18754 42560
rect 21836 42557 21864 42588
rect 22526 42585 22538 42588
rect 22572 42585 22584 42619
rect 22526 42579 22584 42585
rect 22646 42576 22652 42628
rect 22704 42616 22710 42628
rect 24412 42616 24440 42647
rect 26418 42644 26424 42656
rect 26476 42644 26482 42696
rect 30837 42687 30895 42693
rect 30837 42653 30849 42687
rect 30883 42653 30895 42687
rect 30837 42647 30895 42653
rect 31104 42687 31162 42693
rect 31104 42653 31116 42687
rect 31150 42684 31162 42687
rect 31570 42684 31576 42696
rect 31150 42656 31576 42684
rect 31150 42653 31162 42656
rect 31104 42647 31162 42653
rect 22704 42588 24440 42616
rect 27249 42619 27307 42625
rect 22704 42576 22710 42588
rect 27249 42585 27261 42619
rect 27295 42616 27307 42619
rect 27338 42616 27344 42628
rect 27295 42588 27344 42616
rect 27295 42585 27307 42588
rect 27249 42579 27307 42585
rect 27338 42576 27344 42588
rect 27396 42576 27402 42628
rect 30852 42616 30880 42647
rect 31570 42644 31576 42656
rect 31628 42644 31634 42696
rect 32677 42687 32735 42693
rect 32677 42653 32689 42687
rect 32723 42684 32735 42687
rect 32766 42684 32772 42696
rect 32723 42656 32772 42684
rect 32723 42653 32735 42656
rect 32677 42647 32735 42653
rect 32766 42644 32772 42656
rect 32824 42644 32830 42696
rect 32944 42687 33002 42693
rect 32944 42653 32956 42687
rect 32990 42684 33002 42687
rect 34146 42684 34152 42696
rect 32990 42656 34152 42684
rect 32990 42653 33002 42656
rect 32944 42647 33002 42653
rect 34146 42644 34152 42656
rect 34204 42644 34210 42696
rect 35345 42687 35403 42693
rect 35345 42653 35357 42687
rect 35391 42653 35403 42687
rect 35345 42647 35403 42653
rect 35612 42687 35670 42693
rect 35612 42653 35624 42687
rect 35658 42684 35670 42687
rect 36354 42684 36360 42696
rect 35658 42656 36360 42684
rect 35658 42653 35670 42656
rect 35612 42647 35670 42653
rect 32122 42616 32128 42628
rect 30852 42588 32128 42616
rect 32122 42576 32128 42588
rect 32180 42576 32186 42628
rect 32784 42616 32812 42644
rect 34698 42616 34704 42628
rect 32784 42588 34704 42616
rect 34698 42576 34704 42588
rect 34756 42616 34762 42628
rect 35360 42616 35388 42647
rect 36354 42644 36360 42656
rect 36412 42644 36418 42696
rect 37366 42644 37372 42696
rect 37424 42684 37430 42696
rect 37826 42684 37832 42696
rect 37424 42656 37832 42684
rect 37424 42644 37430 42656
rect 37826 42644 37832 42656
rect 37884 42684 37890 42696
rect 37921 42687 37979 42693
rect 37921 42684 37933 42687
rect 37884 42656 37933 42684
rect 37884 42644 37890 42656
rect 37921 42653 37933 42656
rect 37967 42653 37979 42687
rect 37921 42647 37979 42653
rect 38188 42687 38246 42693
rect 38188 42653 38200 42687
rect 38234 42684 38246 42687
rect 40034 42684 40040 42696
rect 38234 42656 40040 42684
rect 38234 42653 38246 42656
rect 38188 42647 38246 42653
rect 40034 42644 40040 42656
rect 40092 42644 40098 42696
rect 40402 42644 40408 42696
rect 40460 42684 40466 42696
rect 40770 42693 40776 42696
rect 40497 42687 40555 42693
rect 40497 42684 40509 42687
rect 40460 42656 40509 42684
rect 40460 42644 40466 42656
rect 40497 42653 40509 42656
rect 40543 42653 40555 42687
rect 40764 42684 40776 42693
rect 40731 42656 40776 42684
rect 40497 42647 40555 42653
rect 40764 42647 40776 42656
rect 40512 42616 40540 42647
rect 40770 42644 40776 42647
rect 40828 42644 40834 42696
rect 42337 42687 42395 42693
rect 42337 42653 42349 42687
rect 42383 42684 42395 42687
rect 42426 42684 42432 42696
rect 42383 42656 42432 42684
rect 42383 42653 42395 42656
rect 42337 42647 42395 42653
rect 42352 42616 42380 42647
rect 42426 42644 42432 42656
rect 42484 42644 42490 42696
rect 44450 42644 44456 42696
rect 44508 42684 44514 42696
rect 47854 42693 47860 42696
rect 45005 42687 45063 42693
rect 45005 42684 45017 42687
rect 44508 42656 45017 42684
rect 44508 42644 44514 42656
rect 45005 42653 45017 42656
rect 45051 42653 45063 42687
rect 47848 42684 47860 42693
rect 47815 42656 47860 42684
rect 45005 42647 45063 42653
rect 47848 42647 47860 42656
rect 47854 42644 47860 42647
rect 47912 42644 47918 42696
rect 50424 42687 50482 42693
rect 50424 42653 50436 42687
rect 50470 42684 50482 42687
rect 51442 42684 51448 42696
rect 50470 42656 51448 42684
rect 50470 42653 50482 42656
rect 50424 42647 50482 42653
rect 51442 42644 51448 42656
rect 51500 42644 51506 42696
rect 57048 42687 57106 42693
rect 57048 42653 57060 42687
rect 57094 42684 57106 42687
rect 57882 42684 57888 42696
rect 57094 42656 57888 42684
rect 57094 42653 57106 42656
rect 57048 42647 57106 42653
rect 57882 42644 57888 42656
rect 57940 42644 57946 42696
rect 34756 42588 35388 42616
rect 40052 42588 42380 42616
rect 42604 42619 42662 42625
rect 34756 42576 34762 42588
rect 40052 42560 40080 42588
rect 42604 42585 42616 42619
rect 42650 42616 42662 42619
rect 43806 42616 43812 42628
rect 42650 42588 43812 42616
rect 42650 42585 42662 42588
rect 42604 42579 42662 42585
rect 43806 42576 43812 42588
rect 43864 42576 43870 42628
rect 45272 42619 45330 42625
rect 45272 42585 45284 42619
rect 45318 42616 45330 42619
rect 46750 42616 46756 42628
rect 45318 42588 46756 42616
rect 45318 42585 45330 42588
rect 45272 42579 45330 42585
rect 46750 42576 46756 42588
rect 46808 42576 46814 42628
rect 53644 42619 53702 42625
rect 53644 42585 53656 42619
rect 53690 42616 53702 42619
rect 55122 42616 55128 42628
rect 53690 42588 55128 42616
rect 53690 42585 53702 42588
rect 53644 42579 53702 42585
rect 55122 42576 55128 42588
rect 55180 42576 55186 42628
rect 21821 42551 21879 42557
rect 21821 42517 21833 42551
rect 21867 42517 21879 42551
rect 25774 42548 25780 42560
rect 25735 42520 25780 42548
rect 21821 42511 21879 42517
rect 25774 42508 25780 42520
rect 25832 42508 25838 42560
rect 27706 42508 27712 42560
rect 27764 42548 27770 42560
rect 28537 42551 28595 42557
rect 28537 42548 28549 42551
rect 27764 42520 28549 42548
rect 27764 42508 27770 42520
rect 28537 42517 28549 42520
rect 28583 42517 28595 42551
rect 28537 42511 28595 42517
rect 32030 42508 32036 42560
rect 32088 42548 32094 42560
rect 32217 42551 32275 42557
rect 32217 42548 32229 42551
rect 32088 42520 32229 42548
rect 32088 42508 32094 42520
rect 32217 42517 32229 42520
rect 32263 42517 32275 42551
rect 34054 42548 34060 42560
rect 34015 42520 34060 42548
rect 32217 42511 32275 42517
rect 34054 42508 34060 42520
rect 34112 42508 34118 42560
rect 36538 42508 36544 42560
rect 36596 42548 36602 42560
rect 36725 42551 36783 42557
rect 36725 42548 36737 42551
rect 36596 42520 36737 42548
rect 36596 42508 36602 42520
rect 36725 42517 36737 42520
rect 36771 42517 36783 42551
rect 36725 42511 36783 42517
rect 39114 42508 39120 42560
rect 39172 42548 39178 42560
rect 39301 42551 39359 42557
rect 39301 42548 39313 42551
rect 39172 42520 39313 42548
rect 39172 42508 39178 42520
rect 39301 42517 39313 42520
rect 39347 42517 39359 42551
rect 39301 42511 39359 42517
rect 40034 42508 40040 42560
rect 40092 42508 40098 42560
rect 41874 42548 41880 42560
rect 41835 42520 41880 42548
rect 41874 42508 41880 42520
rect 41932 42508 41938 42560
rect 43717 42551 43775 42557
rect 43717 42517 43729 42551
rect 43763 42548 43775 42551
rect 45094 42548 45100 42560
rect 43763 42520 45100 42548
rect 43763 42517 43775 42520
rect 43717 42511 43775 42517
rect 45094 42508 45100 42520
rect 45152 42508 45158 42560
rect 48866 42508 48872 42560
rect 48924 42548 48930 42560
rect 48961 42551 49019 42557
rect 48961 42548 48973 42551
rect 48924 42520 48973 42548
rect 48924 42508 48930 42520
rect 48961 42517 48973 42520
rect 49007 42517 49019 42551
rect 48961 42511 49019 42517
rect 51350 42508 51356 42560
rect 51408 42548 51414 42560
rect 51537 42551 51595 42557
rect 51537 42548 51549 42551
rect 51408 42520 51549 42548
rect 51408 42508 51414 42520
rect 51537 42517 51549 42520
rect 51583 42517 51595 42551
rect 54754 42548 54760 42560
rect 54715 42520 54760 42548
rect 51537 42511 51595 42517
rect 54754 42508 54760 42520
rect 54812 42508 54818 42560
rect 1104 42458 59340 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 59340 42458
rect 1104 42384 59340 42406
rect 10962 42344 10968 42356
rect 10923 42316 10968 42344
rect 10962 42304 10968 42316
rect 11020 42304 11026 42356
rect 13354 42304 13360 42356
rect 13412 42344 13418 42356
rect 14277 42347 14335 42353
rect 14277 42344 14289 42347
rect 13412 42316 14289 42344
rect 13412 42304 13418 42316
rect 14277 42313 14289 42316
rect 14323 42313 14335 42347
rect 14277 42307 14335 42313
rect 18785 42347 18843 42353
rect 18785 42313 18797 42347
rect 18831 42344 18843 42347
rect 19334 42344 19340 42356
rect 18831 42316 19340 42344
rect 18831 42313 18843 42316
rect 18785 42307 18843 42313
rect 19334 42304 19340 42316
rect 19392 42304 19398 42356
rect 21266 42344 21272 42356
rect 21227 42316 21272 42344
rect 21266 42304 21272 42316
rect 21324 42304 21330 42356
rect 24029 42347 24087 42353
rect 24029 42313 24041 42347
rect 24075 42344 24087 42347
rect 24946 42344 24952 42356
rect 24075 42316 24952 42344
rect 24075 42313 24087 42316
rect 24029 42307 24087 42313
rect 24946 42304 24952 42316
rect 25004 42304 25010 42356
rect 28902 42304 28908 42356
rect 28960 42344 28966 42356
rect 29089 42347 29147 42353
rect 29089 42344 29101 42347
rect 28960 42316 29101 42344
rect 28960 42304 28966 42316
rect 29089 42313 29101 42316
rect 29135 42313 29147 42347
rect 44450 42344 44456 42356
rect 44411 42316 44456 42344
rect 29089 42307 29147 42313
rect 44450 42304 44456 42316
rect 44508 42304 44514 42356
rect 46750 42344 46756 42356
rect 46711 42316 46756 42344
rect 46750 42304 46756 42316
rect 46808 42304 46814 42356
rect 55122 42344 55128 42356
rect 55083 42316 55128 42344
rect 55122 42304 55128 42316
rect 55180 42304 55186 42356
rect 56502 42304 56508 42356
rect 56560 42344 56566 42356
rect 56873 42347 56931 42353
rect 56873 42344 56885 42347
rect 56560 42316 56885 42344
rect 56560 42304 56566 42316
rect 56873 42313 56885 42316
rect 56919 42313 56931 42347
rect 56873 42307 56931 42313
rect 7460 42279 7518 42285
rect 7460 42245 7472 42279
rect 7506 42276 7518 42279
rect 12802 42276 12808 42288
rect 7506 42248 12808 42276
rect 7506 42245 7518 42248
rect 7460 42239 7518 42245
rect 12802 42236 12808 42248
rect 12860 42236 12866 42288
rect 13164 42279 13222 42285
rect 13164 42245 13176 42279
rect 13210 42276 13222 42279
rect 13538 42276 13544 42288
rect 13210 42248 13544 42276
rect 13210 42245 13222 42248
rect 13164 42239 13222 42245
rect 13538 42236 13544 42248
rect 13596 42236 13602 42288
rect 17672 42279 17730 42285
rect 17672 42245 17684 42279
rect 17718 42276 17730 42279
rect 18690 42276 18696 42288
rect 17718 42248 18696 42276
rect 17718 42245 17730 42248
rect 17672 42239 17730 42245
rect 18690 42236 18696 42248
rect 18748 42236 18754 42288
rect 22916 42279 22974 42285
rect 22916 42245 22928 42279
rect 22962 42276 22974 42279
rect 25682 42276 25688 42288
rect 22962 42248 25688 42276
rect 22962 42245 22974 42248
rect 22916 42239 22974 42245
rect 25682 42236 25688 42248
rect 25740 42236 25746 42288
rect 51626 42276 51632 42288
rect 50816 42248 51632 42276
rect 3136 42211 3194 42217
rect 3136 42177 3148 42211
rect 3182 42208 3194 42211
rect 5442 42208 5448 42220
rect 3182 42180 5448 42208
rect 3182 42177 3194 42180
rect 3136 42171 3194 42177
rect 5442 42168 5448 42180
rect 5500 42168 5506 42220
rect 6822 42168 6828 42220
rect 6880 42208 6886 42220
rect 7193 42211 7251 42217
rect 7193 42208 7205 42211
rect 6880 42180 7205 42208
rect 6880 42168 6886 42180
rect 7193 42177 7205 42180
rect 7239 42177 7251 42211
rect 7193 42171 7251 42177
rect 9852 42211 9910 42217
rect 9852 42177 9864 42211
rect 9898 42208 9910 42211
rect 11606 42208 11612 42220
rect 9898 42180 11612 42208
rect 9898 42177 9910 42180
rect 9852 42171 9910 42177
rect 11606 42168 11612 42180
rect 11664 42168 11670 42220
rect 12897 42211 12955 42217
rect 12897 42177 12909 42211
rect 12943 42208 12955 42211
rect 14090 42208 14096 42220
rect 12943 42180 14096 42208
rect 12943 42177 12955 42180
rect 12897 42171 12955 42177
rect 14090 42168 14096 42180
rect 14148 42208 14154 42220
rect 14737 42211 14795 42217
rect 14737 42208 14749 42211
rect 14148 42180 14749 42208
rect 14148 42168 14154 42180
rect 14737 42177 14749 42180
rect 14783 42177 14795 42211
rect 14737 42171 14795 42177
rect 15004 42211 15062 42217
rect 15004 42177 15016 42211
rect 15050 42208 15062 42211
rect 18598 42208 18604 42220
rect 15050 42180 18604 42208
rect 15050 42177 15062 42180
rect 15004 42171 15062 42177
rect 18598 42168 18604 42180
rect 18656 42168 18662 42220
rect 19889 42211 19947 42217
rect 19889 42177 19901 42211
rect 19935 42208 19947 42211
rect 19978 42208 19984 42220
rect 19935 42180 19984 42208
rect 19935 42177 19947 42180
rect 19889 42171 19947 42177
rect 19978 42168 19984 42180
rect 20036 42168 20042 42220
rect 20156 42211 20214 42217
rect 20156 42177 20168 42211
rect 20202 42208 20214 42211
rect 21542 42208 21548 42220
rect 20202 42180 21548 42208
rect 20202 42177 20214 42180
rect 20156 42171 20214 42177
rect 21542 42168 21548 42180
rect 21600 42168 21606 42220
rect 22646 42208 22652 42220
rect 22607 42180 22652 42208
rect 22646 42168 22652 42180
rect 22704 42208 22710 42220
rect 24489 42211 24547 42217
rect 24489 42208 24501 42211
rect 22704 42180 24501 42208
rect 22704 42168 22710 42180
rect 24489 42177 24501 42180
rect 24535 42177 24547 42211
rect 24489 42171 24547 42177
rect 24756 42211 24814 42217
rect 24756 42177 24768 42211
rect 24802 42208 24814 42211
rect 26142 42208 26148 42220
rect 24802 42180 26148 42208
rect 24802 42177 24814 42180
rect 24756 42171 24814 42177
rect 26142 42168 26148 42180
rect 26200 42168 26206 42220
rect 27976 42211 28034 42217
rect 27976 42177 27988 42211
rect 28022 42208 28034 42211
rect 28994 42208 29000 42220
rect 28022 42180 29000 42208
rect 28022 42177 28034 42180
rect 27976 42171 28034 42177
rect 28994 42168 29000 42180
rect 29052 42168 29058 42220
rect 34238 42168 34244 42220
rect 34296 42208 34302 42220
rect 34957 42211 35015 42217
rect 34957 42208 34969 42211
rect 34296 42180 34969 42208
rect 34296 42168 34302 42180
rect 34957 42177 34969 42180
rect 35003 42177 35015 42211
rect 34957 42171 35015 42177
rect 37826 42168 37832 42220
rect 37884 42208 37890 42220
rect 38749 42211 38807 42217
rect 38749 42208 38761 42211
rect 37884 42180 38761 42208
rect 37884 42168 37890 42180
rect 38749 42177 38761 42180
rect 38795 42177 38807 42211
rect 38749 42171 38807 42177
rect 39016 42211 39074 42217
rect 39016 42177 39028 42211
rect 39062 42208 39074 42211
rect 40218 42208 40224 42220
rect 39062 42180 40224 42208
rect 39062 42177 39074 42180
rect 39016 42171 39074 42177
rect 40218 42168 40224 42180
rect 40276 42168 40282 42220
rect 40402 42168 40408 42220
rect 40460 42208 40466 42220
rect 43165 42211 43223 42217
rect 43165 42208 43177 42211
rect 40460 42180 43177 42208
rect 40460 42168 40466 42180
rect 43165 42177 43177 42180
rect 43211 42177 43223 42211
rect 43165 42171 43223 42177
rect 45186 42168 45192 42220
rect 45244 42208 45250 42220
rect 45373 42211 45431 42217
rect 45373 42208 45385 42211
rect 45244 42180 45385 42208
rect 45244 42168 45250 42180
rect 45373 42177 45385 42180
rect 45419 42177 45431 42211
rect 45373 42171 45431 42177
rect 45640 42211 45698 42217
rect 45640 42177 45652 42211
rect 45686 42208 45698 42211
rect 46382 42208 46388 42220
rect 45686 42180 46388 42208
rect 45686 42177 45698 42180
rect 45640 42171 45698 42177
rect 46382 42168 46388 42180
rect 46440 42168 46446 42220
rect 48314 42168 48320 42220
rect 48372 42208 48378 42220
rect 48961 42211 49019 42217
rect 48961 42208 48973 42211
rect 48372 42180 48973 42208
rect 48372 42168 48378 42180
rect 48961 42177 48973 42180
rect 49007 42177 49019 42211
rect 48961 42171 49019 42177
rect 49228 42211 49286 42217
rect 49228 42177 49240 42211
rect 49274 42208 49286 42211
rect 50154 42208 50160 42220
rect 49274 42180 50160 42208
rect 49274 42177 49286 42180
rect 49228 42171 49286 42177
rect 50154 42168 50160 42180
rect 50212 42168 50218 42220
rect 50816 42217 50844 42248
rect 51626 42236 51632 42248
rect 51684 42236 51690 42288
rect 55582 42276 55588 42288
rect 55543 42248 55588 42276
rect 55582 42236 55588 42248
rect 55640 42236 55646 42288
rect 50801 42211 50859 42217
rect 50801 42177 50813 42211
rect 50847 42177 50859 42211
rect 50801 42171 50859 42177
rect 51068 42211 51126 42217
rect 51068 42177 51080 42211
rect 51114 42208 51126 42211
rect 53650 42208 53656 42220
rect 51114 42180 53656 42208
rect 51114 42177 51126 42180
rect 51068 42171 51126 42177
rect 53650 42168 53656 42180
rect 53708 42168 53714 42220
rect 54012 42211 54070 42217
rect 54012 42177 54024 42211
rect 54058 42208 54070 42211
rect 56226 42208 56232 42220
rect 54058 42180 56232 42208
rect 54058 42177 54070 42180
rect 54012 42171 54070 42177
rect 56226 42168 56232 42180
rect 56284 42168 56290 42220
rect 2869 42143 2927 42149
rect 2869 42109 2881 42143
rect 2915 42109 2927 42143
rect 2869 42103 2927 42109
rect 2884 42004 2912 42103
rect 8938 42100 8944 42152
rect 8996 42140 9002 42152
rect 9582 42140 9588 42152
rect 8996 42112 9588 42140
rect 8996 42100 9002 42112
rect 9582 42100 9588 42112
rect 9640 42100 9646 42152
rect 17310 42100 17316 42152
rect 17368 42140 17374 42152
rect 17405 42143 17463 42149
rect 17405 42140 17417 42143
rect 17368 42112 17417 42140
rect 17368 42100 17374 42112
rect 17405 42109 17417 42112
rect 17451 42109 17463 42143
rect 27706 42140 27712 42152
rect 27667 42112 27712 42140
rect 17405 42103 17463 42109
rect 27706 42100 27712 42112
rect 27764 42100 27770 42152
rect 34698 42140 34704 42152
rect 34659 42112 34704 42140
rect 34698 42100 34704 42112
rect 34756 42100 34762 42152
rect 53374 42100 53380 42152
rect 53432 42140 53438 42152
rect 53745 42143 53803 42149
rect 53745 42140 53757 42143
rect 53432 42112 53757 42140
rect 53432 42100 53438 42112
rect 53745 42109 53757 42112
rect 53791 42109 53803 42143
rect 53745 42103 53803 42109
rect 3786 42004 3792 42016
rect 2884 41976 3792 42004
rect 3786 41964 3792 41976
rect 3844 41964 3850 42016
rect 4062 41964 4068 42016
rect 4120 42004 4126 42016
rect 4249 42007 4307 42013
rect 4249 42004 4261 42007
rect 4120 41976 4261 42004
rect 4120 41964 4126 41976
rect 4249 41973 4261 41976
rect 4295 41973 4307 42007
rect 8570 42004 8576 42016
rect 8531 41976 8576 42004
rect 4249 41967 4307 41973
rect 8570 41964 8576 41976
rect 8628 41964 8634 42016
rect 16114 42004 16120 42016
rect 16075 41976 16120 42004
rect 16114 41964 16120 41976
rect 16172 41964 16178 42016
rect 25866 42004 25872 42016
rect 25827 41976 25872 42004
rect 25866 41964 25872 41976
rect 25924 41964 25930 42016
rect 36078 42004 36084 42016
rect 36039 41976 36084 42004
rect 36078 41964 36084 41976
rect 36136 41964 36142 42016
rect 40129 42007 40187 42013
rect 40129 41973 40141 42007
rect 40175 42004 40187 42007
rect 40310 42004 40316 42016
rect 40175 41976 40316 42004
rect 40175 41973 40187 41976
rect 40129 41967 40187 41973
rect 40310 41964 40316 41976
rect 40368 41964 40374 42016
rect 49694 41964 49700 42016
rect 49752 42004 49758 42016
rect 50341 42007 50399 42013
rect 50341 42004 50353 42007
rect 49752 41976 50353 42004
rect 49752 41964 49758 41976
rect 50341 41973 50353 41976
rect 50387 41973 50399 42007
rect 52178 42004 52184 42016
rect 52139 41976 52184 42004
rect 50341 41967 50399 41973
rect 52178 41964 52184 41976
rect 52236 41964 52242 42016
rect 1104 41914 59340 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 59340 41914
rect 1104 41840 59340 41862
rect 5166 41800 5172 41812
rect 5127 41772 5172 41800
rect 5166 41760 5172 41772
rect 5224 41760 5230 41812
rect 8294 41760 8300 41812
rect 8352 41800 8358 41812
rect 8389 41803 8447 41809
rect 8389 41800 8401 41803
rect 8352 41772 8401 41800
rect 8352 41760 8358 41772
rect 8389 41769 8401 41772
rect 8435 41769 8447 41803
rect 11606 41800 11612 41812
rect 11567 41772 11612 41800
rect 8389 41763 8447 41769
rect 11606 41760 11612 41772
rect 11664 41760 11670 41812
rect 21542 41800 21548 41812
rect 12084 41772 14504 41800
rect 21503 41772 21548 41800
rect 11330 41692 11336 41744
rect 11388 41732 11394 41744
rect 12084 41732 12112 41772
rect 11388 41704 12112 41732
rect 11388 41692 11394 41704
rect 6822 41624 6828 41676
rect 6880 41664 6886 41676
rect 7009 41667 7067 41673
rect 7009 41664 7021 41667
rect 6880 41636 7021 41664
rect 6880 41624 6886 41636
rect 7009 41633 7021 41636
rect 7055 41633 7067 41667
rect 7009 41627 7067 41633
rect 11422 41624 11428 41676
rect 11480 41664 11486 41676
rect 12069 41667 12127 41673
rect 12069 41664 12081 41667
rect 11480 41636 12081 41664
rect 11480 41624 11486 41636
rect 12069 41633 12081 41636
rect 12115 41633 12127 41667
rect 12069 41627 12127 41633
rect 3786 41596 3792 41608
rect 3747 41568 3792 41596
rect 3786 41556 3792 41568
rect 3844 41556 3850 41608
rect 4062 41605 4068 41608
rect 4056 41596 4068 41605
rect 4023 41568 4068 41596
rect 4056 41559 4068 41568
rect 4062 41556 4068 41559
rect 4120 41556 4126 41608
rect 7276 41599 7334 41605
rect 7276 41565 7288 41599
rect 7322 41596 7334 41599
rect 8570 41596 8576 41608
rect 7322 41568 8576 41596
rect 7322 41565 7334 41568
rect 7276 41559 7334 41565
rect 8570 41556 8576 41568
rect 8628 41556 8634 41608
rect 10229 41599 10287 41605
rect 10229 41565 10241 41599
rect 10275 41596 10287 41599
rect 12336 41599 12394 41605
rect 10275 41568 10456 41596
rect 10275 41565 10287 41568
rect 10229 41559 10287 41565
rect 10428 41460 10456 41568
rect 12336 41565 12348 41599
rect 12382 41596 12394 41599
rect 12618 41596 12624 41608
rect 12382 41568 12624 41596
rect 12382 41565 12394 41568
rect 12336 41559 12394 41565
rect 12618 41556 12624 41568
rect 12676 41556 12682 41608
rect 14476 41605 14504 41772
rect 21542 41760 21548 41772
rect 21600 41760 21606 41812
rect 28994 41800 29000 41812
rect 28955 41772 29000 41800
rect 28994 41760 29000 41772
rect 29052 41760 29058 41812
rect 41782 41760 41788 41812
rect 41840 41800 41846 41812
rect 41877 41803 41935 41809
rect 41877 41800 41889 41803
rect 41840 41772 41889 41800
rect 41840 41760 41846 41772
rect 41877 41769 41889 41772
rect 41923 41769 41935 41803
rect 43806 41800 43812 41812
rect 43767 41772 43812 41800
rect 41877 41763 41935 41769
rect 43806 41760 43812 41772
rect 43864 41760 43870 41812
rect 45186 41800 45192 41812
rect 45020 41772 45192 41800
rect 19978 41624 19984 41676
rect 20036 41664 20042 41676
rect 20165 41667 20223 41673
rect 20165 41664 20177 41667
rect 20036 41636 20177 41664
rect 20036 41624 20042 41636
rect 20165 41633 20177 41636
rect 20211 41633 20223 41667
rect 20165 41627 20223 41633
rect 22002 41624 22008 41676
rect 22060 41664 22066 41676
rect 22465 41667 22523 41673
rect 22465 41664 22477 41667
rect 22060 41636 22477 41664
rect 22060 41624 22066 41636
rect 22465 41633 22477 41636
rect 22511 41633 22523 41667
rect 22465 41627 22523 41633
rect 34698 41624 34704 41676
rect 34756 41664 34762 41676
rect 35342 41664 35348 41676
rect 34756 41636 35348 41664
rect 34756 41624 34762 41636
rect 35342 41624 35348 41636
rect 35400 41624 35406 41676
rect 45020 41673 45048 41772
rect 45186 41760 45192 41772
rect 45244 41760 45250 41812
rect 46382 41800 46388 41812
rect 46343 41772 46388 41800
rect 46382 41760 46388 41772
rect 46440 41760 46446 41812
rect 45005 41667 45063 41673
rect 45005 41633 45017 41667
rect 45051 41633 45063 41667
rect 45005 41627 45063 41633
rect 14461 41599 14519 41605
rect 14461 41565 14473 41599
rect 14507 41565 14519 41599
rect 17310 41596 17316 41608
rect 17271 41568 17316 41596
rect 14461 41559 14519 41565
rect 17310 41556 17316 41568
rect 17368 41556 17374 41608
rect 17580 41599 17638 41605
rect 17580 41565 17592 41599
rect 17626 41596 17638 41599
rect 18782 41596 18788 41608
rect 17626 41568 18788 41596
rect 17626 41565 17638 41568
rect 17580 41559 17638 41565
rect 18782 41556 18788 41568
rect 18840 41556 18846 41608
rect 24946 41556 24952 41608
rect 25004 41596 25010 41608
rect 25777 41599 25835 41605
rect 25777 41596 25789 41599
rect 25004 41568 25789 41596
rect 25004 41556 25010 41568
rect 25777 41565 25789 41568
rect 25823 41565 25835 41599
rect 25777 41559 25835 41565
rect 26044 41599 26102 41605
rect 26044 41565 26056 41599
rect 26090 41596 26102 41599
rect 27430 41596 27436 41608
rect 26090 41568 27436 41596
rect 26090 41565 26102 41568
rect 26044 41559 26102 41565
rect 10496 41531 10554 41537
rect 10496 41497 10508 41531
rect 10542 41528 10554 41531
rect 20432 41531 20490 41537
rect 10542 41500 13492 41528
rect 10542 41497 10554 41500
rect 10496 41491 10554 41497
rect 12158 41460 12164 41472
rect 10428 41432 12164 41460
rect 12158 41420 12164 41432
rect 12216 41420 12222 41472
rect 13464 41469 13492 41500
rect 20432 41497 20444 41531
rect 20478 41528 20490 41531
rect 21266 41528 21272 41540
rect 20478 41500 21272 41528
rect 20478 41497 20490 41500
rect 20432 41491 20490 41497
rect 21266 41488 21272 41500
rect 21324 41488 21330 41540
rect 22732 41531 22790 41537
rect 22732 41497 22744 41531
rect 22778 41528 22790 41531
rect 23750 41528 23756 41540
rect 22778 41500 23756 41528
rect 22778 41497 22790 41500
rect 22732 41491 22790 41497
rect 23750 41488 23756 41500
rect 23808 41488 23814 41540
rect 25792 41528 25820 41559
rect 27430 41556 27436 41568
rect 27488 41556 27494 41608
rect 27617 41599 27675 41605
rect 27617 41565 27629 41599
rect 27663 41596 27675 41599
rect 27706 41596 27712 41608
rect 27663 41568 27712 41596
rect 27663 41565 27675 41568
rect 27617 41559 27675 41565
rect 27632 41528 27660 41559
rect 27706 41556 27712 41568
rect 27764 41556 27770 41608
rect 29549 41599 29607 41605
rect 29549 41565 29561 41599
rect 29595 41596 29607 41599
rect 30190 41596 30196 41608
rect 29595 41568 30196 41596
rect 29595 41565 29607 41568
rect 29549 41559 29607 41565
rect 30190 41556 30196 41568
rect 30248 41556 30254 41608
rect 32122 41596 32128 41608
rect 32083 41568 32128 41596
rect 32122 41556 32128 41568
rect 32180 41556 32186 41608
rect 37826 41596 37832 41608
rect 37787 41568 37832 41596
rect 37826 41556 37832 41568
rect 37884 41596 37890 41608
rect 40494 41596 40500 41608
rect 37884 41568 40500 41596
rect 37884 41556 37890 41568
rect 40494 41556 40500 41568
rect 40552 41556 40558 41608
rect 40764 41599 40822 41605
rect 40764 41565 40776 41599
rect 40810 41596 40822 41599
rect 41046 41596 41052 41608
rect 40810 41568 41052 41596
rect 40810 41565 40822 41568
rect 40764 41559 40822 41565
rect 41046 41556 41052 41568
rect 41104 41556 41110 41608
rect 42426 41596 42432 41608
rect 42387 41568 42432 41596
rect 42426 41556 42432 41568
rect 42484 41556 42490 41608
rect 47673 41599 47731 41605
rect 47673 41565 47685 41599
rect 47719 41596 47731 41599
rect 48314 41596 48320 41608
rect 47719 41568 48320 41596
rect 47719 41565 47731 41568
rect 47673 41559 47731 41565
rect 48314 41556 48320 41568
rect 48372 41556 48378 41608
rect 51074 41556 51080 41608
rect 51132 41596 51138 41608
rect 51537 41599 51595 41605
rect 51537 41596 51549 41599
rect 51132 41568 51549 41596
rect 51132 41556 51138 41568
rect 51537 41565 51549 41568
rect 51583 41596 51595 41599
rect 51626 41596 51632 41608
rect 51583 41568 51632 41596
rect 51583 41565 51595 41568
rect 51537 41559 51595 41565
rect 51626 41556 51632 41568
rect 51684 41556 51690 41608
rect 52730 41556 52736 41608
rect 52788 41596 52794 41608
rect 53374 41596 53380 41608
rect 52788 41568 53380 41596
rect 52788 41556 52794 41568
rect 53374 41556 53380 41568
rect 53432 41556 53438 41608
rect 53644 41599 53702 41605
rect 53644 41565 53656 41599
rect 53690 41596 53702 41599
rect 54754 41596 54760 41608
rect 53690 41568 54760 41596
rect 53690 41565 53702 41568
rect 53644 41559 53702 41565
rect 54754 41556 54760 41568
rect 54812 41556 54818 41608
rect 55953 41599 56011 41605
rect 55953 41565 55965 41599
rect 55999 41565 56011 41599
rect 55953 41559 56011 41565
rect 56220 41599 56278 41605
rect 56220 41565 56232 41599
rect 56266 41596 56278 41599
rect 57330 41596 57336 41608
rect 56266 41568 57336 41596
rect 56266 41565 56278 41568
rect 56220 41559 56278 41565
rect 25792 41500 27660 41528
rect 27884 41531 27942 41537
rect 27884 41497 27896 41531
rect 27930 41528 27942 41531
rect 29638 41528 29644 41540
rect 27930 41500 29644 41528
rect 27930 41497 27942 41500
rect 27884 41491 27942 41497
rect 29638 41488 29644 41500
rect 29696 41488 29702 41540
rect 29816 41531 29874 41537
rect 29816 41497 29828 41531
rect 29862 41528 29874 41531
rect 31110 41528 31116 41540
rect 29862 41500 31116 41528
rect 29862 41497 29874 41500
rect 29816 41491 29874 41497
rect 31110 41488 31116 41500
rect 31168 41488 31174 41540
rect 32398 41537 32404 41540
rect 32392 41491 32404 41537
rect 32456 41528 32462 41540
rect 35612 41531 35670 41537
rect 32456 41500 32492 41528
rect 32398 41488 32404 41491
rect 32456 41488 32462 41500
rect 35612 41497 35624 41531
rect 35658 41528 35670 41531
rect 36538 41528 36544 41540
rect 35658 41500 36544 41528
rect 35658 41497 35670 41500
rect 35612 41491 35670 41497
rect 36538 41488 36544 41500
rect 36596 41488 36602 41540
rect 38096 41531 38154 41537
rect 38096 41497 38108 41531
rect 38142 41528 38154 41531
rect 39114 41528 39120 41540
rect 38142 41500 39120 41528
rect 38142 41497 38154 41500
rect 38096 41491 38154 41497
rect 39114 41488 39120 41500
rect 39172 41488 39178 41540
rect 42696 41531 42754 41537
rect 42696 41497 42708 41531
rect 42742 41528 42754 41531
rect 43714 41528 43720 41540
rect 42742 41500 43720 41528
rect 42742 41497 42754 41500
rect 42696 41491 42754 41497
rect 43714 41488 43720 41500
rect 43772 41488 43778 41540
rect 45272 41531 45330 41537
rect 45272 41497 45284 41531
rect 45318 41528 45330 41531
rect 46566 41528 46572 41540
rect 45318 41500 46572 41528
rect 45318 41497 45330 41500
rect 45272 41491 45330 41497
rect 46566 41488 46572 41500
rect 46624 41488 46630 41540
rect 47940 41531 47998 41537
rect 47940 41497 47952 41531
rect 47986 41528 47998 41531
rect 49326 41528 49332 41540
rect 47986 41500 49332 41528
rect 47986 41497 47998 41500
rect 47940 41491 47998 41497
rect 49326 41488 49332 41500
rect 49384 41488 49390 41540
rect 51804 41531 51862 41537
rect 51804 41497 51816 41531
rect 51850 41528 51862 41531
rect 53742 41528 53748 41540
rect 51850 41500 53748 41528
rect 51850 41497 51862 41500
rect 51804 41491 51862 41497
rect 53742 41488 53748 41500
rect 53800 41488 53806 41540
rect 55674 41488 55680 41540
rect 55732 41528 55738 41540
rect 55968 41528 55996 41559
rect 57330 41556 57336 41568
rect 57388 41556 57394 41608
rect 56502 41528 56508 41540
rect 55732 41500 56508 41528
rect 55732 41488 55738 41500
rect 56502 41488 56508 41500
rect 56560 41488 56566 41540
rect 13449 41463 13507 41469
rect 13449 41429 13461 41463
rect 13495 41429 13507 41463
rect 13449 41423 13507 41429
rect 14090 41420 14096 41472
rect 14148 41460 14154 41472
rect 15749 41463 15807 41469
rect 15749 41460 15761 41463
rect 14148 41432 15761 41460
rect 14148 41420 14154 41432
rect 15749 41429 15761 41432
rect 15795 41429 15807 41463
rect 18690 41460 18696 41472
rect 18651 41432 18696 41460
rect 15749 41423 15807 41429
rect 18690 41420 18696 41432
rect 18748 41420 18754 41472
rect 23198 41420 23204 41472
rect 23256 41460 23262 41472
rect 23845 41463 23903 41469
rect 23845 41460 23857 41463
rect 23256 41432 23857 41460
rect 23256 41420 23262 41432
rect 23845 41429 23857 41432
rect 23891 41429 23903 41463
rect 23845 41423 23903 41429
rect 26602 41420 26608 41472
rect 26660 41460 26666 41472
rect 27157 41463 27215 41469
rect 27157 41460 27169 41463
rect 26660 41432 27169 41460
rect 26660 41420 26666 41432
rect 27157 41429 27169 41432
rect 27203 41429 27215 41463
rect 27157 41423 27215 41429
rect 30374 41420 30380 41472
rect 30432 41460 30438 41472
rect 30929 41463 30987 41469
rect 30929 41460 30941 41463
rect 30432 41432 30941 41460
rect 30432 41420 30438 41432
rect 30929 41429 30941 41432
rect 30975 41429 30987 41463
rect 30929 41423 30987 41429
rect 32030 41420 32036 41472
rect 32088 41460 32094 41472
rect 33505 41463 33563 41469
rect 33505 41460 33517 41463
rect 32088 41432 33517 41460
rect 32088 41420 32094 41432
rect 33505 41429 33517 41432
rect 33551 41429 33563 41463
rect 33505 41423 33563 41429
rect 36262 41420 36268 41472
rect 36320 41460 36326 41472
rect 36725 41463 36783 41469
rect 36725 41460 36737 41463
rect 36320 41432 36737 41460
rect 36320 41420 36326 41432
rect 36725 41429 36737 41432
rect 36771 41429 36783 41463
rect 36725 41423 36783 41429
rect 37734 41420 37740 41472
rect 37792 41460 37798 41472
rect 39209 41463 39267 41469
rect 39209 41460 39221 41463
rect 37792 41432 39221 41460
rect 37792 41420 37798 41432
rect 39209 41429 39221 41432
rect 39255 41429 39267 41463
rect 49050 41460 49056 41472
rect 49011 41432 49056 41460
rect 39209 41423 39267 41429
rect 49050 41420 49056 41432
rect 49108 41420 49114 41472
rect 52914 41460 52920 41472
rect 52875 41432 52920 41460
rect 52914 41420 52920 41432
rect 52972 41420 52978 41472
rect 54754 41460 54760 41472
rect 54715 41432 54760 41460
rect 54754 41420 54760 41432
rect 54812 41420 54818 41472
rect 57330 41460 57336 41472
rect 57291 41432 57336 41460
rect 57330 41420 57336 41432
rect 57388 41420 57394 41472
rect 1104 41370 59340 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 59340 41370
rect 1104 41296 59340 41318
rect 3605 41259 3663 41265
rect 3605 41225 3617 41259
rect 3651 41225 3663 41259
rect 5442 41256 5448 41268
rect 5403 41228 5448 41256
rect 3605 41219 3663 41225
rect 3620 41188 3648 41219
rect 5442 41216 5448 41228
rect 5500 41216 5506 41268
rect 21266 41256 21272 41268
rect 21227 41228 21272 41256
rect 21266 41216 21272 41228
rect 21324 41216 21330 41268
rect 29638 41256 29644 41268
rect 29599 41228 29644 41256
rect 29638 41216 29644 41228
rect 29696 41216 29702 41268
rect 36538 41216 36544 41268
rect 36596 41256 36602 41268
rect 36725 41259 36783 41265
rect 36725 41256 36737 41259
rect 36596 41228 36737 41256
rect 36596 41216 36602 41228
rect 36725 41225 36737 41228
rect 36771 41225 36783 41259
rect 36725 41219 36783 41225
rect 43714 41216 43720 41268
rect 43772 41256 43778 41268
rect 43809 41259 43867 41265
rect 43809 41256 43821 41259
rect 43772 41228 43821 41256
rect 43772 41216 43778 41228
rect 43809 41225 43821 41228
rect 43855 41225 43867 41259
rect 46566 41256 46572 41268
rect 46527 41228 46572 41256
rect 43809 41219 43867 41225
rect 46566 41216 46572 41228
rect 46624 41216 46630 41268
rect 50154 41216 50160 41268
rect 50212 41256 50218 41268
rect 50341 41259 50399 41265
rect 50341 41256 50353 41259
rect 50212 41228 50353 41256
rect 50212 41216 50218 41228
rect 50341 41225 50353 41228
rect 50387 41225 50399 41259
rect 50341 41219 50399 41225
rect 53742 41216 53748 41268
rect 53800 41256 53806 41268
rect 54389 41259 54447 41265
rect 54389 41256 54401 41259
rect 53800 41228 54401 41256
rect 53800 41216 53806 41228
rect 54389 41225 54401 41228
rect 54435 41225 54447 41259
rect 54389 41219 54447 41225
rect 4310 41191 4368 41197
rect 4310 41188 4322 41191
rect 2240 41160 3372 41188
rect 3620 41160 4322 41188
rect 2240 41129 2268 41160
rect 2225 41123 2283 41129
rect 2225 41089 2237 41123
rect 2271 41089 2283 41123
rect 2225 41083 2283 41089
rect 2492 41123 2550 41129
rect 2492 41089 2504 41123
rect 2538 41120 2550 41123
rect 3234 41120 3240 41132
rect 2538 41092 3240 41120
rect 2538 41089 2550 41092
rect 2492 41083 2550 41089
rect 3234 41080 3240 41092
rect 3292 41080 3298 41132
rect 3344 41052 3372 41160
rect 4310 41157 4322 41160
rect 4356 41157 4368 41191
rect 4310 41151 4368 41157
rect 6724 41191 6782 41197
rect 6724 41157 6736 41191
rect 6770 41188 6782 41191
rect 7650 41188 7656 41200
rect 6770 41160 7656 41188
rect 6770 41157 6782 41160
rect 6724 41151 6782 41157
rect 7650 41148 7656 41160
rect 7708 41148 7714 41200
rect 9490 41197 9496 41200
rect 9484 41188 9496 41197
rect 9451 41160 9496 41188
rect 9484 41151 9496 41160
rect 9490 41148 9496 41151
rect 9548 41148 9554 41200
rect 14090 41188 14096 41200
rect 12912 41160 14096 41188
rect 12158 41080 12164 41132
rect 12216 41120 12222 41132
rect 12912 41129 12940 41160
rect 14090 41148 14096 41160
rect 14148 41148 14154 41200
rect 15004 41191 15062 41197
rect 15004 41157 15016 41191
rect 15050 41188 15062 41191
rect 16114 41188 16120 41200
rect 15050 41160 16120 41188
rect 15050 41157 15062 41160
rect 15004 41151 15062 41157
rect 16114 41148 16120 41160
rect 16172 41148 16178 41200
rect 17948 41191 18006 41197
rect 17948 41157 17960 41191
rect 17994 41188 18006 41191
rect 18690 41188 18696 41200
rect 17994 41160 18696 41188
rect 17994 41157 18006 41160
rect 17948 41151 18006 41157
rect 18690 41148 18696 41160
rect 18748 41148 18754 41200
rect 23468 41191 23526 41197
rect 23468 41157 23480 41191
rect 23514 41188 23526 41191
rect 25866 41188 25872 41200
rect 23514 41160 25872 41188
rect 23514 41157 23526 41160
rect 23468 41151 23526 41157
rect 25866 41148 25872 41160
rect 25924 41148 25930 41200
rect 51068 41191 51126 41197
rect 51068 41157 51080 41191
rect 51114 41188 51126 41191
rect 52178 41188 52184 41200
rect 51114 41160 52184 41188
rect 51114 41157 51126 41160
rect 51068 41151 51126 41157
rect 52178 41148 52184 41160
rect 52236 41148 52242 41200
rect 53276 41191 53334 41197
rect 53276 41157 53288 41191
rect 53322 41188 53334 41191
rect 54754 41188 54760 41200
rect 53322 41160 54760 41188
rect 53322 41157 53334 41160
rect 53276 41151 53334 41157
rect 54754 41148 54760 41160
rect 54812 41148 54818 41200
rect 55944 41191 56002 41197
rect 55944 41157 55956 41191
rect 55990 41188 56002 41191
rect 57330 41188 57336 41200
rect 55990 41160 57336 41188
rect 55990 41157 56002 41160
rect 55944 41151 56002 41157
rect 57330 41148 57336 41160
rect 57388 41148 57394 41200
rect 12897 41123 12955 41129
rect 12897 41120 12909 41123
rect 12216 41092 12909 41120
rect 12216 41080 12222 41092
rect 12897 41089 12909 41092
rect 12943 41089 12955 41123
rect 12897 41083 12955 41089
rect 13164 41123 13222 41129
rect 13164 41089 13176 41123
rect 13210 41120 13222 41123
rect 14826 41120 14832 41132
rect 13210 41092 14832 41120
rect 13210 41089 13222 41092
rect 13164 41083 13222 41089
rect 14826 41080 14832 41092
rect 14884 41080 14890 41132
rect 19889 41123 19947 41129
rect 19889 41089 19901 41123
rect 19935 41120 19947 41123
rect 19978 41120 19984 41132
rect 19935 41092 19984 41120
rect 19935 41089 19947 41092
rect 19889 41083 19947 41089
rect 19978 41080 19984 41092
rect 20036 41080 20042 41132
rect 20156 41123 20214 41129
rect 20156 41089 20168 41123
rect 20202 41120 20214 41123
rect 21266 41120 21272 41132
rect 20202 41092 21272 41120
rect 20202 41089 20214 41092
rect 20156 41083 20214 41089
rect 21266 41080 21272 41092
rect 21324 41080 21330 41132
rect 22646 41080 22652 41132
rect 22704 41120 22710 41132
rect 23201 41123 23259 41129
rect 23201 41120 23213 41123
rect 22704 41092 23213 41120
rect 22704 41080 22710 41092
rect 23201 41089 23213 41092
rect 23247 41089 23259 41123
rect 23201 41083 23259 41089
rect 25308 41123 25366 41129
rect 25308 41089 25320 41123
rect 25354 41120 25366 41123
rect 27154 41120 27160 41132
rect 25354 41092 27160 41120
rect 25354 41089 25366 41092
rect 25308 41083 25366 41089
rect 27154 41080 27160 41092
rect 27212 41080 27218 41132
rect 28528 41123 28586 41129
rect 28528 41089 28540 41123
rect 28574 41120 28586 41123
rect 28994 41120 29000 41132
rect 28574 41092 29000 41120
rect 28574 41089 28586 41092
rect 28528 41083 28586 41089
rect 28994 41080 29000 41092
rect 29052 41080 29058 41132
rect 30460 41123 30518 41129
rect 30460 41089 30472 41123
rect 30506 41120 30518 41123
rect 31570 41120 31576 41132
rect 30506 41092 31576 41120
rect 30506 41089 30518 41092
rect 30460 41083 30518 41089
rect 31570 41080 31576 41092
rect 31628 41080 31634 41132
rect 32760 41123 32818 41129
rect 32760 41089 32772 41123
rect 32806 41120 32818 41123
rect 34054 41120 34060 41132
rect 32806 41092 34060 41120
rect 32806 41089 32818 41092
rect 32760 41083 32818 41089
rect 34054 41080 34060 41092
rect 34112 41080 34118 41132
rect 35342 41120 35348 41132
rect 35303 41092 35348 41120
rect 35342 41080 35348 41092
rect 35400 41080 35406 41132
rect 35612 41123 35670 41129
rect 35612 41089 35624 41123
rect 35658 41120 35670 41123
rect 36722 41120 36728 41132
rect 35658 41092 36728 41120
rect 35658 41089 35670 41092
rect 35612 41083 35670 41089
rect 36722 41080 36728 41092
rect 36780 41080 36786 41132
rect 38924 41123 38982 41129
rect 38924 41089 38936 41123
rect 38970 41120 38982 41123
rect 40586 41120 40592 41132
rect 38970 41092 40592 41120
rect 38970 41089 38982 41092
rect 38924 41083 38982 41089
rect 40586 41080 40592 41092
rect 40644 41080 40650 41132
rect 40764 41123 40822 41129
rect 40764 41089 40776 41123
rect 40810 41120 40822 41123
rect 41782 41120 41788 41132
rect 40810 41092 41788 41120
rect 40810 41089 40822 41092
rect 40764 41083 40822 41089
rect 41782 41080 41788 41092
rect 41840 41080 41846 41132
rect 42696 41123 42754 41129
rect 42696 41089 42708 41123
rect 42742 41120 42754 41123
rect 43806 41120 43812 41132
rect 42742 41092 43812 41120
rect 42742 41089 42754 41092
rect 42696 41083 42754 41089
rect 43806 41080 43812 41092
rect 43864 41080 43870 41132
rect 45186 41120 45192 41132
rect 45147 41092 45192 41120
rect 45186 41080 45192 41092
rect 45244 41080 45250 41132
rect 45456 41123 45514 41129
rect 45456 41089 45468 41123
rect 45502 41120 45514 41123
rect 46842 41120 46848 41132
rect 45502 41092 46848 41120
rect 45502 41089 45514 41092
rect 45456 41083 45514 41089
rect 46842 41080 46848 41092
rect 46900 41080 46906 41132
rect 48314 41080 48320 41132
rect 48372 41120 48378 41132
rect 48961 41123 49019 41129
rect 48961 41120 48973 41123
rect 48372 41092 48973 41120
rect 48372 41080 48378 41092
rect 48961 41089 48973 41092
rect 49007 41089 49019 41123
rect 48961 41083 49019 41089
rect 49228 41123 49286 41129
rect 49228 41089 49240 41123
rect 49274 41120 49286 41123
rect 51534 41120 51540 41132
rect 49274 41092 51540 41120
rect 49274 41089 49286 41092
rect 49228 41083 49286 41089
rect 51534 41080 51540 41092
rect 51592 41080 51598 41132
rect 55674 41120 55680 41132
rect 55635 41092 55680 41120
rect 55674 41080 55680 41092
rect 55732 41080 55738 41132
rect 3786 41052 3792 41064
rect 3344 41024 3792 41052
rect 3786 41012 3792 41024
rect 3844 41052 3850 41064
rect 4065 41055 4123 41061
rect 4065 41052 4077 41055
rect 3844 41024 4077 41052
rect 3844 41012 3850 41024
rect 4065 41021 4077 41024
rect 4111 41021 4123 41055
rect 6454 41052 6460 41064
rect 6415 41024 6460 41052
rect 4065 41015 4123 41021
rect 6454 41012 6460 41024
rect 6512 41012 6518 41064
rect 8938 41012 8944 41064
rect 8996 41052 9002 41064
rect 9217 41055 9275 41061
rect 9217 41052 9229 41055
rect 8996 41024 9229 41052
rect 8996 41012 9002 41024
rect 9217 41021 9229 41024
rect 9263 41021 9275 41055
rect 9217 41015 9275 41021
rect 14090 41012 14096 41064
rect 14148 41052 14154 41064
rect 14734 41052 14740 41064
rect 14148 41024 14740 41052
rect 14148 41012 14154 41024
rect 14734 41012 14740 41024
rect 14792 41012 14798 41064
rect 17310 41012 17316 41064
rect 17368 41052 17374 41064
rect 17681 41055 17739 41061
rect 17681 41052 17693 41055
rect 17368 41024 17693 41052
rect 17368 41012 17374 41024
rect 17681 41021 17693 41024
rect 17727 41021 17739 41055
rect 17681 41015 17739 41021
rect 24946 41012 24952 41064
rect 25004 41052 25010 41064
rect 25041 41055 25099 41061
rect 25041 41052 25053 41055
rect 25004 41024 25053 41052
rect 25004 41012 25010 41024
rect 25041 41021 25053 41024
rect 25087 41021 25099 41055
rect 25041 41015 25099 41021
rect 27706 41012 27712 41064
rect 27764 41052 27770 41064
rect 28261 41055 28319 41061
rect 28261 41052 28273 41055
rect 27764 41024 28273 41052
rect 27764 41012 27770 41024
rect 28261 41021 28273 41024
rect 28307 41021 28319 41055
rect 30190 41052 30196 41064
rect 30151 41024 30196 41052
rect 28261 41015 28319 41021
rect 30190 41012 30196 41024
rect 30248 41012 30254 41064
rect 32122 41012 32128 41064
rect 32180 41052 32186 41064
rect 32490 41052 32496 41064
rect 32180 41024 32496 41052
rect 32180 41012 32186 41024
rect 32490 41012 32496 41024
rect 32548 41012 32554 41064
rect 38657 41055 38715 41061
rect 38657 41021 38669 41055
rect 38703 41021 38715 41055
rect 38657 41015 38715 41021
rect 16022 40944 16028 40996
rect 16080 40984 16086 40996
rect 16117 40987 16175 40993
rect 16117 40984 16129 40987
rect 16080 40956 16129 40984
rect 16080 40944 16086 40956
rect 16117 40953 16129 40956
rect 16163 40953 16175 40987
rect 16117 40947 16175 40953
rect 7834 40916 7840 40928
rect 7795 40888 7840 40916
rect 7834 40876 7840 40888
rect 7892 40876 7898 40928
rect 10594 40916 10600 40928
rect 10555 40888 10600 40916
rect 10594 40876 10600 40888
rect 10652 40876 10658 40928
rect 14274 40916 14280 40928
rect 14235 40888 14280 40916
rect 14274 40876 14280 40888
rect 14332 40876 14338 40928
rect 19058 40916 19064 40928
rect 19019 40888 19064 40916
rect 19058 40876 19064 40888
rect 19116 40876 19122 40928
rect 24578 40916 24584 40928
rect 24539 40888 24584 40916
rect 24578 40876 24584 40888
rect 24636 40876 24642 40928
rect 26418 40916 26424 40928
rect 26379 40888 26424 40916
rect 26418 40876 26424 40888
rect 26476 40876 26482 40928
rect 30006 40876 30012 40928
rect 30064 40916 30070 40928
rect 31573 40919 31631 40925
rect 31573 40916 31585 40919
rect 30064 40888 31585 40916
rect 30064 40876 30070 40888
rect 31573 40885 31585 40888
rect 31619 40885 31631 40919
rect 31573 40879 31631 40885
rect 31754 40876 31760 40928
rect 31812 40916 31818 40928
rect 33873 40919 33931 40925
rect 33873 40916 33885 40919
rect 31812 40888 33885 40916
rect 31812 40876 31818 40888
rect 33873 40885 33885 40888
rect 33919 40885 33931 40919
rect 38672 40916 38700 41015
rect 39942 41012 39948 41064
rect 40000 41052 40006 41064
rect 40497 41055 40555 41061
rect 40497 41052 40509 41055
rect 40000 41024 40509 41052
rect 40000 41012 40006 41024
rect 40497 41021 40509 41024
rect 40543 41021 40555 41055
rect 42426 41052 42432 41064
rect 42387 41024 42432 41052
rect 40497 41015 40555 41021
rect 42426 41012 42432 41024
rect 42484 41012 42490 41064
rect 50801 41055 50859 41061
rect 50801 41021 50813 41055
rect 50847 41021 50859 41055
rect 50801 41015 50859 41021
rect 39390 40916 39396 40928
rect 38672 40888 39396 40916
rect 33873 40879 33931 40885
rect 39390 40876 39396 40888
rect 39448 40876 39454 40928
rect 40034 40916 40040 40928
rect 39995 40888 40040 40916
rect 40034 40876 40040 40888
rect 40092 40876 40098 40928
rect 40126 40876 40132 40928
rect 40184 40916 40190 40928
rect 41877 40919 41935 40925
rect 41877 40916 41889 40919
rect 40184 40888 41889 40916
rect 40184 40876 40190 40888
rect 41877 40885 41889 40888
rect 41923 40885 41935 40919
rect 50816 40916 50844 41015
rect 52730 41012 52736 41064
rect 52788 41052 52794 41064
rect 53009 41055 53067 41061
rect 53009 41052 53021 41055
rect 52788 41024 53021 41052
rect 52788 41012 52794 41024
rect 53009 41021 53021 41024
rect 53055 41021 53067 41055
rect 53009 41015 53067 41021
rect 51074 40916 51080 40928
rect 50816 40888 51080 40916
rect 41877 40879 41935 40885
rect 51074 40876 51080 40888
rect 51132 40876 51138 40928
rect 52178 40916 52184 40928
rect 52139 40888 52184 40916
rect 52178 40876 52184 40888
rect 52236 40876 52242 40928
rect 57054 40916 57060 40928
rect 57015 40888 57060 40916
rect 57054 40876 57060 40888
rect 57112 40876 57118 40928
rect 1104 40826 59340 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 59340 40826
rect 1104 40752 59340 40774
rect 3234 40712 3240 40724
rect 3195 40684 3240 40712
rect 3234 40672 3240 40684
rect 3292 40672 3298 40724
rect 10870 40672 10876 40724
rect 10928 40712 10934 40724
rect 10965 40715 11023 40721
rect 10965 40712 10977 40715
rect 10928 40684 10977 40712
rect 10928 40672 10934 40684
rect 10965 40681 10977 40684
rect 11011 40681 11023 40715
rect 12802 40712 12808 40724
rect 12763 40684 12808 40712
rect 10965 40675 11023 40681
rect 12802 40672 12808 40684
rect 12860 40672 12866 40724
rect 18598 40672 18604 40724
rect 18656 40712 18662 40724
rect 18693 40715 18751 40721
rect 18693 40712 18705 40715
rect 18656 40684 18705 40712
rect 18656 40672 18662 40684
rect 18693 40681 18705 40684
rect 18739 40681 18751 40715
rect 18693 40675 18751 40681
rect 23750 40672 23756 40724
rect 23808 40712 23814 40724
rect 23845 40715 23903 40721
rect 23845 40712 23857 40715
rect 23808 40684 23857 40712
rect 23808 40672 23814 40684
rect 23845 40681 23857 40684
rect 23891 40681 23903 40715
rect 27154 40712 27160 40724
rect 27115 40684 27160 40712
rect 23845 40675 23903 40681
rect 27154 40672 27160 40684
rect 27212 40672 27218 40724
rect 28994 40712 29000 40724
rect 28955 40684 29000 40712
rect 28994 40672 29000 40684
rect 29052 40672 29058 40724
rect 30190 40672 30196 40724
rect 30248 40712 30254 40724
rect 32122 40712 32128 40724
rect 30248 40684 32128 40712
rect 30248 40672 30254 40684
rect 15286 40576 15292 40588
rect 15247 40548 15292 40576
rect 15286 40536 15292 40548
rect 15344 40536 15350 40588
rect 24946 40536 24952 40588
rect 25004 40576 25010 40588
rect 30576 40585 30604 40684
rect 32122 40672 32128 40684
rect 32180 40672 32186 40724
rect 41782 40712 41788 40724
rect 41743 40684 41788 40712
rect 41782 40672 41788 40684
rect 41840 40672 41846 40724
rect 43806 40712 43812 40724
rect 43767 40684 43812 40712
rect 43806 40672 43812 40684
rect 43864 40672 43870 40724
rect 45186 40712 45192 40724
rect 45020 40684 45192 40712
rect 25777 40579 25835 40585
rect 25777 40576 25789 40579
rect 25004 40548 25789 40576
rect 25004 40536 25010 40548
rect 25777 40545 25789 40548
rect 25823 40545 25835 40579
rect 25777 40539 25835 40545
rect 30561 40579 30619 40585
rect 30561 40545 30573 40579
rect 30607 40545 30619 40579
rect 37921 40579 37979 40585
rect 37921 40576 37933 40579
rect 30561 40539 30619 40545
rect 37844 40548 37933 40576
rect 1857 40511 1915 40517
rect 1857 40477 1869 40511
rect 1903 40508 1915 40511
rect 2866 40508 2872 40520
rect 1903 40480 2872 40508
rect 1903 40477 1915 40480
rect 1857 40471 1915 40477
rect 2866 40468 2872 40480
rect 2924 40468 2930 40520
rect 5810 40468 5816 40520
rect 5868 40508 5874 40520
rect 6181 40511 6239 40517
rect 6181 40508 6193 40511
rect 5868 40480 6193 40508
rect 5868 40468 5874 40480
rect 6181 40477 6193 40480
rect 6227 40477 6239 40511
rect 6181 40471 6239 40477
rect 6448 40511 6506 40517
rect 6448 40477 6460 40511
rect 6494 40508 6506 40511
rect 7834 40508 7840 40520
rect 6494 40480 7840 40508
rect 6494 40477 6506 40480
rect 6448 40471 6506 40477
rect 7834 40468 7840 40480
rect 7892 40468 7898 40520
rect 8938 40468 8944 40520
rect 8996 40508 9002 40520
rect 9585 40511 9643 40517
rect 9585 40508 9597 40511
rect 8996 40480 9597 40508
rect 8996 40468 9002 40480
rect 9585 40477 9597 40480
rect 9631 40477 9643 40511
rect 9585 40471 9643 40477
rect 9852 40511 9910 40517
rect 9852 40477 9864 40511
rect 9898 40508 9910 40511
rect 10594 40508 10600 40520
rect 9898 40480 10600 40508
rect 9898 40477 9910 40480
rect 9852 40471 9910 40477
rect 10594 40468 10600 40480
rect 10652 40468 10658 40520
rect 11425 40511 11483 40517
rect 11425 40477 11437 40511
rect 11471 40477 11483 40511
rect 11425 40471 11483 40477
rect 2124 40443 2182 40449
rect 2124 40409 2136 40443
rect 2170 40440 2182 40443
rect 3234 40440 3240 40452
rect 2170 40412 3240 40440
rect 2170 40409 2182 40412
rect 2124 40403 2182 40409
rect 3234 40400 3240 40412
rect 3292 40400 3298 40452
rect 11440 40440 11468 40471
rect 11514 40468 11520 40520
rect 11572 40508 11578 40520
rect 11681 40511 11739 40517
rect 11681 40508 11693 40511
rect 11572 40480 11693 40508
rect 11572 40468 11578 40480
rect 11681 40477 11693 40480
rect 11727 40477 11739 40511
rect 11681 40471 11739 40477
rect 12158 40440 12164 40452
rect 11440 40412 12164 40440
rect 12158 40400 12164 40412
rect 12216 40400 12222 40452
rect 15304 40440 15332 40536
rect 15556 40511 15614 40517
rect 15556 40477 15568 40511
rect 15602 40508 15614 40511
rect 16850 40508 16856 40520
rect 15602 40480 16856 40508
rect 15602 40477 15614 40480
rect 15556 40471 15614 40477
rect 16850 40468 16856 40480
rect 16908 40468 16914 40520
rect 17310 40508 17316 40520
rect 17271 40480 17316 40508
rect 17310 40468 17316 40480
rect 17368 40468 17374 40520
rect 17580 40511 17638 40517
rect 17580 40477 17592 40511
rect 17626 40508 17638 40511
rect 19058 40508 19064 40520
rect 17626 40480 19064 40508
rect 17626 40477 17638 40480
rect 17580 40471 17638 40477
rect 19058 40468 19064 40480
rect 19116 40468 19122 40520
rect 22465 40511 22523 40517
rect 22465 40477 22477 40511
rect 22511 40508 22523 40511
rect 22554 40508 22560 40520
rect 22511 40480 22560 40508
rect 22511 40477 22523 40480
rect 22465 40471 22523 40477
rect 22554 40468 22560 40480
rect 22612 40468 22618 40520
rect 22732 40511 22790 40517
rect 22732 40477 22744 40511
rect 22778 40508 22790 40511
rect 24578 40508 24584 40520
rect 22778 40480 24584 40508
rect 22778 40477 22790 40480
rect 22732 40471 22790 40477
rect 24578 40468 24584 40480
rect 24636 40468 24642 40520
rect 26044 40511 26102 40517
rect 26044 40477 26056 40511
rect 26090 40508 26102 40511
rect 26602 40508 26608 40520
rect 26090 40480 26608 40508
rect 26090 40477 26102 40480
rect 26044 40471 26102 40477
rect 26602 40468 26608 40480
rect 26660 40468 26666 40520
rect 27617 40511 27675 40517
rect 27617 40477 27629 40511
rect 27663 40508 27675 40511
rect 27706 40508 27712 40520
rect 27663 40480 27712 40508
rect 27663 40477 27675 40480
rect 27617 40471 27675 40477
rect 27706 40468 27712 40480
rect 27764 40468 27770 40520
rect 30828 40511 30886 40517
rect 30828 40477 30840 40511
rect 30874 40508 30886 40511
rect 32030 40508 32036 40520
rect 30874 40480 32036 40508
rect 30874 40477 30886 40480
rect 30828 40471 30886 40477
rect 32030 40468 32036 40480
rect 32088 40468 32094 40520
rect 35986 40468 35992 40520
rect 36044 40508 36050 40520
rect 36081 40511 36139 40517
rect 36081 40508 36093 40511
rect 36044 40480 36093 40508
rect 36044 40468 36050 40480
rect 36081 40477 36093 40480
rect 36127 40477 36139 40511
rect 36081 40471 36139 40477
rect 36348 40511 36406 40517
rect 36348 40477 36360 40511
rect 36394 40508 36406 40511
rect 37734 40508 37740 40520
rect 36394 40480 37740 40508
rect 36394 40477 36406 40480
rect 36348 40471 36406 40477
rect 17328 40440 17356 40468
rect 15304 40412 17356 40440
rect 19613 40443 19671 40449
rect 19613 40409 19625 40443
rect 19659 40440 19671 40443
rect 20530 40440 20536 40452
rect 19659 40412 20536 40440
rect 19659 40409 19671 40412
rect 19613 40403 19671 40409
rect 20530 40400 20536 40412
rect 20588 40400 20594 40452
rect 27884 40443 27942 40449
rect 27884 40409 27896 40443
rect 27930 40440 27942 40443
rect 29730 40440 29736 40452
rect 27930 40412 29736 40440
rect 27930 40409 27942 40412
rect 27884 40403 27942 40409
rect 29730 40400 29736 40412
rect 29788 40400 29794 40452
rect 32306 40400 32312 40452
rect 32364 40440 32370 40452
rect 32401 40443 32459 40449
rect 32401 40440 32413 40443
rect 32364 40412 32413 40440
rect 32364 40400 32370 40412
rect 32401 40409 32413 40412
rect 32447 40440 32459 40443
rect 32950 40440 32956 40452
rect 32447 40412 32956 40440
rect 32447 40409 32459 40412
rect 32401 40403 32459 40409
rect 32950 40400 32956 40412
rect 33008 40400 33014 40452
rect 34149 40443 34207 40449
rect 34149 40409 34161 40443
rect 34195 40440 34207 40443
rect 34330 40440 34336 40452
rect 34195 40412 34336 40440
rect 34195 40409 34207 40412
rect 34149 40403 34207 40409
rect 34330 40400 34336 40412
rect 34388 40400 34394 40452
rect 36096 40440 36124 40471
rect 37734 40468 37740 40480
rect 37792 40468 37798 40520
rect 37844 40452 37872 40548
rect 37921 40545 37933 40548
rect 37967 40545 37979 40579
rect 37921 40539 37979 40545
rect 39390 40536 39396 40588
rect 39448 40576 39454 40588
rect 39942 40576 39948 40588
rect 39448 40548 39948 40576
rect 39448 40536 39454 40548
rect 39942 40536 39948 40548
rect 40000 40576 40006 40588
rect 45020 40585 45048 40684
rect 45186 40672 45192 40684
rect 45244 40672 45250 40724
rect 46198 40672 46204 40724
rect 46256 40712 46262 40724
rect 46385 40715 46443 40721
rect 46385 40712 46397 40715
rect 46256 40684 46397 40712
rect 46256 40672 46262 40684
rect 46385 40681 46397 40684
rect 46431 40681 46443 40715
rect 51074 40712 51080 40724
rect 46385 40675 46443 40681
rect 50448 40684 51080 40712
rect 50448 40585 50476 40684
rect 51074 40672 51080 40684
rect 51132 40672 51138 40724
rect 53650 40712 53656 40724
rect 53611 40684 53656 40712
rect 53650 40672 53656 40684
rect 53708 40672 53714 40724
rect 55674 40712 55680 40724
rect 55324 40684 55680 40712
rect 40405 40579 40463 40585
rect 40405 40576 40417 40579
rect 40000 40548 40417 40576
rect 40000 40536 40006 40548
rect 40405 40545 40417 40548
rect 40451 40545 40463 40579
rect 40405 40539 40463 40545
rect 45005 40579 45063 40585
rect 45005 40545 45017 40579
rect 45051 40545 45063 40579
rect 45005 40539 45063 40545
rect 50433 40579 50491 40585
rect 50433 40545 50445 40579
rect 50479 40545 50491 40579
rect 50433 40539 50491 40545
rect 38188 40511 38246 40517
rect 38188 40477 38200 40511
rect 38234 40508 38246 40511
rect 40034 40508 40040 40520
rect 38234 40480 40040 40508
rect 38234 40477 38246 40480
rect 38188 40471 38246 40477
rect 40034 40468 40040 40480
rect 40092 40468 40098 40520
rect 40420 40508 40448 40539
rect 51626 40536 51632 40588
rect 51684 40576 51690 40588
rect 52273 40579 52331 40585
rect 52273 40576 52285 40579
rect 51684 40548 52285 40576
rect 51684 40536 51690 40548
rect 52273 40545 52285 40548
rect 52319 40545 52331 40579
rect 52273 40539 52331 40545
rect 53374 40536 53380 40588
rect 53432 40576 53438 40588
rect 55324 40585 55352 40684
rect 55674 40672 55680 40684
rect 55732 40672 55738 40724
rect 56226 40672 56232 40724
rect 56284 40712 56290 40724
rect 56689 40715 56747 40721
rect 56689 40712 56701 40715
rect 56284 40684 56701 40712
rect 56284 40672 56290 40684
rect 56689 40681 56701 40684
rect 56735 40681 56747 40715
rect 56689 40675 56747 40681
rect 55309 40579 55367 40585
rect 55309 40576 55321 40579
rect 53432 40548 55321 40576
rect 53432 40536 53438 40548
rect 55309 40545 55321 40548
rect 55355 40545 55367 40579
rect 55309 40539 55367 40545
rect 42426 40508 42432 40520
rect 40420 40480 42432 40508
rect 42426 40468 42432 40480
rect 42484 40468 42490 40520
rect 43070 40508 43076 40520
rect 42536 40480 43076 40508
rect 37826 40440 37832 40452
rect 36096 40412 37832 40440
rect 37826 40400 37832 40412
rect 37884 40400 37890 40452
rect 40672 40443 40730 40449
rect 40672 40409 40684 40443
rect 40718 40440 40730 40443
rect 42536 40440 42564 40480
rect 43070 40468 43076 40480
rect 43128 40468 43134 40520
rect 45094 40468 45100 40520
rect 45152 40508 45158 40520
rect 45261 40511 45319 40517
rect 45261 40508 45273 40511
rect 45152 40480 45273 40508
rect 45152 40468 45158 40480
rect 45261 40477 45273 40480
rect 45307 40477 45319 40511
rect 45261 40471 45319 40477
rect 48225 40511 48283 40517
rect 48225 40477 48237 40511
rect 48271 40508 48283 40511
rect 48314 40508 48320 40520
rect 48271 40480 48320 40508
rect 48271 40477 48283 40480
rect 48225 40471 48283 40477
rect 48314 40468 48320 40480
rect 48372 40468 48378 40520
rect 48492 40511 48550 40517
rect 48492 40477 48504 40511
rect 48538 40508 48550 40511
rect 49694 40508 49700 40520
rect 48538 40480 49700 40508
rect 48538 40477 48550 40480
rect 48492 40471 48550 40477
rect 49694 40468 49700 40480
rect 49752 40468 49758 40520
rect 50700 40511 50758 40517
rect 50700 40477 50712 40511
rect 50746 40508 50758 40511
rect 52178 40508 52184 40520
rect 50746 40480 52184 40508
rect 50746 40477 50758 40480
rect 50700 40471 50758 40477
rect 52178 40468 52184 40480
rect 52236 40468 52242 40520
rect 52540 40511 52598 40517
rect 52540 40477 52552 40511
rect 52586 40508 52598 40511
rect 52914 40508 52920 40520
rect 52586 40480 52920 40508
rect 52586 40477 52598 40480
rect 52540 40471 52598 40477
rect 52914 40468 52920 40480
rect 52972 40468 52978 40520
rect 55576 40511 55634 40517
rect 55576 40477 55588 40511
rect 55622 40508 55634 40511
rect 57054 40508 57060 40520
rect 55622 40480 57060 40508
rect 55622 40477 55634 40480
rect 55576 40471 55634 40477
rect 57054 40468 57060 40480
rect 57112 40468 57118 40520
rect 40718 40412 42564 40440
rect 42696 40443 42754 40449
rect 40718 40409 40730 40412
rect 40672 40403 40730 40409
rect 42696 40409 42708 40443
rect 42742 40440 42754 40443
rect 43714 40440 43720 40452
rect 42742 40412 43720 40440
rect 42742 40409 42754 40412
rect 42696 40403 42754 40409
rect 43714 40400 43720 40412
rect 43772 40400 43778 40452
rect 7558 40372 7564 40384
rect 7519 40344 7564 40372
rect 7558 40332 7564 40344
rect 7616 40332 7622 40384
rect 15286 40332 15292 40384
rect 15344 40372 15350 40384
rect 16669 40375 16727 40381
rect 16669 40372 16681 40375
rect 15344 40344 16681 40372
rect 15344 40332 15350 40344
rect 16669 40341 16681 40344
rect 16715 40341 16727 40375
rect 21082 40372 21088 40384
rect 21043 40344 21088 40372
rect 16669 40335 16727 40341
rect 21082 40332 21088 40344
rect 21140 40332 21146 40384
rect 31938 40372 31944 40384
rect 31899 40344 31944 40372
rect 31938 40332 31944 40344
rect 31996 40332 32002 40384
rect 37458 40372 37464 40384
rect 37419 40344 37464 40372
rect 37458 40332 37464 40344
rect 37516 40332 37522 40384
rect 39298 40372 39304 40384
rect 39259 40344 39304 40372
rect 39298 40332 39304 40344
rect 39356 40332 39362 40384
rect 49602 40372 49608 40384
rect 49563 40344 49608 40372
rect 49602 40332 49608 40344
rect 49660 40332 49666 40384
rect 51810 40372 51816 40384
rect 51771 40344 51816 40372
rect 51810 40332 51816 40344
rect 51868 40332 51874 40384
rect 1104 40282 59340 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 59340 40282
rect 1104 40208 59340 40230
rect 18049 40171 18107 40177
rect 18049 40137 18061 40171
rect 18095 40168 18107 40171
rect 19334 40168 19340 40180
rect 18095 40140 19340 40168
rect 18095 40137 18107 40140
rect 18049 40131 18107 40137
rect 19334 40128 19340 40140
rect 19392 40128 19398 40180
rect 21266 40168 21272 40180
rect 21227 40140 21272 40168
rect 21266 40128 21272 40140
rect 21324 40128 21330 40180
rect 26142 40168 26148 40180
rect 26103 40140 26148 40168
rect 26142 40128 26148 40140
rect 26200 40128 26206 40180
rect 29730 40168 29736 40180
rect 29691 40140 29736 40168
rect 29730 40128 29736 40140
rect 29788 40128 29794 40180
rect 31570 40168 31576 40180
rect 31531 40140 31576 40168
rect 31570 40128 31576 40140
rect 31628 40128 31634 40180
rect 36722 40168 36728 40180
rect 36683 40140 36728 40168
rect 36722 40128 36728 40140
rect 36780 40128 36786 40180
rect 40586 40128 40592 40180
rect 40644 40168 40650 40180
rect 40773 40171 40831 40177
rect 40773 40168 40785 40171
rect 40644 40140 40785 40168
rect 40644 40128 40650 40140
rect 40773 40137 40785 40140
rect 40819 40137 40831 40171
rect 40773 40131 40831 40137
rect 43714 40128 43720 40180
rect 43772 40168 43778 40180
rect 43809 40171 43867 40177
rect 43809 40168 43821 40171
rect 43772 40140 43821 40168
rect 43772 40128 43778 40140
rect 43809 40137 43821 40140
rect 43855 40137 43867 40171
rect 51534 40168 51540 40180
rect 51495 40140 51540 40168
rect 43809 40131 43867 40137
rect 51534 40128 51540 40140
rect 51592 40128 51598 40180
rect 2866 40100 2872 40112
rect 2240 40072 2872 40100
rect 2240 40041 2268 40072
rect 2866 40060 2872 40072
rect 2924 40100 2930 40112
rect 3786 40100 3792 40112
rect 2924 40072 3792 40100
rect 2924 40060 2930 40072
rect 3786 40060 3792 40072
rect 3844 40060 3850 40112
rect 4065 40103 4123 40109
rect 4065 40069 4077 40103
rect 4111 40100 4123 40103
rect 5626 40100 5632 40112
rect 4111 40072 5632 40100
rect 4111 40069 4123 40072
rect 4065 40063 4123 40069
rect 5626 40060 5632 40072
rect 5684 40060 5690 40112
rect 17310 40100 17316 40112
rect 16684 40072 17316 40100
rect 2225 40035 2283 40041
rect 2225 40001 2237 40035
rect 2271 40001 2283 40035
rect 2225 39995 2283 40001
rect 2492 40035 2550 40041
rect 2492 40001 2504 40035
rect 2538 40032 2550 40035
rect 3970 40032 3976 40044
rect 2538 40004 3976 40032
rect 2538 40001 2550 40004
rect 2492 39995 2550 40001
rect 3970 39992 3976 40004
rect 4028 39992 4034 40044
rect 6365 40035 6423 40041
rect 6365 40001 6377 40035
rect 6411 40032 6423 40035
rect 6454 40032 6460 40044
rect 6411 40004 6460 40032
rect 6411 40001 6423 40004
rect 6365 39995 6423 40001
rect 5810 39964 5816 39976
rect 5771 39936 5816 39964
rect 5810 39924 5816 39936
rect 5868 39924 5874 39976
rect 3602 39828 3608 39840
rect 3563 39800 3608 39828
rect 3602 39788 3608 39800
rect 3660 39788 3666 39840
rect 6380 39828 6408 39995
rect 6454 39992 6460 40004
rect 6512 39992 6518 40044
rect 6632 40035 6690 40041
rect 6632 40001 6644 40035
rect 6678 40032 6690 40035
rect 7558 40032 7564 40044
rect 6678 40004 7564 40032
rect 6678 40001 6690 40004
rect 6632 39995 6690 40001
rect 7558 39992 7564 40004
rect 7616 39992 7622 40044
rect 7834 39992 7840 40044
rect 7892 40032 7898 40044
rect 8461 40035 8519 40041
rect 8461 40032 8473 40035
rect 7892 40004 8473 40032
rect 7892 39992 7898 40004
rect 8461 40001 8473 40004
rect 8507 40001 8519 40035
rect 12158 40032 12164 40044
rect 12119 40004 12164 40032
rect 8461 39995 8519 40001
rect 12158 39992 12164 40004
rect 12216 39992 12222 40044
rect 12428 40035 12486 40041
rect 12428 40001 12440 40035
rect 12474 40032 12486 40035
rect 14274 40032 14280 40044
rect 12474 40004 14280 40032
rect 12474 40001 12486 40004
rect 12428 39995 12486 40001
rect 14274 39992 14280 40004
rect 14332 39992 14338 40044
rect 14734 40032 14740 40044
rect 14695 40004 14740 40032
rect 14734 39992 14740 40004
rect 14792 39992 14798 40044
rect 15004 40035 15062 40041
rect 15004 40001 15016 40035
rect 15050 40032 15062 40035
rect 15286 40032 15292 40044
rect 15050 40004 15292 40032
rect 15050 40001 15062 40004
rect 15004 39995 15062 40001
rect 15286 39992 15292 40004
rect 15344 39992 15350 40044
rect 16684 40041 16712 40072
rect 17310 40060 17316 40072
rect 17368 40060 17374 40112
rect 24946 40060 24952 40112
rect 25004 40060 25010 40112
rect 32490 40060 32496 40112
rect 32548 40100 32554 40112
rect 34330 40100 34336 40112
rect 32548 40072 34336 40100
rect 32548 40060 32554 40072
rect 16669 40035 16727 40041
rect 16669 40001 16681 40035
rect 16715 40001 16727 40035
rect 16669 39995 16727 40001
rect 16936 40035 16994 40041
rect 16936 40001 16948 40035
rect 16982 40032 16994 40035
rect 18046 40032 18052 40044
rect 16982 40004 18052 40032
rect 16982 40001 16994 40004
rect 16936 39995 16994 40001
rect 18046 39992 18052 40004
rect 18104 39992 18110 40044
rect 19889 40035 19947 40041
rect 19889 40001 19901 40035
rect 19935 40032 19947 40035
rect 19978 40032 19984 40044
rect 19935 40004 19984 40032
rect 19935 40001 19947 40004
rect 19889 39995 19947 40001
rect 19978 39992 19984 40004
rect 20036 39992 20042 40044
rect 20156 40035 20214 40041
rect 20156 40001 20168 40035
rect 20202 40032 20214 40035
rect 23014 40032 23020 40044
rect 20202 40004 23020 40032
rect 20202 40001 20214 40004
rect 20156 39995 20214 40001
rect 23014 39992 23020 40004
rect 23072 39992 23078 40044
rect 23198 40041 23204 40044
rect 23192 40032 23204 40041
rect 23159 40004 23204 40032
rect 23192 39995 23204 40004
rect 23198 39992 23204 39995
rect 23256 39992 23262 40044
rect 24765 40035 24823 40041
rect 24765 40001 24777 40035
rect 24811 40032 24823 40035
rect 24964 40032 24992 40060
rect 32784 40044 32812 40072
rect 34330 40060 34336 40072
rect 34388 40060 34394 40112
rect 35986 40100 35992 40112
rect 35544 40072 35992 40100
rect 24811 40004 24992 40032
rect 25032 40035 25090 40041
rect 24811 40001 24823 40004
rect 24765 39995 24823 40001
rect 25032 40001 25044 40035
rect 25078 40032 25090 40035
rect 26418 40032 26424 40044
rect 25078 40004 26424 40032
rect 25078 40001 25090 40004
rect 25032 39995 25090 40001
rect 26418 39992 26424 40004
rect 26476 39992 26482 40044
rect 27706 39992 27712 40044
rect 27764 40032 27770 40044
rect 28353 40035 28411 40041
rect 28353 40032 28365 40035
rect 27764 40004 28365 40032
rect 27764 39992 27770 40004
rect 28353 40001 28365 40004
rect 28399 40001 28411 40035
rect 28353 39995 28411 40001
rect 28620 40035 28678 40041
rect 28620 40001 28632 40035
rect 28666 40032 28678 40035
rect 30282 40032 30288 40044
rect 28666 40004 30288 40032
rect 28666 40001 28678 40004
rect 28620 39995 28678 40001
rect 30282 39992 30288 40004
rect 30340 39992 30346 40044
rect 30460 40035 30518 40041
rect 30460 40001 30472 40035
rect 30506 40032 30518 40035
rect 31570 40032 31576 40044
rect 30506 40004 31576 40032
rect 30506 40001 30518 40004
rect 30460 39995 30518 40001
rect 31570 39992 31576 40004
rect 31628 39992 31634 40044
rect 32766 40032 32772 40044
rect 32679 40004 32772 40032
rect 32766 39992 32772 40004
rect 32824 39992 32830 40044
rect 33036 40035 33094 40041
rect 33036 40001 33048 40035
rect 33082 40032 33094 40035
rect 35345 40035 35403 40041
rect 33082 40004 34468 40032
rect 33082 40001 33094 40004
rect 33036 39995 33094 40001
rect 8202 39964 8208 39976
rect 7576 39936 8208 39964
rect 7576 39828 7604 39936
rect 8202 39924 8208 39936
rect 8260 39924 8266 39976
rect 22554 39924 22560 39976
rect 22612 39964 22618 39976
rect 22925 39967 22983 39973
rect 22925 39964 22937 39967
rect 22612 39936 22937 39964
rect 22612 39924 22618 39936
rect 22925 39933 22937 39936
rect 22971 39933 22983 39967
rect 30190 39964 30196 39976
rect 30151 39936 30196 39964
rect 22925 39927 22983 39933
rect 30190 39924 30196 39936
rect 30248 39924 30254 39976
rect 7742 39828 7748 39840
rect 6380 39800 7604 39828
rect 7703 39800 7748 39828
rect 7742 39788 7748 39800
rect 7800 39788 7806 39840
rect 8386 39788 8392 39840
rect 8444 39828 8450 39840
rect 9585 39831 9643 39837
rect 9585 39828 9597 39831
rect 8444 39800 9597 39828
rect 8444 39788 8450 39800
rect 9585 39797 9597 39800
rect 9631 39797 9643 39831
rect 13538 39828 13544 39840
rect 13499 39800 13544 39828
rect 9585 39791 9643 39797
rect 13538 39788 13544 39800
rect 13596 39788 13602 39840
rect 16114 39828 16120 39840
rect 16075 39800 16120 39828
rect 16114 39788 16120 39800
rect 16172 39788 16178 39840
rect 24302 39828 24308 39840
rect 24263 39800 24308 39828
rect 24302 39788 24308 39800
rect 24360 39788 24366 39840
rect 34146 39828 34152 39840
rect 34107 39800 34152 39828
rect 34146 39788 34152 39800
rect 34204 39788 34210 39840
rect 34440 39828 34468 40004
rect 35345 40001 35357 40035
rect 35391 40032 35403 40035
rect 35544 40032 35572 40072
rect 35986 40060 35992 40072
rect 36044 40060 36050 40112
rect 47946 40100 47952 40112
rect 47859 40072 47952 40100
rect 47946 40060 47952 40072
rect 48004 40100 48010 40112
rect 49786 40100 49792 40112
rect 48004 40072 49792 40100
rect 48004 40060 48010 40072
rect 49786 40060 49792 40072
rect 49844 40060 49850 40112
rect 51074 40100 51080 40112
rect 50172 40072 51080 40100
rect 35391 40004 35572 40032
rect 35612 40035 35670 40041
rect 35391 40001 35403 40004
rect 35345 39995 35403 40001
rect 35612 40001 35624 40035
rect 35658 40032 35670 40035
rect 37366 40032 37372 40044
rect 35658 40004 37372 40032
rect 35658 40001 35670 40004
rect 35612 39995 35670 40001
rect 37366 39992 37372 40004
rect 37424 39992 37430 40044
rect 37820 40035 37878 40041
rect 37820 40001 37832 40035
rect 37866 40032 37878 40035
rect 39390 40032 39396 40044
rect 37866 40004 39068 40032
rect 39351 40004 39396 40032
rect 37866 40001 37878 40004
rect 37820 39995 37878 40001
rect 37553 39967 37611 39973
rect 37553 39933 37565 39967
rect 37599 39933 37611 39967
rect 37553 39927 37611 39933
rect 36078 39828 36084 39840
rect 34440 39800 36084 39828
rect 36078 39788 36084 39800
rect 36136 39788 36142 39840
rect 37568 39828 37596 39927
rect 38746 39828 38752 39840
rect 37568 39800 38752 39828
rect 38746 39788 38752 39800
rect 38804 39788 38810 39840
rect 38930 39828 38936 39840
rect 38891 39800 38936 39828
rect 38930 39788 38936 39800
rect 38988 39788 38994 39840
rect 39040 39828 39068 40004
rect 39390 39992 39396 40004
rect 39448 39992 39454 40044
rect 39660 40035 39718 40041
rect 39660 40001 39672 40035
rect 39706 40032 39718 40035
rect 40126 40032 40132 40044
rect 39706 40004 40132 40032
rect 39706 40001 39718 40004
rect 39660 39995 39718 40001
rect 40126 39992 40132 40004
rect 40184 39992 40190 40044
rect 42426 40032 42432 40044
rect 42387 40004 42432 40032
rect 42426 39992 42432 40004
rect 42484 39992 42490 40044
rect 42696 40035 42754 40041
rect 42696 40001 42708 40035
rect 42742 40032 42754 40035
rect 43806 40032 43812 40044
rect 42742 40004 43812 40032
rect 42742 40001 42754 40004
rect 42696 39995 42754 40001
rect 43806 39992 43812 40004
rect 43864 39992 43870 40044
rect 45186 39992 45192 40044
rect 45244 40032 45250 40044
rect 45649 40035 45707 40041
rect 45649 40032 45661 40035
rect 45244 40004 45661 40032
rect 45244 39992 45250 40004
rect 45649 40001 45661 40004
rect 45695 40001 45707 40035
rect 45649 39995 45707 40001
rect 45916 40035 45974 40041
rect 45916 40001 45928 40035
rect 45962 40032 45974 40035
rect 47762 40032 47768 40044
rect 45962 40004 47768 40032
rect 45962 40001 45974 40004
rect 45916 39995 45974 40001
rect 47762 39992 47768 40004
rect 47820 39992 47826 40044
rect 50172 40041 50200 40072
rect 51074 40060 51080 40072
rect 51132 40060 51138 40112
rect 50157 40035 50215 40041
rect 50157 40001 50169 40035
rect 50203 40001 50215 40035
rect 50157 39995 50215 40001
rect 50424 40035 50482 40041
rect 50424 40001 50436 40035
rect 50470 40032 50482 40035
rect 51810 40032 51816 40044
rect 50470 40004 51816 40032
rect 50470 40001 50482 40004
rect 50424 39995 50482 40001
rect 51810 39992 51816 40004
rect 51868 39992 51874 40044
rect 40310 39828 40316 39840
rect 39040 39800 40316 39828
rect 40310 39788 40316 39800
rect 40368 39788 40374 39840
rect 47026 39828 47032 39840
rect 46987 39800 47032 39828
rect 47026 39788 47032 39800
rect 47084 39788 47090 39840
rect 48222 39788 48228 39840
rect 48280 39828 48286 39840
rect 49237 39831 49295 39837
rect 49237 39828 49249 39831
rect 48280 39800 49249 39828
rect 48280 39788 48286 39800
rect 49237 39797 49249 39800
rect 49283 39797 49295 39831
rect 49237 39791 49295 39797
rect 49786 39788 49792 39840
rect 49844 39828 49850 39840
rect 53098 39828 53104 39840
rect 49844 39800 53104 39828
rect 49844 39788 49850 39800
rect 53098 39788 53104 39800
rect 53156 39828 53162 39840
rect 54662 39828 54668 39840
rect 53156 39800 54668 39828
rect 53156 39788 53162 39800
rect 54662 39788 54668 39800
rect 54720 39788 54726 39840
rect 1104 39738 59340 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 59340 39738
rect 1104 39664 59340 39686
rect 3234 39624 3240 39636
rect 3195 39596 3240 39624
rect 3234 39584 3240 39596
rect 3292 39584 3298 39636
rect 3970 39584 3976 39636
rect 4028 39624 4034 39636
rect 5169 39627 5227 39633
rect 5169 39624 5181 39627
rect 4028 39596 5181 39624
rect 4028 39584 4034 39596
rect 5169 39593 5181 39596
rect 5215 39593 5227 39627
rect 5169 39587 5227 39593
rect 7745 39627 7803 39633
rect 7745 39593 7757 39627
rect 7791 39624 7803 39627
rect 7834 39624 7840 39636
rect 7791 39596 7840 39624
rect 7791 39593 7803 39596
rect 7745 39587 7803 39593
rect 7834 39584 7840 39596
rect 7892 39584 7898 39636
rect 11330 39584 11336 39636
rect 11388 39624 11394 39636
rect 11517 39627 11575 39633
rect 11517 39624 11529 39627
rect 11388 39596 11529 39624
rect 11388 39584 11394 39596
rect 11517 39593 11529 39596
rect 11563 39593 11575 39627
rect 18046 39624 18052 39636
rect 11517 39587 11575 39593
rect 11716 39596 17908 39624
rect 18007 39596 18052 39624
rect 8294 39448 8300 39500
rect 8352 39488 8358 39500
rect 8938 39488 8944 39500
rect 8352 39460 8944 39488
rect 8352 39448 8358 39460
rect 8938 39448 8944 39460
rect 8996 39448 9002 39500
rect 1857 39423 1915 39429
rect 1857 39389 1869 39423
rect 1903 39389 1915 39423
rect 1857 39383 1915 39389
rect 2124 39423 2182 39429
rect 2124 39389 2136 39423
rect 2170 39420 2182 39423
rect 3602 39420 3608 39432
rect 2170 39392 3608 39420
rect 2170 39389 2182 39392
rect 2124 39383 2182 39389
rect 1872 39352 1900 39383
rect 3602 39380 3608 39392
rect 3660 39380 3666 39432
rect 3786 39420 3792 39432
rect 3747 39392 3792 39420
rect 3786 39380 3792 39392
rect 3844 39380 3850 39432
rect 5810 39380 5816 39432
rect 5868 39420 5874 39432
rect 6365 39423 6423 39429
rect 6365 39420 6377 39423
rect 5868 39392 6377 39420
rect 5868 39380 5874 39392
rect 6365 39389 6377 39392
rect 6411 39389 6423 39423
rect 6365 39383 6423 39389
rect 6632 39423 6690 39429
rect 6632 39389 6644 39423
rect 6678 39420 6690 39423
rect 7742 39420 7748 39432
rect 6678 39392 7748 39420
rect 6678 39389 6690 39392
rect 6632 39383 6690 39389
rect 3804 39352 3832 39380
rect 4062 39361 4068 39364
rect 1872 39324 3832 39352
rect 4056 39315 4068 39361
rect 4120 39352 4126 39364
rect 6380 39352 6408 39383
rect 7742 39380 7748 39392
rect 7800 39380 7806 39432
rect 6822 39352 6828 39364
rect 4120 39324 4156 39352
rect 6380 39324 6828 39352
rect 4062 39312 4068 39315
rect 4120 39312 4126 39324
rect 6822 39312 6828 39324
rect 6880 39312 6886 39364
rect 8478 39312 8484 39364
rect 8536 39352 8542 39364
rect 9186 39355 9244 39361
rect 9186 39352 9198 39355
rect 8536 39324 9198 39352
rect 8536 39312 8542 39324
rect 9186 39321 9198 39324
rect 9232 39321 9244 39355
rect 11532 39352 11560 39587
rect 11716 39429 11744 39596
rect 17880 39556 17908 39596
rect 18046 39584 18052 39596
rect 18104 39584 18110 39636
rect 20806 39624 20812 39636
rect 18156 39596 20812 39624
rect 18156 39556 18184 39596
rect 20806 39584 20812 39596
rect 20864 39584 20870 39636
rect 27157 39627 27215 39633
rect 27157 39593 27169 39627
rect 27203 39624 27215 39627
rect 29638 39624 29644 39636
rect 27203 39596 29644 39624
rect 27203 39593 27215 39596
rect 27157 39587 27215 39593
rect 29638 39584 29644 39596
rect 29696 39584 29702 39636
rect 32309 39627 32367 39633
rect 32309 39593 32321 39627
rect 32355 39624 32367 39627
rect 32398 39624 32404 39636
rect 32355 39596 32404 39624
rect 32355 39593 32367 39596
rect 32309 39587 32367 39593
rect 32398 39584 32404 39596
rect 32456 39584 32462 39636
rect 34054 39584 34060 39636
rect 34112 39624 34118 39636
rect 34149 39627 34207 39633
rect 34149 39624 34161 39627
rect 34112 39596 34161 39624
rect 34112 39584 34118 39596
rect 34149 39593 34161 39596
rect 34195 39593 34207 39627
rect 34149 39587 34207 39593
rect 37366 39584 37372 39636
rect 37424 39624 37430 39636
rect 37461 39627 37519 39633
rect 37461 39624 37473 39627
rect 37424 39596 37473 39624
rect 37424 39584 37430 39596
rect 37461 39593 37473 39596
rect 37507 39593 37519 39627
rect 37461 39587 37519 39593
rect 39114 39584 39120 39636
rect 39172 39624 39178 39636
rect 39301 39627 39359 39633
rect 39301 39624 39313 39627
rect 39172 39596 39313 39624
rect 39172 39584 39178 39596
rect 39301 39593 39313 39596
rect 39347 39593 39359 39627
rect 39301 39587 39359 39593
rect 40313 39627 40371 39633
rect 40313 39593 40325 39627
rect 40359 39624 40371 39627
rect 40402 39624 40408 39636
rect 40359 39596 40408 39624
rect 40359 39593 40371 39596
rect 40313 39587 40371 39593
rect 40402 39584 40408 39596
rect 40460 39584 40466 39636
rect 43806 39624 43812 39636
rect 43767 39596 43812 39624
rect 43806 39584 43812 39596
rect 43864 39584 43870 39636
rect 47762 39624 47768 39636
rect 47723 39596 47768 39624
rect 47762 39584 47768 39596
rect 47820 39584 47826 39636
rect 17880 39528 18184 39556
rect 12158 39488 12164 39500
rect 12119 39460 12164 39488
rect 12158 39448 12164 39460
rect 12216 39448 12222 39500
rect 32766 39488 32772 39500
rect 32727 39460 32772 39488
rect 32766 39448 32772 39460
rect 32824 39448 32830 39500
rect 34330 39448 34336 39500
rect 34388 39488 34394 39500
rect 36081 39491 36139 39497
rect 36081 39488 36093 39491
rect 34388 39460 36093 39488
rect 34388 39448 34394 39460
rect 36081 39457 36093 39460
rect 36127 39457 36139 39491
rect 36081 39451 36139 39457
rect 37826 39448 37832 39500
rect 37884 39488 37890 39500
rect 37921 39491 37979 39497
rect 37921 39488 37933 39491
rect 37884 39460 37933 39488
rect 37884 39448 37890 39460
rect 37921 39457 37933 39460
rect 37967 39457 37979 39491
rect 42426 39488 42432 39500
rect 42387 39460 42432 39488
rect 37921 39451 37979 39457
rect 42426 39448 42432 39460
rect 42484 39448 42490 39500
rect 47946 39448 47952 39500
rect 48004 39488 48010 39500
rect 48222 39488 48228 39500
rect 48004 39460 48228 39488
rect 48004 39448 48010 39460
rect 48222 39448 48228 39460
rect 48280 39448 48286 39500
rect 11701 39423 11759 39429
rect 11701 39389 11713 39423
rect 11747 39389 11759 39423
rect 11701 39383 11759 39389
rect 12428 39423 12486 39429
rect 12428 39389 12440 39423
rect 12474 39420 12486 39423
rect 13538 39420 13544 39432
rect 12474 39392 13544 39420
rect 12474 39389 12486 39392
rect 12428 39383 12486 39389
rect 13538 39380 13544 39392
rect 13596 39380 13602 39432
rect 14185 39423 14243 39429
rect 14185 39389 14197 39423
rect 14231 39389 14243 39423
rect 14185 39383 14243 39389
rect 14452 39423 14510 39429
rect 14452 39389 14464 39423
rect 14498 39420 14510 39423
rect 16114 39420 16120 39432
rect 14498 39392 16120 39420
rect 14498 39389 14510 39392
rect 14452 39383 14510 39389
rect 13354 39352 13360 39364
rect 11532 39324 13360 39352
rect 9186 39315 9244 39321
rect 13354 39312 13360 39324
rect 13412 39312 13418 39364
rect 14200 39352 14228 39383
rect 16114 39380 16120 39392
rect 16172 39380 16178 39432
rect 16669 39423 16727 39429
rect 16669 39389 16681 39423
rect 16715 39420 16727 39423
rect 17310 39420 17316 39432
rect 16715 39392 17316 39420
rect 16715 39389 16727 39392
rect 16669 39383 16727 39389
rect 17310 39380 17316 39392
rect 17368 39420 17374 39432
rect 18506 39420 18512 39432
rect 17368 39392 18512 39420
rect 17368 39380 17374 39392
rect 18506 39380 18512 39392
rect 18564 39420 18570 39432
rect 19245 39423 19303 39429
rect 19245 39420 19257 39423
rect 18564 39392 19257 39420
rect 18564 39380 18570 39392
rect 19245 39389 19257 39392
rect 19291 39389 19303 39423
rect 19245 39383 19303 39389
rect 19334 39380 19340 39432
rect 19392 39420 19398 39432
rect 19501 39423 19559 39429
rect 19501 39420 19513 39423
rect 19392 39392 19513 39420
rect 19392 39380 19398 39392
rect 19501 39389 19513 39392
rect 19547 39389 19559 39423
rect 19501 39383 19559 39389
rect 22465 39423 22523 39429
rect 22465 39389 22477 39423
rect 22511 39420 22523 39423
rect 22554 39420 22560 39432
rect 22511 39392 22560 39420
rect 22511 39389 22523 39392
rect 22465 39383 22523 39389
rect 22554 39380 22560 39392
rect 22612 39380 22618 39432
rect 22732 39423 22790 39429
rect 22732 39389 22744 39423
rect 22778 39420 22790 39423
rect 24302 39420 24308 39432
rect 22778 39392 24308 39420
rect 22778 39389 22790 39392
rect 22732 39383 22790 39389
rect 24302 39380 24308 39392
rect 24360 39380 24366 39432
rect 24394 39380 24400 39432
rect 24452 39420 24458 39432
rect 25777 39423 25835 39429
rect 25777 39420 25789 39423
rect 24452 39392 25789 39420
rect 24452 39380 24458 39392
rect 25777 39389 25789 39392
rect 25823 39420 25835 39423
rect 27617 39423 27675 39429
rect 27617 39420 27629 39423
rect 25823 39392 27629 39420
rect 25823 39389 25835 39392
rect 25777 39383 25835 39389
rect 27617 39389 27629 39392
rect 27663 39389 27675 39423
rect 27617 39383 27675 39389
rect 30190 39380 30196 39432
rect 30248 39420 30254 39432
rect 30929 39423 30987 39429
rect 30929 39420 30941 39423
rect 30248 39392 30941 39420
rect 30248 39380 30254 39392
rect 30929 39389 30941 39392
rect 30975 39389 30987 39423
rect 30929 39383 30987 39389
rect 31196 39423 31254 39429
rect 31196 39389 31208 39423
rect 31242 39420 31254 39423
rect 31754 39420 31760 39432
rect 31242 39392 31760 39420
rect 31242 39389 31254 39392
rect 31196 39383 31254 39389
rect 14734 39352 14740 39364
rect 14200 39324 14740 39352
rect 14734 39312 14740 39324
rect 14792 39312 14798 39364
rect 16936 39355 16994 39361
rect 16936 39321 16948 39355
rect 16982 39352 16994 39355
rect 18322 39352 18328 39364
rect 16982 39324 18328 39352
rect 16982 39321 16994 39324
rect 16936 39315 16994 39321
rect 18322 39312 18328 39324
rect 18380 39312 18386 39364
rect 26044 39355 26102 39361
rect 26044 39321 26056 39355
rect 26090 39352 26102 39355
rect 27522 39352 27528 39364
rect 26090 39324 27528 39352
rect 26090 39321 26102 39324
rect 26044 39315 26102 39321
rect 27522 39312 27528 39324
rect 27580 39312 27586 39364
rect 27884 39355 27942 39361
rect 27884 39321 27896 39355
rect 27930 39352 27942 39355
rect 30282 39352 30288 39364
rect 27930 39324 30288 39352
rect 27930 39321 27942 39324
rect 27884 39315 27942 39321
rect 30282 39312 30288 39324
rect 30340 39312 30346 39364
rect 30944 39352 30972 39383
rect 31754 39380 31760 39392
rect 31812 39380 31818 39432
rect 33036 39423 33094 39429
rect 33036 39389 33048 39423
rect 33082 39420 33094 39423
rect 34146 39420 34152 39432
rect 33082 39392 34152 39420
rect 33082 39389 33094 39392
rect 33036 39383 33094 39389
rect 34146 39380 34152 39392
rect 34204 39380 34210 39432
rect 36348 39423 36406 39429
rect 36348 39389 36360 39423
rect 36394 39420 36406 39423
rect 37458 39420 37464 39432
rect 36394 39392 37464 39420
rect 36394 39389 36406 39392
rect 36348 39383 36406 39389
rect 37458 39380 37464 39392
rect 37516 39380 37522 39432
rect 38188 39423 38246 39429
rect 38188 39389 38200 39423
rect 38234 39420 38246 39423
rect 38930 39420 38936 39432
rect 38234 39392 38936 39420
rect 38234 39389 38246 39392
rect 38188 39383 38246 39389
rect 38930 39380 38936 39392
rect 38988 39380 38994 39432
rect 40310 39380 40316 39432
rect 40368 39420 40374 39432
rect 40497 39423 40555 39429
rect 40497 39420 40509 39423
rect 40368 39392 40509 39420
rect 40368 39380 40374 39392
rect 40497 39389 40509 39392
rect 40543 39420 40555 39423
rect 40954 39420 40960 39432
rect 40543 39392 40960 39420
rect 40543 39389 40555 39392
rect 40497 39383 40555 39389
rect 40954 39380 40960 39392
rect 41012 39420 41018 39432
rect 46198 39420 46204 39432
rect 41012 39392 46204 39420
rect 41012 39380 41018 39392
rect 46198 39380 46204 39392
rect 46256 39380 46262 39432
rect 46385 39423 46443 39429
rect 46385 39389 46397 39423
rect 46431 39420 46443 39423
rect 47964 39420 47992 39448
rect 46431 39392 47992 39420
rect 48492 39423 48550 39429
rect 46431 39389 46443 39392
rect 46385 39383 46443 39389
rect 48492 39389 48504 39423
rect 48538 39420 48550 39423
rect 49602 39420 49608 39432
rect 48538 39392 49608 39420
rect 48538 39389 48550 39392
rect 48492 39383 48550 39389
rect 49602 39380 49608 39392
rect 49660 39380 49666 39432
rect 50893 39423 50951 39429
rect 50893 39389 50905 39423
rect 50939 39420 50951 39423
rect 52730 39420 52736 39432
rect 50939 39392 52736 39420
rect 50939 39389 50951 39392
rect 50893 39383 50951 39389
rect 52730 39380 52736 39392
rect 52788 39420 52794 39432
rect 53466 39420 53472 39432
rect 52788 39392 53472 39420
rect 52788 39380 52794 39392
rect 53466 39380 53472 39392
rect 53524 39380 53530 39432
rect 32766 39352 32772 39364
rect 30944 39324 32772 39352
rect 32766 39312 32772 39324
rect 32824 39312 32830 39364
rect 42696 39355 42754 39361
rect 42696 39321 42708 39355
rect 42742 39352 42754 39355
rect 43714 39352 43720 39364
rect 42742 39324 43720 39352
rect 42742 39321 42754 39324
rect 42696 39315 42754 39321
rect 43714 39312 43720 39324
rect 43772 39312 43778 39364
rect 46652 39355 46710 39361
rect 46652 39321 46664 39355
rect 46698 39352 46710 39355
rect 49050 39352 49056 39364
rect 46698 39324 49056 39352
rect 46698 39321 46710 39324
rect 46652 39315 46710 39321
rect 49050 39312 49056 39324
rect 49108 39312 49114 39364
rect 51160 39355 51218 39361
rect 51160 39321 51172 39355
rect 51206 39352 51218 39355
rect 52822 39352 52828 39364
rect 51206 39324 52828 39352
rect 51206 39321 51218 39324
rect 51160 39315 51218 39321
rect 52822 39312 52828 39324
rect 52880 39312 52886 39364
rect 53006 39361 53012 39364
rect 53000 39315 53012 39361
rect 53064 39352 53070 39364
rect 53064 39324 53100 39352
rect 53006 39312 53012 39315
rect 53064 39312 53070 39324
rect 10318 39284 10324 39296
rect 10279 39256 10324 39284
rect 10318 39244 10324 39256
rect 10376 39244 10382 39296
rect 13538 39284 13544 39296
rect 13499 39256 13544 39284
rect 13538 39244 13544 39256
rect 13596 39244 13602 39296
rect 14826 39244 14832 39296
rect 14884 39284 14890 39296
rect 15565 39287 15623 39293
rect 15565 39284 15577 39287
rect 14884 39256 15577 39284
rect 14884 39244 14890 39256
rect 15565 39253 15577 39256
rect 15611 39253 15623 39287
rect 20622 39284 20628 39296
rect 20583 39256 20628 39284
rect 15565 39247 15623 39253
rect 20622 39244 20628 39256
rect 20680 39244 20686 39296
rect 23842 39284 23848 39296
rect 23803 39256 23848 39284
rect 23842 39244 23848 39256
rect 23900 39244 23906 39296
rect 27614 39244 27620 39296
rect 27672 39284 27678 39296
rect 28997 39287 29055 39293
rect 28997 39284 29009 39287
rect 27672 39256 29009 39284
rect 27672 39244 27678 39256
rect 28997 39253 29009 39256
rect 29043 39253 29055 39287
rect 49602 39284 49608 39296
rect 49563 39256 49608 39284
rect 28997 39247 29055 39253
rect 49602 39244 49608 39256
rect 49660 39244 49666 39296
rect 52270 39284 52276 39296
rect 52231 39256 52276 39284
rect 52270 39244 52276 39256
rect 52328 39244 52334 39296
rect 53926 39244 53932 39296
rect 53984 39284 53990 39296
rect 54113 39287 54171 39293
rect 54113 39284 54125 39287
rect 53984 39256 54125 39284
rect 53984 39244 53990 39256
rect 54113 39253 54125 39256
rect 54159 39253 54171 39287
rect 54113 39247 54171 39253
rect 1104 39194 59340 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 59340 39194
rect 1104 39120 59340 39142
rect 8478 39080 8484 39092
rect 8439 39052 8484 39080
rect 8478 39040 8484 39052
rect 8536 39040 8542 39092
rect 18322 39080 18328 39092
rect 18283 39052 18328 39080
rect 18322 39040 18328 39052
rect 18380 39040 18386 39092
rect 23014 39040 23020 39092
rect 23072 39080 23078 39092
rect 24213 39083 24271 39089
rect 24213 39080 24225 39083
rect 23072 39052 24225 39080
rect 23072 39040 23078 39052
rect 24213 39049 24225 39052
rect 24259 39049 24271 39083
rect 24213 39043 24271 39049
rect 28353 39083 28411 39089
rect 28353 39049 28365 39083
rect 28399 39080 28411 39083
rect 28442 39080 28448 39092
rect 28399 39052 28448 39080
rect 28399 39049 28411 39052
rect 28353 39043 28411 39049
rect 28442 39040 28448 39052
rect 28500 39040 28506 39092
rect 31570 39080 31576 39092
rect 31531 39052 31576 39080
rect 31570 39040 31576 39052
rect 31628 39040 31634 39092
rect 34238 39080 34244 39092
rect 34199 39052 34244 39080
rect 34238 39040 34244 39052
rect 34296 39040 34302 39092
rect 40218 39080 40224 39092
rect 40179 39052 40224 39080
rect 40218 39040 40224 39052
rect 40276 39040 40282 39092
rect 43714 39040 43720 39092
rect 43772 39080 43778 39092
rect 43809 39083 43867 39089
rect 43809 39080 43821 39083
rect 43772 39052 43821 39080
rect 43772 39040 43778 39052
rect 43809 39049 43821 39052
rect 43855 39049 43867 39083
rect 49326 39080 49332 39092
rect 49287 39052 49332 39080
rect 43809 39043 43867 39049
rect 49326 39040 49332 39052
rect 49384 39040 49390 39092
rect 56689 39083 56747 39089
rect 56689 39080 56701 39083
rect 55186 39052 56701 39080
rect 7368 39015 7426 39021
rect 7368 38981 7380 39015
rect 7414 39012 7426 39015
rect 8386 39012 8392 39024
rect 7414 38984 8392 39012
rect 7414 38981 7426 38984
rect 7368 38975 7426 38981
rect 8386 38972 8392 38984
rect 8444 38972 8450 39024
rect 9208 39015 9266 39021
rect 9208 38981 9220 39015
rect 9254 39012 9266 39015
rect 10318 39012 10324 39024
rect 9254 38984 10324 39012
rect 9254 38981 9266 38984
rect 9208 38975 9266 38981
rect 10318 38972 10324 38984
rect 10376 38972 10382 39024
rect 12428 39015 12486 39021
rect 12428 38981 12440 39015
rect 12474 39012 12486 39015
rect 13538 39012 13544 39024
rect 12474 38984 13544 39012
rect 12474 38981 12486 38984
rect 12428 38975 12486 38981
rect 13538 38972 13544 38984
rect 13596 38972 13602 39024
rect 19052 39015 19110 39021
rect 19052 38981 19064 39015
rect 19098 39012 19110 39015
rect 20622 39012 20628 39024
rect 19098 38984 20628 39012
rect 19098 38981 19110 38984
rect 19052 38975 19110 38981
rect 20622 38972 20628 38984
rect 20680 38972 20686 39024
rect 23100 39015 23158 39021
rect 23100 38981 23112 39015
rect 23146 39012 23158 39015
rect 23842 39012 23848 39024
rect 23146 38984 23848 39012
rect 23146 38981 23158 38984
rect 23100 38975 23158 38981
rect 23842 38972 23848 38984
rect 23900 38972 23906 39024
rect 27706 39012 27712 39024
rect 26988 38984 27712 39012
rect 4056 38947 4114 38953
rect 4056 38913 4068 38947
rect 4102 38944 4114 38947
rect 5718 38944 5724 38956
rect 4102 38916 5724 38944
rect 4102 38913 4114 38916
rect 4056 38907 4114 38913
rect 5718 38904 5724 38916
rect 5776 38904 5782 38956
rect 6822 38904 6828 38956
rect 6880 38944 6886 38956
rect 7101 38947 7159 38953
rect 7101 38944 7113 38947
rect 6880 38916 7113 38944
rect 6880 38904 6886 38916
rect 7101 38913 7113 38916
rect 7147 38913 7159 38947
rect 8938 38944 8944 38956
rect 8899 38916 8944 38944
rect 7101 38907 7159 38913
rect 8938 38904 8944 38916
rect 8996 38904 9002 38956
rect 12158 38944 12164 38956
rect 12119 38916 12164 38944
rect 12158 38904 12164 38916
rect 12216 38904 12222 38956
rect 17212 38947 17270 38953
rect 17212 38913 17224 38947
rect 17258 38944 17270 38947
rect 18046 38944 18052 38956
rect 17258 38916 18052 38944
rect 17258 38913 17270 38916
rect 17212 38907 17270 38913
rect 18046 38904 18052 38916
rect 18104 38904 18110 38956
rect 20806 38944 20812 38956
rect 20719 38916 20812 38944
rect 20806 38904 20812 38916
rect 20864 38904 20870 38956
rect 22833 38947 22891 38953
rect 22833 38913 22845 38947
rect 22879 38944 22891 38947
rect 24394 38944 24400 38956
rect 22879 38916 24400 38944
rect 22879 38913 22891 38916
rect 22833 38907 22891 38913
rect 24394 38904 24400 38916
rect 24452 38904 24458 38956
rect 26988 38953 27016 38984
rect 27706 38972 27712 38984
rect 27764 38972 27770 39024
rect 30460 39015 30518 39021
rect 30460 38981 30472 39015
rect 30506 39012 30518 39015
rect 31938 39012 31944 39024
rect 30506 38984 31944 39012
rect 30506 38981 30518 38984
rect 30460 38975 30518 38981
rect 31938 38972 31944 38984
rect 31996 38972 32002 39024
rect 33128 39015 33186 39021
rect 33128 38981 33140 39015
rect 33174 39012 33186 39015
rect 36262 39012 36268 39024
rect 33174 38984 36268 39012
rect 33174 38981 33186 38984
rect 33128 38975 33186 38981
rect 36262 38972 36268 38984
rect 36320 38972 36326 39024
rect 39108 39015 39166 39021
rect 39108 38981 39120 39015
rect 39154 39012 39166 39015
rect 39298 39012 39304 39024
rect 39154 38984 39304 39012
rect 39154 38981 39166 38984
rect 39108 38975 39166 38981
rect 39298 38972 39304 38984
rect 39356 38972 39362 39024
rect 45640 39015 45698 39021
rect 45640 38981 45652 39015
rect 45686 39012 45698 39015
rect 47026 39012 47032 39024
rect 45686 38984 47032 39012
rect 45686 38981 45698 38984
rect 45640 38975 45698 38981
rect 47026 38972 47032 38984
rect 47084 38972 47090 39024
rect 48216 39015 48274 39021
rect 48216 38981 48228 39015
rect 48262 39012 48274 39015
rect 49602 39012 49608 39024
rect 48262 38984 49608 39012
rect 48262 38981 48274 38984
rect 48216 38975 48274 38981
rect 49602 38972 49608 38984
rect 49660 38972 49666 39024
rect 51534 39012 51540 39024
rect 50540 38984 51540 39012
rect 26973 38947 27031 38953
rect 26973 38913 26985 38947
rect 27019 38913 27031 38947
rect 26973 38907 27031 38913
rect 27240 38947 27298 38953
rect 27240 38913 27252 38947
rect 27286 38944 27298 38947
rect 28534 38944 28540 38956
rect 27286 38916 28540 38944
rect 27286 38913 27298 38916
rect 27240 38907 27298 38913
rect 28534 38904 28540 38916
rect 28592 38904 28598 38956
rect 30190 38944 30196 38956
rect 30151 38916 30196 38944
rect 30190 38904 30196 38916
rect 30248 38904 30254 38956
rect 32766 38904 32772 38956
rect 32824 38944 32830 38956
rect 32861 38947 32919 38953
rect 32861 38944 32873 38947
rect 32824 38916 32873 38944
rect 32824 38904 32830 38916
rect 32861 38913 32873 38916
rect 32907 38913 32919 38947
rect 32861 38907 32919 38913
rect 34968 38947 35026 38953
rect 34968 38913 34980 38947
rect 35014 38944 35026 38947
rect 36078 38944 36084 38956
rect 35014 38916 36084 38944
rect 35014 38913 35026 38916
rect 34968 38907 35026 38913
rect 36078 38904 36084 38916
rect 36136 38904 36142 38956
rect 38746 38904 38752 38956
rect 38804 38944 38810 38956
rect 38841 38947 38899 38953
rect 38841 38944 38853 38947
rect 38804 38916 38853 38944
rect 38804 38904 38810 38916
rect 38841 38913 38853 38916
rect 38887 38913 38899 38947
rect 38841 38907 38899 38913
rect 42696 38947 42754 38953
rect 42696 38913 42708 38947
rect 42742 38944 42754 38947
rect 43990 38944 43996 38956
rect 42742 38916 43996 38944
rect 42742 38913 42754 38916
rect 42696 38907 42754 38913
rect 43990 38904 43996 38916
rect 44048 38904 44054 38956
rect 45186 38904 45192 38956
rect 45244 38944 45250 38956
rect 45373 38947 45431 38953
rect 45373 38944 45385 38947
rect 45244 38916 45385 38944
rect 45244 38904 45250 38916
rect 45373 38913 45385 38916
rect 45419 38913 45431 38947
rect 45373 38907 45431 38913
rect 46198 38904 46204 38956
rect 46256 38944 46262 38956
rect 50540 38953 50568 38984
rect 51534 38972 51540 38984
rect 51592 38972 51598 39024
rect 53736 39015 53794 39021
rect 53736 38981 53748 39015
rect 53782 39012 53794 39015
rect 55186 39012 55214 39052
rect 56689 39049 56701 39052
rect 56735 39049 56747 39083
rect 56689 39043 56747 39049
rect 53782 38984 55214 39012
rect 53782 38981 53794 38984
rect 53736 38975 53794 38981
rect 49973 38947 50031 38953
rect 49973 38944 49985 38947
rect 46256 38916 49985 38944
rect 46256 38904 46262 38916
rect 49973 38913 49985 38916
rect 50019 38913 50031 38947
rect 49973 38907 50031 38913
rect 50525 38947 50583 38953
rect 50525 38913 50537 38947
rect 50571 38913 50583 38947
rect 50525 38907 50583 38913
rect 50792 38947 50850 38953
rect 50792 38913 50804 38947
rect 50838 38944 50850 38947
rect 52086 38944 52092 38956
rect 50838 38916 52092 38944
rect 50838 38913 50850 38916
rect 50792 38907 50850 38913
rect 52086 38904 52092 38916
rect 52144 38904 52150 38956
rect 53466 38944 53472 38956
rect 53427 38916 53472 38944
rect 53466 38904 53472 38916
rect 53524 38904 53530 38956
rect 55576 38947 55634 38953
rect 55576 38913 55588 38947
rect 55622 38944 55634 38947
rect 56686 38944 56692 38956
rect 55622 38916 56692 38944
rect 55622 38913 55634 38916
rect 55576 38907 55634 38913
rect 56686 38904 56692 38916
rect 56744 38904 56750 38956
rect 3786 38876 3792 38888
rect 3699 38848 3792 38876
rect 3786 38836 3792 38848
rect 3844 38836 3850 38888
rect 16666 38836 16672 38888
rect 16724 38876 16730 38888
rect 16945 38879 17003 38885
rect 16945 38876 16957 38879
rect 16724 38848 16957 38876
rect 16724 38836 16730 38848
rect 16945 38845 16957 38848
rect 16991 38845 17003 38879
rect 16945 38839 17003 38845
rect 18506 38836 18512 38888
rect 18564 38876 18570 38888
rect 18785 38879 18843 38885
rect 18785 38876 18797 38879
rect 18564 38848 18797 38876
rect 18564 38836 18570 38848
rect 18785 38845 18797 38848
rect 18831 38845 18843 38879
rect 18785 38839 18843 38845
rect 3804 38740 3832 38836
rect 4982 38740 4988 38752
rect 3804 38712 4988 38740
rect 4982 38700 4988 38712
rect 5040 38700 5046 38752
rect 5166 38740 5172 38752
rect 5127 38712 5172 38740
rect 5166 38700 5172 38712
rect 5224 38700 5230 38752
rect 10318 38740 10324 38752
rect 10279 38712 10324 38740
rect 10318 38700 10324 38712
rect 10376 38700 10382 38752
rect 13538 38740 13544 38752
rect 13499 38712 13544 38740
rect 13538 38700 13544 38712
rect 13596 38700 13602 38752
rect 19518 38700 19524 38752
rect 19576 38740 19582 38752
rect 20165 38743 20223 38749
rect 20165 38740 20177 38743
rect 19576 38712 20177 38740
rect 19576 38700 19582 38712
rect 20165 38709 20177 38712
rect 20211 38709 20223 38743
rect 20165 38703 20223 38709
rect 20530 38700 20536 38752
rect 20588 38740 20594 38752
rect 20625 38743 20683 38749
rect 20625 38740 20637 38743
rect 20588 38712 20637 38740
rect 20588 38700 20594 38712
rect 20625 38709 20637 38712
rect 20671 38709 20683 38743
rect 20824 38740 20852 38904
rect 34698 38876 34704 38888
rect 34659 38848 34704 38876
rect 34698 38836 34704 38848
rect 34756 38836 34762 38888
rect 42426 38876 42432 38888
rect 42387 38848 42432 38876
rect 42426 38836 42432 38848
rect 42484 38836 42490 38888
rect 47486 38836 47492 38888
rect 47544 38876 47550 38888
rect 47946 38876 47952 38888
rect 47544 38848 47952 38876
rect 47544 38836 47550 38848
rect 47946 38836 47952 38848
rect 48004 38836 48010 38888
rect 55306 38876 55312 38888
rect 55186 38848 55312 38876
rect 55186 38808 55214 38848
rect 55306 38836 55312 38848
rect 55364 38836 55370 38888
rect 54404 38780 55214 38808
rect 30834 38740 30840 38752
rect 20824 38712 30840 38740
rect 20625 38703 20683 38709
rect 30834 38700 30840 38712
rect 30892 38700 30898 38752
rect 36081 38743 36139 38749
rect 36081 38709 36093 38743
rect 36127 38740 36139 38743
rect 36630 38740 36636 38752
rect 36127 38712 36636 38740
rect 36127 38709 36139 38712
rect 36081 38703 36139 38709
rect 36630 38700 36636 38712
rect 36688 38700 36694 38752
rect 46750 38740 46756 38752
rect 46711 38712 46756 38740
rect 46750 38700 46756 38712
rect 46808 38700 46814 38752
rect 49786 38740 49792 38752
rect 49747 38712 49792 38740
rect 49786 38700 49792 38712
rect 49844 38700 49850 38752
rect 49878 38700 49884 38752
rect 49936 38740 49942 38752
rect 51905 38743 51963 38749
rect 51905 38740 51917 38743
rect 49936 38712 51917 38740
rect 49936 38700 49942 38712
rect 51905 38709 51917 38712
rect 51951 38709 51963 38743
rect 51905 38703 51963 38709
rect 53742 38700 53748 38752
rect 53800 38740 53806 38752
rect 54404 38740 54432 38780
rect 54846 38740 54852 38752
rect 53800 38712 54432 38740
rect 54807 38712 54852 38740
rect 53800 38700 53806 38712
rect 54846 38700 54852 38712
rect 54904 38700 54910 38752
rect 1104 38650 59340 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 59340 38650
rect 1104 38576 59340 38598
rect 27522 38496 27528 38548
rect 27580 38536 27586 38548
rect 27617 38539 27675 38545
rect 27617 38536 27629 38539
rect 27580 38508 27629 38536
rect 27580 38496 27586 38508
rect 27617 38505 27629 38508
rect 27663 38505 27675 38539
rect 31110 38536 31116 38548
rect 31071 38508 31116 38536
rect 27617 38499 27675 38505
rect 31110 38496 31116 38508
rect 31168 38496 31174 38548
rect 36078 38536 36084 38548
rect 36039 38508 36084 38536
rect 36078 38496 36084 38508
rect 36136 38496 36142 38548
rect 46842 38536 46848 38548
rect 46803 38508 46848 38536
rect 46842 38496 46848 38508
rect 46900 38496 46906 38548
rect 52917 38539 52975 38545
rect 52917 38505 52929 38539
rect 52963 38536 52975 38539
rect 53006 38536 53012 38548
rect 52963 38508 53012 38536
rect 52963 38505 52975 38508
rect 52917 38499 52975 38505
rect 53006 38496 53012 38508
rect 53064 38496 53070 38548
rect 53742 38536 53748 38548
rect 53392 38508 53748 38536
rect 47486 38400 47492 38412
rect 47447 38372 47492 38400
rect 47486 38360 47492 38372
rect 47544 38360 47550 38412
rect 53392 38409 53420 38508
rect 53742 38496 53748 38508
rect 53800 38496 53806 38548
rect 56686 38536 56692 38548
rect 56647 38508 56692 38536
rect 56686 38496 56692 38508
rect 56744 38496 56750 38548
rect 53377 38403 53435 38409
rect 53377 38369 53389 38403
rect 53423 38369 53435 38403
rect 53377 38363 53435 38369
rect 4982 38332 4988 38344
rect 4943 38304 4988 38332
rect 4982 38292 4988 38304
rect 5040 38292 5046 38344
rect 8938 38332 8944 38344
rect 8899 38304 8944 38332
rect 8938 38292 8944 38304
rect 8996 38292 9002 38344
rect 9208 38335 9266 38341
rect 9208 38301 9220 38335
rect 9254 38332 9266 38335
rect 10318 38332 10324 38344
rect 9254 38304 10324 38332
rect 9254 38301 9266 38304
rect 9208 38295 9266 38301
rect 10318 38292 10324 38304
rect 10376 38292 10382 38344
rect 12069 38335 12127 38341
rect 12069 38301 12081 38335
rect 12115 38332 12127 38335
rect 12158 38332 12164 38344
rect 12115 38304 12164 38332
rect 12115 38301 12127 38304
rect 12069 38295 12127 38301
rect 12158 38292 12164 38304
rect 12216 38292 12222 38344
rect 12336 38335 12394 38341
rect 12336 38301 12348 38335
rect 12382 38332 12394 38335
rect 13538 38332 13544 38344
rect 12382 38304 13544 38332
rect 12382 38301 12394 38304
rect 12336 38295 12394 38301
rect 13538 38292 13544 38304
rect 13596 38292 13602 38344
rect 14645 38335 14703 38341
rect 14645 38301 14657 38335
rect 14691 38332 14703 38335
rect 14734 38332 14740 38344
rect 14691 38304 14740 38332
rect 14691 38301 14703 38304
rect 14645 38295 14703 38301
rect 14734 38292 14740 38304
rect 14792 38332 14798 38344
rect 19518 38341 19524 38344
rect 16485 38335 16543 38341
rect 16485 38332 16497 38335
rect 14792 38304 16497 38332
rect 14792 38292 14798 38304
rect 16485 38301 16497 38304
rect 16531 38301 16543 38335
rect 16485 38295 16543 38301
rect 19245 38335 19303 38341
rect 19245 38301 19257 38335
rect 19291 38301 19303 38335
rect 19512 38332 19524 38341
rect 19479 38304 19524 38332
rect 19245 38295 19303 38301
rect 19512 38295 19524 38304
rect 5252 38267 5310 38273
rect 5252 38233 5264 38267
rect 5298 38264 5310 38267
rect 5810 38264 5816 38276
rect 5298 38236 5816 38264
rect 5298 38233 5310 38236
rect 5252 38227 5310 38233
rect 5810 38224 5816 38236
rect 5868 38224 5874 38276
rect 14912 38267 14970 38273
rect 14912 38233 14924 38267
rect 14958 38264 14970 38267
rect 15838 38264 15844 38276
rect 14958 38236 15844 38264
rect 14958 38233 14970 38236
rect 14912 38227 14970 38233
rect 15838 38224 15844 38236
rect 15896 38224 15902 38276
rect 16752 38267 16810 38273
rect 16752 38233 16764 38267
rect 16798 38264 16810 38267
rect 17954 38264 17960 38276
rect 16798 38236 17960 38264
rect 16798 38233 16810 38236
rect 16752 38227 16810 38233
rect 17954 38224 17960 38236
rect 18012 38224 18018 38276
rect 18506 38224 18512 38276
rect 18564 38264 18570 38276
rect 19260 38264 19288 38295
rect 19518 38292 19524 38295
rect 19576 38292 19582 38344
rect 21082 38332 21088 38344
rect 20995 38304 21088 38332
rect 21082 38292 21088 38304
rect 21140 38332 21146 38344
rect 21818 38332 21824 38344
rect 21140 38304 21824 38332
rect 21140 38292 21146 38304
rect 21818 38292 21824 38304
rect 21876 38292 21882 38344
rect 24394 38332 24400 38344
rect 24355 38304 24400 38332
rect 24394 38292 24400 38304
rect 24452 38292 24458 38344
rect 26234 38292 26240 38344
rect 26292 38332 26298 38344
rect 30006 38341 30012 38344
rect 29733 38335 29791 38341
rect 26292 38304 26337 38332
rect 26292 38292 26298 38304
rect 29733 38301 29745 38335
rect 29779 38301 29791 38335
rect 30000 38332 30012 38341
rect 29967 38304 30012 38332
rect 29733 38295 29791 38301
rect 30000 38295 30012 38304
rect 21100 38264 21128 38292
rect 18564 38236 21128 38264
rect 21352 38267 21410 38273
rect 18564 38224 18570 38236
rect 21352 38233 21364 38267
rect 21398 38264 21410 38267
rect 22370 38264 22376 38276
rect 21398 38236 22376 38264
rect 21398 38233 21410 38236
rect 21352 38227 21410 38233
rect 22370 38224 22376 38236
rect 22428 38224 22434 38276
rect 24664 38267 24722 38273
rect 24664 38233 24676 38267
rect 24710 38264 24722 38267
rect 26504 38267 26562 38273
rect 24710 38236 26464 38264
rect 24710 38233 24722 38236
rect 24664 38227 24722 38233
rect 6362 38196 6368 38208
rect 6323 38168 6368 38196
rect 6362 38156 6368 38168
rect 6420 38156 6426 38208
rect 10318 38196 10324 38208
rect 10279 38168 10324 38196
rect 10318 38156 10324 38168
rect 10376 38156 10382 38208
rect 13446 38196 13452 38208
rect 13407 38168 13452 38196
rect 13446 38156 13452 38168
rect 13504 38156 13510 38208
rect 16025 38199 16083 38205
rect 16025 38165 16037 38199
rect 16071 38196 16083 38199
rect 16942 38196 16948 38208
rect 16071 38168 16948 38196
rect 16071 38165 16083 38168
rect 16025 38159 16083 38165
rect 16942 38156 16948 38168
rect 17000 38156 17006 38208
rect 17862 38196 17868 38208
rect 17823 38168 17868 38196
rect 17862 38156 17868 38168
rect 17920 38156 17926 38208
rect 20622 38196 20628 38208
rect 20583 38168 20628 38196
rect 20622 38156 20628 38168
rect 20680 38156 20686 38208
rect 22186 38156 22192 38208
rect 22244 38196 22250 38208
rect 22465 38199 22523 38205
rect 22465 38196 22477 38199
rect 22244 38168 22477 38196
rect 22244 38156 22250 38168
rect 22465 38165 22477 38168
rect 22511 38165 22523 38199
rect 22465 38159 22523 38165
rect 25777 38199 25835 38205
rect 25777 38165 25789 38199
rect 25823 38196 25835 38199
rect 26326 38196 26332 38208
rect 25823 38168 26332 38196
rect 25823 38165 25835 38168
rect 25777 38159 25835 38165
rect 26326 38156 26332 38168
rect 26384 38156 26390 38208
rect 26436 38196 26464 38236
rect 26504 38233 26516 38267
rect 26550 38264 26562 38267
rect 27706 38264 27712 38276
rect 26550 38236 27712 38264
rect 26550 38233 26562 38236
rect 26504 38227 26562 38233
rect 27706 38224 27712 38236
rect 27764 38224 27770 38276
rect 29748 38264 29776 38295
rect 30006 38292 30012 38295
rect 30064 38292 30070 38344
rect 31754 38292 31760 38344
rect 31812 38332 31818 38344
rect 32493 38335 32551 38341
rect 32493 38332 32505 38335
rect 31812 38304 32505 38332
rect 31812 38292 31818 38304
rect 32493 38301 32505 38304
rect 32539 38301 32551 38335
rect 34698 38332 34704 38344
rect 34659 38304 34704 38332
rect 32493 38295 32551 38301
rect 34698 38292 34704 38304
rect 34756 38292 34762 38344
rect 36541 38335 36599 38341
rect 36541 38301 36553 38335
rect 36587 38332 36599 38335
rect 38746 38332 38752 38344
rect 36587 38304 38752 38332
rect 36587 38301 36599 38304
rect 36541 38295 36599 38301
rect 38746 38292 38752 38304
rect 38804 38292 38810 38344
rect 42426 38292 42432 38344
rect 42484 38332 42490 38344
rect 42889 38335 42947 38341
rect 42889 38332 42901 38335
rect 42484 38304 42901 38332
rect 42484 38292 42490 38304
rect 42889 38301 42901 38304
rect 42935 38301 42947 38335
rect 42889 38295 42947 38301
rect 45186 38292 45192 38344
rect 45244 38332 45250 38344
rect 45465 38335 45523 38341
rect 45465 38332 45477 38335
rect 45244 38304 45477 38332
rect 45244 38292 45250 38304
rect 45465 38301 45477 38304
rect 45511 38301 45523 38335
rect 45465 38295 45523 38301
rect 45732 38335 45790 38341
rect 45732 38301 45744 38335
rect 45778 38332 45790 38335
rect 46750 38332 46756 38344
rect 45778 38304 46756 38332
rect 45778 38301 45790 38304
rect 45732 38295 45790 38301
rect 30190 38264 30196 38276
rect 29748 38236 30196 38264
rect 30190 38224 30196 38236
rect 30248 38224 30254 38276
rect 32760 38267 32818 38273
rect 32760 38233 32772 38267
rect 32806 38264 32818 38267
rect 33502 38264 33508 38276
rect 32806 38236 33508 38264
rect 32806 38233 32818 38236
rect 32760 38227 32818 38233
rect 33502 38224 33508 38236
rect 33560 38224 33566 38276
rect 34968 38267 35026 38273
rect 34968 38233 34980 38267
rect 35014 38264 35026 38267
rect 35342 38264 35348 38276
rect 35014 38236 35348 38264
rect 35014 38233 35026 38236
rect 34968 38227 35026 38233
rect 35342 38224 35348 38236
rect 35400 38224 35406 38276
rect 36808 38267 36866 38273
rect 36808 38233 36820 38267
rect 36854 38264 36866 38267
rect 37550 38264 37556 38276
rect 36854 38236 37556 38264
rect 36854 38233 36866 38236
rect 36808 38227 36866 38233
rect 37550 38224 37556 38236
rect 37608 38224 37614 38276
rect 43156 38267 43214 38273
rect 43156 38233 43168 38267
rect 43202 38264 43214 38267
rect 44450 38264 44456 38276
rect 43202 38236 44456 38264
rect 43202 38233 43214 38236
rect 43156 38227 43214 38233
rect 44450 38224 44456 38236
rect 44508 38224 44514 38276
rect 45480 38264 45508 38295
rect 46750 38292 46756 38304
rect 46808 38292 46814 38344
rect 51534 38332 51540 38344
rect 51447 38304 51540 38332
rect 51534 38292 51540 38304
rect 51592 38332 51598 38344
rect 53392 38332 53420 38363
rect 51592 38304 53420 38332
rect 53644 38335 53702 38341
rect 51592 38292 51598 38304
rect 53644 38301 53656 38335
rect 53690 38332 53702 38335
rect 54846 38332 54852 38344
rect 53690 38304 54852 38332
rect 53690 38301 53702 38304
rect 53644 38295 53702 38301
rect 54846 38292 54852 38304
rect 54904 38292 54910 38344
rect 55306 38332 55312 38344
rect 55267 38304 55312 38332
rect 55306 38292 55312 38304
rect 55364 38292 55370 38344
rect 47486 38264 47492 38276
rect 45480 38236 47492 38264
rect 47486 38224 47492 38236
rect 47544 38224 47550 38276
rect 47756 38267 47814 38273
rect 47756 38233 47768 38267
rect 47802 38264 47814 38267
rect 51442 38264 51448 38276
rect 47802 38236 51448 38264
rect 47802 38233 47814 38236
rect 47756 38227 47814 38233
rect 51442 38224 51448 38236
rect 51500 38224 51506 38276
rect 51804 38267 51862 38273
rect 51804 38233 51816 38267
rect 51850 38264 51862 38267
rect 53742 38264 53748 38276
rect 51850 38236 53748 38264
rect 51850 38233 51862 38236
rect 51804 38227 51862 38233
rect 53742 38224 53748 38236
rect 53800 38224 53806 38276
rect 55576 38267 55634 38273
rect 55576 38233 55588 38267
rect 55622 38264 55634 38267
rect 56686 38264 56692 38276
rect 55622 38236 56692 38264
rect 55622 38233 55634 38236
rect 55576 38227 55634 38233
rect 56686 38224 56692 38236
rect 56744 38224 56750 38276
rect 27798 38196 27804 38208
rect 26436 38168 27804 38196
rect 27798 38156 27804 38168
rect 27856 38156 27862 38208
rect 33873 38199 33931 38205
rect 33873 38165 33885 38199
rect 33919 38196 33931 38199
rect 34790 38196 34796 38208
rect 33919 38168 34796 38196
rect 33919 38165 33931 38168
rect 33873 38159 33931 38165
rect 34790 38156 34796 38168
rect 34848 38156 34854 38208
rect 37918 38196 37924 38208
rect 37879 38168 37924 38196
rect 37918 38156 37924 38168
rect 37976 38156 37982 38208
rect 44266 38196 44272 38208
rect 44227 38168 44272 38196
rect 44266 38156 44272 38168
rect 44324 38156 44330 38208
rect 47026 38156 47032 38208
rect 47084 38196 47090 38208
rect 48869 38199 48927 38205
rect 48869 38196 48881 38199
rect 47084 38168 48881 38196
rect 47084 38156 47090 38168
rect 48869 38165 48881 38168
rect 48915 38165 48927 38199
rect 48869 38159 48927 38165
rect 53834 38156 53840 38208
rect 53892 38196 53898 38208
rect 54757 38199 54815 38205
rect 54757 38196 54769 38199
rect 53892 38168 54769 38196
rect 53892 38156 53898 38168
rect 54757 38165 54769 38168
rect 54803 38165 54815 38199
rect 54757 38159 54815 38165
rect 1104 38106 59340 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 59340 38106
rect 1104 38032 59340 38054
rect 3973 37995 4031 38001
rect 3973 37961 3985 37995
rect 4019 37992 4031 37995
rect 4062 37992 4068 38004
rect 4019 37964 4068 37992
rect 4019 37961 4031 37964
rect 3973 37955 4031 37961
rect 4062 37952 4068 37964
rect 4120 37952 4126 38004
rect 5718 37952 5724 38004
rect 5776 37992 5782 38004
rect 5813 37995 5871 38001
rect 5813 37992 5825 37995
rect 5776 37964 5825 37992
rect 5776 37952 5782 37964
rect 5813 37961 5825 37964
rect 5859 37961 5871 37995
rect 15838 37992 15844 38004
rect 15799 37964 15844 37992
rect 5813 37955 5871 37961
rect 15838 37952 15844 37964
rect 15896 37952 15902 38004
rect 18046 37992 18052 38004
rect 18007 37964 18052 37992
rect 18046 37952 18052 37964
rect 18104 37952 18110 38004
rect 28534 37992 28540 38004
rect 28495 37964 28540 37992
rect 28534 37952 28540 37964
rect 28592 37952 28598 38004
rect 30282 37952 30288 38004
rect 30340 37992 30346 38004
rect 30469 37995 30527 38001
rect 30469 37992 30481 37995
rect 30340 37964 30481 37992
rect 30340 37952 30346 37964
rect 30469 37961 30481 37964
rect 30515 37961 30527 37995
rect 33502 37992 33508 38004
rect 33463 37964 33508 37992
rect 30469 37955 30527 37961
rect 33502 37952 33508 37964
rect 33560 37952 33566 38004
rect 35342 37992 35348 38004
rect 35303 37964 35348 37992
rect 35342 37952 35348 37964
rect 35400 37952 35406 38004
rect 44450 37992 44456 38004
rect 44411 37964 44456 37992
rect 44450 37952 44456 37964
rect 44508 37952 44514 38004
rect 4700 37927 4758 37933
rect 4700 37893 4712 37927
rect 4746 37924 4758 37927
rect 6362 37924 6368 37936
rect 4746 37896 6368 37924
rect 4746 37893 4758 37896
rect 4700 37887 4758 37893
rect 6362 37884 6368 37896
rect 6420 37884 6426 37936
rect 8656 37927 8714 37933
rect 8656 37893 8668 37927
rect 8702 37924 8714 37927
rect 10318 37924 10324 37936
rect 8702 37896 10324 37924
rect 8702 37893 8714 37896
rect 8656 37887 8714 37893
rect 10318 37884 10324 37896
rect 10376 37884 10382 37936
rect 12060 37927 12118 37933
rect 12060 37893 12072 37927
rect 12106 37924 12118 37927
rect 13446 37924 13452 37936
rect 12106 37896 13452 37924
rect 12106 37893 12118 37896
rect 12060 37887 12118 37893
rect 13446 37884 13452 37896
rect 13504 37884 13510 37936
rect 16936 37927 16994 37933
rect 14476 37896 16574 37924
rect 2860 37859 2918 37865
rect 2860 37825 2872 37859
rect 2906 37856 2918 37859
rect 5166 37856 5172 37868
rect 2906 37828 5172 37856
rect 2906 37825 2918 37828
rect 2860 37819 2918 37825
rect 5166 37816 5172 37828
rect 5224 37816 5230 37868
rect 14476 37865 14504 37896
rect 14461 37859 14519 37865
rect 14461 37825 14473 37859
rect 14507 37825 14519 37859
rect 14461 37819 14519 37825
rect 14728 37859 14786 37865
rect 14728 37825 14740 37859
rect 14774 37856 14786 37859
rect 15286 37856 15292 37868
rect 14774 37828 15292 37856
rect 14774 37825 14786 37828
rect 14728 37819 14786 37825
rect 15286 37816 15292 37828
rect 15344 37816 15350 37868
rect 2593 37791 2651 37797
rect 2593 37757 2605 37791
rect 2639 37757 2651 37791
rect 2593 37751 2651 37757
rect 4433 37791 4491 37797
rect 4433 37757 4445 37791
rect 4479 37757 4491 37791
rect 4433 37751 4491 37757
rect 2608 37652 2636 37751
rect 4448 37652 4476 37751
rect 6638 37748 6644 37800
rect 6696 37788 6702 37800
rect 8389 37791 8447 37797
rect 8389 37788 8401 37791
rect 6696 37760 8401 37788
rect 6696 37748 6702 37760
rect 8389 37757 8401 37760
rect 8435 37757 8447 37791
rect 8389 37751 8447 37757
rect 11514 37748 11520 37800
rect 11572 37788 11578 37800
rect 11793 37791 11851 37797
rect 11793 37788 11805 37791
rect 11572 37760 11805 37788
rect 11572 37748 11578 37760
rect 11793 37757 11805 37760
rect 11839 37757 11851 37791
rect 16546 37788 16574 37896
rect 16936 37893 16948 37927
rect 16982 37924 16994 37927
rect 17862 37924 17868 37936
rect 16982 37896 17868 37924
rect 16982 37893 16994 37896
rect 16936 37887 16994 37893
rect 17862 37884 17868 37896
rect 17920 37884 17926 37936
rect 18776 37927 18834 37933
rect 18776 37893 18788 37927
rect 18822 37924 18834 37927
rect 20622 37924 20628 37936
rect 18822 37896 20628 37924
rect 18822 37893 18834 37896
rect 18776 37887 18834 37893
rect 20622 37884 20628 37896
rect 20680 37884 20686 37936
rect 24394 37924 24400 37936
rect 23676 37896 24400 37924
rect 18506 37856 18512 37868
rect 18467 37828 18512 37856
rect 18506 37816 18512 37828
rect 18564 37816 18570 37868
rect 21818 37856 21824 37868
rect 21779 37828 21824 37856
rect 21818 37816 21824 37828
rect 21876 37816 21882 37868
rect 22088 37859 22146 37865
rect 22088 37825 22100 37859
rect 22134 37856 22146 37859
rect 23198 37856 23204 37868
rect 22134 37828 23204 37856
rect 22134 37825 22146 37828
rect 22088 37819 22146 37825
rect 23198 37816 23204 37828
rect 23256 37816 23262 37868
rect 23676 37865 23704 37896
rect 24394 37884 24400 37896
rect 24452 37884 24458 37936
rect 27424 37927 27482 37933
rect 27424 37893 27436 37927
rect 27470 37924 27482 37927
rect 27614 37924 27620 37936
rect 27470 37896 27620 37924
rect 27470 37893 27482 37896
rect 27424 37887 27482 37893
rect 27614 37884 27620 37896
rect 27672 37884 27678 37936
rect 34698 37924 34704 37936
rect 32140 37896 34704 37924
rect 23661 37859 23719 37865
rect 23661 37825 23673 37859
rect 23707 37825 23719 37859
rect 23661 37819 23719 37825
rect 23928 37859 23986 37865
rect 23928 37825 23940 37859
rect 23974 37856 23986 37859
rect 24946 37856 24952 37868
rect 23974 37828 24952 37856
rect 23974 37825 23986 37828
rect 23928 37819 23986 37825
rect 24946 37816 24952 37828
rect 25004 37816 25010 37868
rect 29356 37859 29414 37865
rect 29356 37825 29368 37859
rect 29402 37856 29414 37859
rect 30926 37856 30932 37868
rect 29402 37828 30932 37856
rect 29402 37825 29414 37828
rect 29356 37819 29414 37825
rect 30926 37816 30932 37828
rect 30984 37816 30990 37868
rect 16666 37788 16672 37800
rect 16546 37760 16672 37788
rect 11793 37751 11851 37757
rect 16666 37748 16672 37760
rect 16724 37748 16730 37800
rect 26234 37748 26240 37800
rect 26292 37788 26298 37800
rect 27157 37791 27215 37797
rect 27157 37788 27169 37791
rect 26292 37760 27169 37788
rect 26292 37748 26298 37760
rect 27157 37757 27169 37760
rect 27203 37757 27215 37791
rect 29086 37788 29092 37800
rect 29047 37760 29092 37788
rect 27157 37751 27215 37757
rect 29086 37748 29092 37760
rect 29144 37748 29150 37800
rect 31754 37748 31760 37800
rect 31812 37788 31818 37800
rect 32140 37797 32168 37896
rect 32392 37859 32450 37865
rect 32392 37825 32404 37859
rect 32438 37856 32450 37859
rect 33134 37856 33140 37868
rect 32438 37828 33140 37856
rect 32438 37825 32450 37828
rect 32392 37819 32450 37825
rect 33134 37816 33140 37828
rect 33192 37816 33198 37868
rect 33980 37865 34008 37896
rect 34698 37884 34704 37896
rect 34756 37884 34762 37936
rect 38746 37924 38752 37936
rect 37292 37896 38752 37924
rect 33965 37859 34023 37865
rect 33965 37825 33977 37859
rect 34011 37825 34023 37859
rect 33965 37819 34023 37825
rect 34232 37859 34290 37865
rect 34232 37825 34244 37859
rect 34278 37856 34290 37859
rect 35342 37856 35348 37868
rect 34278 37828 35348 37856
rect 34278 37825 34290 37828
rect 34232 37819 34290 37825
rect 35342 37816 35348 37828
rect 35400 37816 35406 37868
rect 37292 37865 37320 37896
rect 38746 37884 38752 37896
rect 38804 37924 38810 37936
rect 49228 37927 49286 37933
rect 38804 37896 39160 37924
rect 38804 37884 38810 37896
rect 39132 37868 39160 37896
rect 43088 37896 45554 37924
rect 37277 37859 37335 37865
rect 37277 37825 37289 37859
rect 37323 37825 37335 37859
rect 37277 37819 37335 37825
rect 37544 37859 37602 37865
rect 37544 37825 37556 37859
rect 37590 37856 37602 37859
rect 38654 37856 38660 37868
rect 37590 37828 38660 37856
rect 37590 37825 37602 37828
rect 37544 37819 37602 37825
rect 38654 37816 38660 37828
rect 38712 37816 38718 37868
rect 39114 37856 39120 37868
rect 39027 37828 39120 37856
rect 39114 37816 39120 37828
rect 39172 37816 39178 37868
rect 39390 37865 39396 37868
rect 39384 37819 39396 37865
rect 39448 37856 39454 37868
rect 43088 37865 43116 37896
rect 43073 37859 43131 37865
rect 39448 37828 39484 37856
rect 39390 37816 39396 37819
rect 39448 37816 39454 37828
rect 43073 37825 43085 37859
rect 43119 37825 43131 37859
rect 43073 37819 43131 37825
rect 43340 37859 43398 37865
rect 43340 37825 43352 37859
rect 43386 37856 43398 37859
rect 44450 37856 44456 37868
rect 43386 37828 44456 37856
rect 43386 37825 43398 37828
rect 43340 37819 43398 37825
rect 44450 37816 44456 37828
rect 44508 37816 44514 37868
rect 45526 37800 45554 37896
rect 49228 37893 49240 37927
rect 49274 37924 49286 37927
rect 49878 37924 49884 37936
rect 49274 37896 49884 37924
rect 49274 37893 49286 37896
rect 49228 37887 49286 37893
rect 49878 37884 49884 37896
rect 49936 37884 49942 37936
rect 51068 37927 51126 37933
rect 51068 37893 51080 37927
rect 51114 37924 51126 37927
rect 52270 37924 52276 37936
rect 51114 37896 52276 37924
rect 51114 37893 51126 37896
rect 51068 37887 51126 37893
rect 52270 37884 52276 37896
rect 52328 37884 52334 37936
rect 54662 37884 54668 37936
rect 54720 37924 54726 37936
rect 54757 37927 54815 37933
rect 54757 37924 54769 37927
rect 54720 37896 54769 37924
rect 54720 37884 54726 37896
rect 54757 37893 54769 37896
rect 54803 37893 54815 37927
rect 54757 37887 54815 37893
rect 45824 37859 45882 37865
rect 45824 37825 45836 37859
rect 45870 37856 45882 37859
rect 47118 37856 47124 37868
rect 45870 37828 47124 37856
rect 45870 37825 45882 37828
rect 45824 37819 45882 37825
rect 47118 37816 47124 37828
rect 47176 37816 47182 37868
rect 47486 37816 47492 37868
rect 47544 37856 47550 37868
rect 48222 37856 48228 37868
rect 47544 37828 48228 37856
rect 47544 37816 47550 37828
rect 48222 37816 48228 37828
rect 48280 37856 48286 37868
rect 48961 37859 49019 37865
rect 48961 37856 48973 37859
rect 48280 37828 48973 37856
rect 48280 37816 48286 37828
rect 48961 37825 48973 37828
rect 49007 37825 49019 37859
rect 48961 37819 49019 37825
rect 32125 37791 32183 37797
rect 32125 37788 32137 37791
rect 31812 37760 32137 37788
rect 31812 37748 31818 37760
rect 32125 37757 32137 37760
rect 32171 37757 32183 37791
rect 45526 37760 45560 37800
rect 32125 37751 32183 37757
rect 45554 37748 45560 37760
rect 45612 37788 45618 37800
rect 50798 37788 50804 37800
rect 45612 37760 45657 37788
rect 50759 37760 50804 37788
rect 45612 37748 45618 37760
rect 50798 37748 50804 37760
rect 50856 37748 50862 37800
rect 4614 37652 4620 37664
rect 2608 37624 4620 37652
rect 4614 37612 4620 37624
rect 4672 37612 4678 37664
rect 9766 37652 9772 37664
rect 9727 37624 9772 37652
rect 9766 37612 9772 37624
rect 9824 37612 9830 37664
rect 13170 37652 13176 37664
rect 13131 37624 13176 37652
rect 13170 37612 13176 37624
rect 13228 37612 13234 37664
rect 19886 37652 19892 37664
rect 19847 37624 19892 37652
rect 19886 37612 19892 37624
rect 19944 37612 19950 37664
rect 22094 37612 22100 37664
rect 22152 37652 22158 37664
rect 23201 37655 23259 37661
rect 23201 37652 23213 37655
rect 22152 37624 23213 37652
rect 22152 37612 22158 37624
rect 23201 37621 23213 37624
rect 23247 37621 23259 37655
rect 25038 37652 25044 37664
rect 24999 37624 25044 37652
rect 23201 37615 23259 37621
rect 25038 37612 25044 37624
rect 25096 37612 25102 37664
rect 38657 37655 38715 37661
rect 38657 37621 38669 37655
rect 38703 37652 38715 37655
rect 38746 37652 38752 37664
rect 38703 37624 38752 37652
rect 38703 37621 38715 37624
rect 38657 37615 38715 37621
rect 38746 37612 38752 37624
rect 38804 37612 38810 37664
rect 40494 37652 40500 37664
rect 40455 37624 40500 37652
rect 40494 37612 40500 37624
rect 40552 37612 40558 37664
rect 46934 37652 46940 37664
rect 46895 37624 46940 37652
rect 46934 37612 46940 37624
rect 46992 37612 46998 37664
rect 49878 37612 49884 37664
rect 49936 37652 49942 37664
rect 50341 37655 50399 37661
rect 50341 37652 50353 37655
rect 49936 37624 50353 37652
rect 49936 37612 49942 37624
rect 50341 37621 50353 37624
rect 50387 37621 50399 37655
rect 52178 37652 52184 37664
rect 52139 37624 52184 37652
rect 50341 37615 50399 37621
rect 52178 37612 52184 37624
rect 52236 37612 52242 37664
rect 55306 37612 55312 37664
rect 55364 37652 55370 37664
rect 56045 37655 56103 37661
rect 56045 37652 56057 37655
rect 55364 37624 56057 37652
rect 55364 37612 55370 37624
rect 56045 37621 56057 37624
rect 56091 37621 56103 37655
rect 56045 37615 56103 37621
rect 1104 37562 59340 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 59340 37562
rect 1104 37488 59340 37510
rect 17954 37408 17960 37460
rect 18012 37448 18018 37460
rect 18049 37451 18107 37457
rect 18049 37448 18061 37451
rect 18012 37420 18061 37448
rect 18012 37408 18018 37420
rect 18049 37417 18061 37420
rect 18095 37417 18107 37451
rect 18049 37411 18107 37417
rect 22370 37408 22376 37460
rect 22428 37448 22434 37460
rect 22465 37451 22523 37457
rect 22465 37448 22477 37451
rect 22428 37420 22477 37448
rect 22428 37408 22434 37420
rect 22465 37417 22477 37420
rect 22511 37417 22523 37451
rect 22465 37411 22523 37417
rect 27617 37451 27675 37457
rect 27617 37417 27629 37451
rect 27663 37448 27675 37451
rect 27706 37448 27712 37460
rect 27663 37420 27712 37448
rect 27663 37417 27675 37420
rect 27617 37411 27675 37417
rect 27706 37408 27712 37420
rect 27764 37408 27770 37460
rect 30926 37448 30932 37460
rect 30887 37420 30932 37448
rect 30926 37408 30932 37420
rect 30984 37408 30990 37460
rect 33134 37448 33140 37460
rect 33095 37420 33140 37448
rect 33134 37408 33140 37420
rect 33192 37408 33198 37460
rect 37550 37408 37556 37460
rect 37608 37448 37614 37460
rect 37921 37451 37979 37457
rect 37921 37448 37933 37451
rect 37608 37420 37933 37448
rect 37608 37408 37614 37420
rect 37921 37417 37933 37420
rect 37967 37417 37979 37451
rect 37921 37411 37979 37417
rect 42426 37408 42432 37460
rect 42484 37448 42490 37460
rect 42521 37451 42579 37457
rect 42521 37448 42533 37451
rect 42484 37420 42533 37448
rect 42484 37408 42490 37420
rect 42521 37417 42533 37420
rect 42567 37417 42579 37451
rect 55306 37448 55312 37460
rect 42521 37411 42579 37417
rect 55186 37420 55312 37448
rect 8938 37312 8944 37324
rect 8899 37284 8944 37312
rect 8938 37272 8944 37284
rect 8996 37272 9002 37324
rect 14734 37272 14740 37324
rect 14792 37312 14798 37324
rect 14829 37315 14887 37321
rect 14829 37312 14841 37315
rect 14792 37284 14841 37312
rect 14792 37272 14798 37284
rect 14829 37281 14841 37284
rect 14875 37281 14887 37315
rect 34698 37312 34704 37324
rect 34659 37284 34704 37312
rect 14829 37275 14887 37281
rect 34698 37272 34704 37284
rect 34756 37272 34762 37324
rect 48222 37312 48228 37324
rect 48183 37284 48228 37312
rect 48222 37272 48228 37284
rect 48280 37272 48286 37324
rect 4982 37204 4988 37256
rect 5040 37244 5046 37256
rect 5169 37247 5227 37253
rect 5169 37244 5181 37247
rect 5040 37216 5181 37244
rect 5040 37204 5046 37216
rect 5169 37213 5181 37216
rect 5215 37244 5227 37247
rect 6822 37244 6828 37256
rect 5215 37216 6828 37244
rect 5215 37213 5227 37216
rect 5169 37207 5227 37213
rect 6822 37204 6828 37216
rect 6880 37244 6886 37256
rect 7009 37247 7067 37253
rect 7009 37244 7021 37247
rect 6880 37216 7021 37244
rect 6880 37204 6886 37216
rect 7009 37213 7021 37216
rect 7055 37213 7067 37247
rect 7009 37207 7067 37213
rect 9208 37247 9266 37253
rect 9208 37213 9220 37247
rect 9254 37244 9266 37247
rect 9766 37244 9772 37256
rect 9254 37216 9772 37244
rect 9254 37213 9266 37216
rect 9208 37207 9266 37213
rect 9766 37204 9772 37216
rect 9824 37204 9830 37256
rect 11514 37244 11520 37256
rect 10152 37216 11520 37244
rect 5436 37179 5494 37185
rect 5436 37145 5448 37179
rect 5482 37176 5494 37179
rect 6730 37176 6736 37188
rect 5482 37148 6736 37176
rect 5482 37145 5494 37148
rect 5436 37139 5494 37145
rect 6730 37136 6736 37148
rect 6788 37136 6794 37188
rect 7276 37179 7334 37185
rect 7276 37145 7288 37179
rect 7322 37176 7334 37179
rect 9674 37176 9680 37188
rect 7322 37148 9680 37176
rect 7322 37145 7334 37148
rect 7276 37139 7334 37145
rect 9674 37136 9680 37148
rect 9732 37136 9738 37188
rect 6546 37108 6552 37120
rect 6507 37080 6552 37108
rect 6546 37068 6552 37080
rect 6604 37068 6610 37120
rect 8389 37111 8447 37117
rect 8389 37077 8401 37111
rect 8435 37108 8447 37111
rect 9030 37108 9036 37120
rect 8435 37080 9036 37108
rect 8435 37077 8447 37080
rect 8389 37071 8447 37077
rect 9030 37068 9036 37080
rect 9088 37068 9094 37120
rect 9122 37068 9128 37120
rect 9180 37108 9186 37120
rect 10152 37108 10180 37216
rect 11514 37204 11520 37216
rect 11572 37204 11578 37256
rect 11784 37247 11842 37253
rect 11784 37213 11796 37247
rect 11830 37244 11842 37247
rect 13170 37244 13176 37256
rect 11830 37216 13176 37244
rect 11830 37213 11842 37216
rect 11784 37207 11842 37213
rect 13170 37204 13176 37216
rect 13228 37204 13234 37256
rect 16666 37244 16672 37256
rect 16627 37216 16672 37244
rect 16666 37204 16672 37216
rect 16724 37204 16730 37256
rect 16942 37253 16948 37256
rect 16936 37207 16948 37253
rect 17000 37244 17006 37256
rect 19245 37247 19303 37253
rect 17000 37216 17036 37244
rect 16942 37204 16948 37207
rect 17000 37204 17006 37216
rect 19245 37213 19257 37247
rect 19291 37213 19303 37247
rect 19245 37207 19303 37213
rect 19512 37247 19570 37253
rect 19512 37213 19524 37247
rect 19558 37244 19570 37247
rect 19886 37244 19892 37256
rect 19558 37216 19892 37244
rect 19558 37213 19570 37216
rect 19512 37207 19570 37213
rect 15096 37179 15154 37185
rect 15096 37145 15108 37179
rect 15142 37176 15154 37179
rect 15286 37176 15292 37188
rect 15142 37148 15292 37176
rect 15142 37145 15154 37148
rect 15096 37139 15154 37145
rect 15286 37136 15292 37148
rect 15344 37136 15350 37188
rect 19260 37176 19288 37207
rect 19886 37204 19892 37216
rect 19944 37204 19950 37256
rect 21082 37244 21088 37256
rect 19987 37216 21088 37244
rect 19987 37176 20015 37216
rect 21082 37204 21088 37216
rect 21140 37204 21146 37256
rect 24394 37244 24400 37256
rect 24307 37216 24400 37244
rect 24394 37204 24400 37216
rect 24452 37204 24458 37256
rect 24664 37247 24722 37253
rect 24664 37213 24676 37247
rect 24710 37244 24722 37247
rect 25038 37244 25044 37256
rect 24710 37216 25044 37244
rect 24710 37213 24722 37216
rect 24664 37207 24722 37213
rect 25038 37204 25044 37216
rect 25096 37204 25102 37256
rect 26226 37247 26284 37253
rect 26226 37244 26238 37247
rect 26206 37213 26238 37244
rect 26272 37213 26284 37247
rect 26206 37207 26284 37213
rect 19260 37148 20015 37176
rect 20254 37136 20260 37188
rect 20312 37176 20318 37188
rect 21330 37179 21388 37185
rect 21330 37176 21342 37179
rect 20312 37148 21342 37176
rect 20312 37136 20318 37148
rect 21330 37145 21342 37148
rect 21376 37145 21388 37179
rect 24412 37176 24440 37204
rect 26206 37176 26234 37207
rect 26326 37204 26332 37256
rect 26384 37244 26390 37256
rect 26493 37247 26551 37253
rect 26493 37244 26505 37247
rect 26384 37216 26505 37244
rect 26384 37204 26390 37216
rect 26493 37213 26505 37216
rect 26539 37213 26551 37247
rect 29546 37244 29552 37256
rect 29507 37216 29552 37244
rect 26493 37207 26551 37213
rect 29546 37204 29552 37216
rect 29604 37204 29610 37256
rect 29638 37204 29644 37256
rect 29696 37244 29702 37256
rect 29805 37247 29863 37253
rect 29805 37244 29817 37247
rect 29696 37216 29817 37244
rect 29696 37204 29702 37216
rect 29805 37213 29817 37216
rect 29851 37213 29863 37247
rect 31754 37244 31760 37256
rect 31715 37216 31760 37244
rect 29805 37207 29863 37213
rect 31754 37204 31760 37216
rect 31812 37204 31818 37256
rect 34790 37204 34796 37256
rect 34848 37244 34854 37256
rect 34957 37247 35015 37253
rect 34957 37244 34969 37247
rect 34848 37216 34969 37244
rect 34848 37204 34854 37216
rect 34957 37213 34969 37216
rect 35003 37213 35015 37247
rect 34957 37207 35015 37213
rect 35434 37204 35440 37256
rect 35492 37244 35498 37256
rect 36541 37247 36599 37253
rect 36541 37244 36553 37247
rect 35492 37216 36553 37244
rect 35492 37204 35498 37216
rect 36541 37213 36553 37216
rect 36587 37213 36599 37247
rect 36541 37207 36599 37213
rect 36630 37204 36636 37256
rect 36688 37244 36694 37256
rect 36797 37247 36855 37253
rect 36797 37244 36809 37247
rect 36688 37216 36809 37244
rect 36688 37204 36694 37216
rect 36797 37213 36809 37216
rect 36843 37213 36855 37247
rect 36797 37207 36855 37213
rect 40402 37204 40408 37256
rect 40460 37244 40466 37256
rect 41233 37247 41291 37253
rect 41233 37244 41245 37247
rect 40460 37216 41245 37244
rect 40460 37204 40466 37216
rect 41233 37213 41245 37216
rect 41279 37213 41291 37247
rect 41233 37207 41291 37213
rect 45554 37204 45560 37256
rect 45612 37244 45618 37256
rect 46385 37247 46443 37253
rect 46385 37244 46397 37247
rect 45612 37216 46397 37244
rect 45612 37204 45618 37216
rect 46385 37213 46397 37216
rect 46431 37213 46443 37247
rect 46385 37207 46443 37213
rect 46652 37247 46710 37253
rect 46652 37213 46664 37247
rect 46698 37244 46710 37247
rect 47026 37244 47032 37256
rect 46698 37216 47032 37244
rect 46698 37213 46710 37216
rect 46652 37207 46710 37213
rect 47026 37204 47032 37216
rect 47084 37204 47090 37256
rect 51537 37247 51595 37253
rect 51537 37213 51549 37247
rect 51583 37244 51595 37247
rect 53377 37247 53435 37253
rect 53377 37244 53389 37247
rect 51583 37216 53389 37244
rect 51583 37213 51595 37216
rect 51537 37207 51595 37213
rect 53377 37213 53389 37216
rect 53423 37244 53435 37247
rect 55186 37244 55214 37420
rect 55306 37408 55312 37420
rect 55364 37408 55370 37460
rect 56686 37448 56692 37460
rect 56647 37420 56692 37448
rect 56686 37408 56692 37420
rect 56744 37408 56750 37460
rect 55306 37244 55312 37256
rect 53423 37216 55214 37244
rect 55267 37216 55312 37244
rect 53423 37213 53435 37216
rect 53377 37207 53435 37213
rect 55306 37204 55312 37216
rect 55364 37204 55370 37256
rect 24412 37148 26234 37176
rect 21330 37139 21388 37145
rect 26206 37120 26234 37148
rect 32024 37179 32082 37185
rect 32024 37145 32036 37179
rect 32070 37176 32082 37179
rect 33502 37176 33508 37188
rect 32070 37148 33508 37176
rect 32070 37145 32082 37148
rect 32024 37139 32082 37145
rect 33502 37136 33508 37148
rect 33560 37136 33566 37188
rect 48492 37179 48550 37185
rect 48492 37145 48504 37179
rect 48538 37176 48550 37179
rect 50154 37176 50160 37188
rect 48538 37148 50160 37176
rect 48538 37145 48550 37148
rect 48492 37139 48550 37145
rect 50154 37136 50160 37148
rect 50212 37136 50218 37188
rect 51804 37179 51862 37185
rect 51804 37145 51816 37179
rect 51850 37176 51862 37179
rect 53644 37179 53702 37185
rect 51850 37148 53604 37176
rect 51850 37145 51862 37148
rect 51804 37139 51862 37145
rect 53576 37120 53604 37148
rect 53644 37145 53656 37179
rect 53690 37176 53702 37179
rect 53834 37176 53840 37188
rect 53690 37148 53840 37176
rect 53690 37145 53702 37148
rect 53644 37139 53702 37145
rect 53834 37136 53840 37148
rect 53892 37136 53898 37188
rect 55576 37179 55634 37185
rect 55576 37145 55588 37179
rect 55622 37176 55634 37179
rect 56410 37176 56416 37188
rect 55622 37148 56416 37176
rect 55622 37145 55634 37148
rect 55576 37139 55634 37145
rect 56410 37136 56416 37148
rect 56468 37136 56474 37188
rect 10318 37108 10324 37120
rect 9180 37080 10180 37108
rect 10279 37080 10324 37108
rect 9180 37068 9186 37080
rect 10318 37068 10324 37080
rect 10376 37068 10382 37120
rect 12894 37108 12900 37120
rect 12855 37080 12900 37108
rect 12894 37068 12900 37080
rect 12952 37068 12958 37120
rect 15654 37068 15660 37120
rect 15712 37108 15718 37120
rect 16209 37111 16267 37117
rect 16209 37108 16221 37111
rect 15712 37080 16221 37108
rect 15712 37068 15718 37080
rect 16209 37077 16221 37080
rect 16255 37077 16267 37111
rect 20622 37108 20628 37120
rect 20583 37080 20628 37108
rect 16209 37071 16267 37077
rect 20622 37068 20628 37080
rect 20680 37068 20686 37120
rect 25774 37108 25780 37120
rect 25735 37080 25780 37108
rect 25774 37068 25780 37080
rect 25832 37068 25838 37120
rect 26206 37080 26240 37120
rect 26234 37068 26240 37080
rect 26292 37068 26298 37120
rect 35342 37068 35348 37120
rect 35400 37108 35406 37120
rect 36081 37111 36139 37117
rect 36081 37108 36093 37111
rect 35400 37080 36093 37108
rect 35400 37068 35406 37080
rect 36081 37077 36093 37080
rect 36127 37077 36139 37111
rect 47762 37108 47768 37120
rect 47723 37080 47768 37108
rect 36081 37071 36139 37077
rect 47762 37068 47768 37080
rect 47820 37068 47826 37120
rect 49605 37111 49663 37117
rect 49605 37077 49617 37111
rect 49651 37108 49663 37111
rect 50062 37108 50068 37120
rect 49651 37080 50068 37108
rect 49651 37077 49663 37080
rect 49605 37071 49663 37077
rect 50062 37068 50068 37080
rect 50120 37068 50126 37120
rect 52822 37068 52828 37120
rect 52880 37108 52886 37120
rect 52917 37111 52975 37117
rect 52917 37108 52929 37111
rect 52880 37080 52929 37108
rect 52880 37068 52886 37080
rect 52917 37077 52929 37080
rect 52963 37077 52975 37111
rect 52917 37071 52975 37077
rect 53558 37068 53564 37120
rect 53616 37068 53622 37120
rect 53742 37068 53748 37120
rect 53800 37108 53806 37120
rect 54757 37111 54815 37117
rect 54757 37108 54769 37111
rect 53800 37080 54769 37108
rect 53800 37068 53806 37080
rect 54757 37077 54769 37080
rect 54803 37077 54815 37111
rect 54757 37071 54815 37077
rect 1104 37018 59340 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 59340 37018
rect 1104 36944 59340 36966
rect 5810 36904 5816 36916
rect 5771 36876 5816 36904
rect 5810 36864 5816 36876
rect 5868 36864 5874 36916
rect 9674 36864 9680 36916
rect 9732 36904 9738 36916
rect 9769 36907 9827 36913
rect 9769 36904 9781 36907
rect 9732 36876 9781 36904
rect 9732 36864 9738 36876
rect 9769 36873 9781 36876
rect 9815 36873 9827 36907
rect 9769 36867 9827 36873
rect 14734 36864 14740 36916
rect 14792 36904 14798 36916
rect 14829 36907 14887 36913
rect 14829 36904 14841 36907
rect 14792 36876 14841 36904
rect 14792 36864 14798 36876
rect 14829 36873 14841 36876
rect 14875 36873 14887 36907
rect 14829 36867 14887 36873
rect 18049 36907 18107 36913
rect 18049 36873 18061 36907
rect 18095 36904 18107 36907
rect 19426 36904 19432 36916
rect 18095 36876 19432 36904
rect 18095 36873 18107 36876
rect 18049 36867 18107 36873
rect 19426 36864 19432 36876
rect 19484 36864 19490 36916
rect 20254 36904 20260 36916
rect 20215 36876 20260 36904
rect 20254 36864 20260 36876
rect 20312 36864 20318 36916
rect 23198 36904 23204 36916
rect 23159 36876 23204 36904
rect 23198 36864 23204 36876
rect 23256 36864 23262 36916
rect 24946 36864 24952 36916
rect 25004 36904 25010 36916
rect 25041 36907 25099 36913
rect 25041 36904 25053 36907
rect 25004 36876 25053 36904
rect 25004 36864 25010 36876
rect 25041 36873 25053 36876
rect 25087 36873 25099 36907
rect 33502 36904 33508 36916
rect 33463 36876 33508 36904
rect 25041 36867 25099 36873
rect 33502 36864 33508 36876
rect 33560 36864 33566 36916
rect 38654 36904 38660 36916
rect 38615 36876 38660 36904
rect 38654 36864 38660 36876
rect 38712 36864 38718 36916
rect 50154 36864 50160 36916
rect 50212 36904 50218 36916
rect 50341 36907 50399 36913
rect 50341 36904 50353 36907
rect 50212 36876 50353 36904
rect 50212 36864 50218 36876
rect 50341 36873 50353 36876
rect 50387 36873 50399 36907
rect 56410 36904 56416 36916
rect 56371 36876 56416 36904
rect 50341 36867 50399 36873
rect 56410 36864 56416 36876
rect 56468 36864 56474 36916
rect 4700 36839 4758 36845
rect 4700 36805 4712 36839
rect 4746 36836 4758 36839
rect 6546 36836 6552 36848
rect 4746 36808 6552 36836
rect 4746 36805 4758 36808
rect 4700 36799 4758 36805
rect 6546 36796 6552 36808
rect 6604 36796 6610 36848
rect 6816 36839 6874 36845
rect 6816 36805 6828 36839
rect 6862 36836 6874 36839
rect 8478 36836 8484 36848
rect 6862 36808 8484 36836
rect 6862 36805 6874 36808
rect 6816 36799 6874 36805
rect 8478 36796 8484 36808
rect 8536 36796 8542 36848
rect 8656 36839 8714 36845
rect 8656 36805 8668 36839
rect 8702 36836 8714 36839
rect 10318 36836 10324 36848
rect 8702 36808 10324 36836
rect 8702 36805 8714 36808
rect 8656 36799 8714 36805
rect 10318 36796 10324 36808
rect 10376 36796 10382 36848
rect 11784 36839 11842 36845
rect 11784 36805 11796 36839
rect 11830 36836 11842 36839
rect 12894 36836 12900 36848
rect 11830 36808 12900 36836
rect 11830 36805 11842 36808
rect 11784 36799 11842 36805
rect 12894 36796 12900 36808
rect 12952 36796 12958 36848
rect 13354 36796 13360 36848
rect 13412 36836 13418 36848
rect 13541 36839 13599 36845
rect 13541 36836 13553 36839
rect 13412 36808 13553 36836
rect 13412 36796 13418 36808
rect 13541 36805 13553 36808
rect 13587 36805 13599 36839
rect 19144 36839 19202 36845
rect 13541 36799 13599 36805
rect 16684 36808 18920 36836
rect 16684 36780 16712 36808
rect 4433 36771 4491 36777
rect 4433 36737 4445 36771
rect 4479 36768 4491 36771
rect 4522 36768 4528 36780
rect 4479 36740 4528 36768
rect 4479 36737 4491 36740
rect 4433 36731 4491 36737
rect 4522 36728 4528 36740
rect 4580 36768 4586 36780
rect 4982 36768 4988 36780
rect 4580 36740 4988 36768
rect 4580 36728 4586 36740
rect 4982 36728 4988 36740
rect 5040 36728 5046 36780
rect 6638 36728 6644 36780
rect 6696 36728 6702 36780
rect 11514 36768 11520 36780
rect 11475 36740 11520 36768
rect 11514 36728 11520 36740
rect 11572 36728 11578 36780
rect 16666 36768 16672 36780
rect 16579 36740 16672 36768
rect 16666 36728 16672 36740
rect 16724 36728 16730 36780
rect 16936 36771 16994 36777
rect 16936 36737 16948 36771
rect 16982 36768 16994 36771
rect 18046 36768 18052 36780
rect 16982 36740 18052 36768
rect 16982 36737 16994 36740
rect 16936 36731 16994 36737
rect 18046 36728 18052 36740
rect 18104 36728 18110 36780
rect 18892 36777 18920 36808
rect 19144 36805 19156 36839
rect 19190 36836 19202 36839
rect 20622 36836 20628 36848
rect 19190 36808 20628 36836
rect 19190 36805 19202 36808
rect 19144 36799 19202 36805
rect 20622 36796 20628 36808
rect 20680 36796 20686 36848
rect 27338 36836 27344 36848
rect 27299 36808 27344 36836
rect 27338 36796 27344 36808
rect 27396 36796 27402 36848
rect 35612 36839 35670 36845
rect 35612 36805 35624 36839
rect 35658 36836 35670 36839
rect 37544 36839 37602 36845
rect 35658 36808 37412 36836
rect 35658 36805 35670 36808
rect 35612 36799 35670 36805
rect 18877 36771 18935 36777
rect 18877 36737 18889 36771
rect 18923 36768 18935 36771
rect 21082 36768 21088 36780
rect 18923 36740 21088 36768
rect 18923 36737 18935 36740
rect 18877 36731 18935 36737
rect 21082 36728 21088 36740
rect 21140 36768 21146 36780
rect 21821 36771 21879 36777
rect 21821 36768 21833 36771
rect 21140 36740 21833 36768
rect 21140 36728 21146 36740
rect 21821 36737 21833 36740
rect 21867 36737 21879 36771
rect 21821 36731 21879 36737
rect 22088 36771 22146 36777
rect 22088 36737 22100 36771
rect 22134 36768 22146 36771
rect 22462 36768 22468 36780
rect 22134 36740 22468 36768
rect 22134 36737 22146 36740
rect 22088 36731 22146 36737
rect 22462 36728 22468 36740
rect 22520 36728 22526 36780
rect 23928 36771 23986 36777
rect 23928 36737 23940 36771
rect 23974 36768 23986 36771
rect 25038 36768 25044 36780
rect 23974 36740 25044 36768
rect 23974 36737 23986 36740
rect 23928 36731 23986 36737
rect 25038 36728 25044 36740
rect 25096 36728 25102 36780
rect 29086 36728 29092 36780
rect 29144 36768 29150 36780
rect 29549 36771 29607 36777
rect 29549 36768 29561 36771
rect 29144 36740 29561 36768
rect 29144 36728 29150 36740
rect 29549 36737 29561 36740
rect 29595 36737 29607 36771
rect 29549 36731 29607 36737
rect 29816 36771 29874 36777
rect 29816 36737 29828 36771
rect 29862 36768 29874 36771
rect 30926 36768 30932 36780
rect 29862 36740 30932 36768
rect 29862 36737 29874 36740
rect 29816 36731 29874 36737
rect 30926 36728 30932 36740
rect 30984 36728 30990 36780
rect 32392 36771 32450 36777
rect 32392 36737 32404 36771
rect 32438 36768 32450 36771
rect 33502 36768 33508 36780
rect 32438 36740 33508 36768
rect 32438 36737 32450 36740
rect 32392 36731 32450 36737
rect 33502 36728 33508 36740
rect 33560 36728 33566 36780
rect 35345 36771 35403 36777
rect 35345 36737 35357 36771
rect 35391 36768 35403 36771
rect 35434 36768 35440 36780
rect 35391 36740 35440 36768
rect 35391 36737 35403 36740
rect 35345 36731 35403 36737
rect 35434 36728 35440 36740
rect 35492 36768 35498 36780
rect 37277 36771 37335 36777
rect 37277 36768 37289 36771
rect 35492 36740 37289 36768
rect 35492 36728 35498 36740
rect 37277 36737 37289 36740
rect 37323 36737 37335 36771
rect 37384 36768 37412 36808
rect 37544 36805 37556 36839
rect 37590 36836 37602 36839
rect 37918 36836 37924 36848
rect 37590 36808 37924 36836
rect 37590 36805 37602 36808
rect 37544 36799 37602 36805
rect 37918 36796 37924 36808
rect 37976 36796 37982 36848
rect 45916 36839 45974 36845
rect 45916 36805 45928 36839
rect 45962 36836 45974 36839
rect 47762 36836 47768 36848
rect 45962 36808 47768 36836
rect 45962 36805 45974 36808
rect 45916 36799 45974 36805
rect 47762 36796 47768 36808
rect 47820 36796 47826 36848
rect 49228 36839 49286 36845
rect 49228 36805 49240 36839
rect 49274 36836 49286 36839
rect 49878 36836 49884 36848
rect 49274 36808 49884 36836
rect 49274 36805 49286 36808
rect 49228 36799 49286 36805
rect 49878 36796 49884 36808
rect 49936 36796 49942 36848
rect 51068 36839 51126 36845
rect 51068 36805 51080 36839
rect 51114 36836 51126 36839
rect 52178 36836 52184 36848
rect 51114 36808 52184 36836
rect 51114 36805 51126 36808
rect 51068 36799 51126 36805
rect 52178 36796 52184 36808
rect 52236 36796 52242 36848
rect 55214 36836 55220 36848
rect 55048 36808 55220 36836
rect 37384 36740 38323 36768
rect 37277 36731 37335 36737
rect 6549 36703 6607 36709
rect 6549 36669 6561 36703
rect 6595 36700 6607 36703
rect 6656 36700 6684 36728
rect 8386 36700 8392 36712
rect 6595 36672 6684 36700
rect 8347 36672 8392 36700
rect 6595 36669 6607 36672
rect 6549 36663 6607 36669
rect 8386 36660 8392 36672
rect 8444 36660 8450 36712
rect 23658 36700 23664 36712
rect 23619 36672 23664 36700
rect 23658 36660 23664 36672
rect 23716 36660 23722 36712
rect 31754 36660 31760 36712
rect 31812 36700 31818 36712
rect 32125 36703 32183 36709
rect 32125 36700 32137 36703
rect 31812 36672 32137 36700
rect 31812 36660 31818 36672
rect 32125 36669 32137 36672
rect 32171 36669 32183 36703
rect 38295 36700 38323 36740
rect 38654 36728 38660 36780
rect 38712 36768 38718 36780
rect 39373 36771 39431 36777
rect 39373 36768 39385 36771
rect 38712 36740 39385 36768
rect 38712 36728 38718 36740
rect 39373 36737 39385 36740
rect 39419 36737 39431 36771
rect 39373 36731 39431 36737
rect 42426 36728 42432 36780
rect 42484 36768 42490 36780
rect 43809 36771 43867 36777
rect 43809 36768 43821 36771
rect 42484 36740 43821 36768
rect 42484 36728 42490 36740
rect 43809 36737 43821 36740
rect 43855 36737 43867 36771
rect 43809 36731 43867 36737
rect 44076 36771 44134 36777
rect 44076 36737 44088 36771
rect 44122 36768 44134 36771
rect 46934 36768 46940 36780
rect 44122 36740 46940 36768
rect 44122 36737 44134 36740
rect 44076 36731 44134 36737
rect 46934 36728 46940 36740
rect 46992 36728 46998 36780
rect 50154 36728 50160 36780
rect 50212 36768 50218 36780
rect 50798 36768 50804 36780
rect 50212 36740 50804 36768
rect 50212 36728 50218 36740
rect 50798 36728 50804 36740
rect 50856 36728 50862 36780
rect 55048 36777 55076 36808
rect 55214 36796 55220 36808
rect 55272 36796 55278 36848
rect 55033 36771 55091 36777
rect 55033 36737 55045 36771
rect 55079 36737 55091 36771
rect 55033 36731 55091 36737
rect 55300 36771 55358 36777
rect 55300 36737 55312 36771
rect 55346 36768 55358 36771
rect 56686 36768 56692 36780
rect 55346 36740 56692 36768
rect 55346 36737 55358 36740
rect 55300 36731 55358 36737
rect 56686 36728 56692 36740
rect 56744 36728 56750 36780
rect 38838 36700 38844 36712
rect 38295 36672 38844 36700
rect 32125 36663 32183 36669
rect 38838 36660 38844 36672
rect 38896 36660 38902 36712
rect 39114 36700 39120 36712
rect 39075 36672 39120 36700
rect 39114 36660 39120 36672
rect 39172 36660 39178 36712
rect 45554 36660 45560 36712
rect 45612 36700 45618 36712
rect 45649 36703 45707 36709
rect 45649 36700 45661 36703
rect 45612 36672 45661 36700
rect 45612 36660 45618 36672
rect 45649 36669 45661 36672
rect 45695 36669 45707 36703
rect 45649 36663 45707 36669
rect 48222 36660 48228 36712
rect 48280 36700 48286 36712
rect 48961 36703 49019 36709
rect 48961 36700 48973 36703
rect 48280 36672 48973 36700
rect 48280 36660 48286 36672
rect 48961 36669 48973 36672
rect 49007 36669 49019 36703
rect 48961 36663 49019 36669
rect 52086 36592 52092 36644
rect 52144 36632 52150 36644
rect 52181 36635 52239 36641
rect 52181 36632 52193 36635
rect 52144 36604 52193 36632
rect 52144 36592 52150 36604
rect 52181 36601 52193 36604
rect 52227 36601 52239 36635
rect 52181 36595 52239 36601
rect 7926 36564 7932 36576
rect 7887 36536 7932 36564
rect 7926 36524 7932 36536
rect 7984 36524 7990 36576
rect 12894 36564 12900 36576
rect 12855 36536 12900 36564
rect 12894 36524 12900 36536
rect 12952 36524 12958 36576
rect 28813 36567 28871 36573
rect 28813 36533 28825 36567
rect 28859 36564 28871 36567
rect 28902 36564 28908 36576
rect 28859 36536 28908 36564
rect 28859 36533 28871 36536
rect 28813 36527 28871 36533
rect 28902 36524 28908 36536
rect 28960 36524 28966 36576
rect 29822 36524 29828 36576
rect 29880 36564 29886 36576
rect 30929 36567 30987 36573
rect 30929 36564 30941 36567
rect 29880 36536 30941 36564
rect 29880 36524 29886 36536
rect 30929 36533 30941 36536
rect 30975 36533 30987 36567
rect 36722 36564 36728 36576
rect 36683 36536 36728 36564
rect 30929 36527 30987 36533
rect 36722 36524 36728 36536
rect 36780 36524 36786 36576
rect 39482 36524 39488 36576
rect 39540 36564 39546 36576
rect 40497 36567 40555 36573
rect 40497 36564 40509 36567
rect 39540 36536 40509 36564
rect 39540 36524 39546 36536
rect 40497 36533 40509 36536
rect 40543 36533 40555 36567
rect 40497 36527 40555 36533
rect 45189 36567 45247 36573
rect 45189 36533 45201 36567
rect 45235 36564 45247 36567
rect 45646 36564 45652 36576
rect 45235 36536 45652 36564
rect 45235 36533 45247 36536
rect 45189 36527 45247 36533
rect 45646 36524 45652 36536
rect 45704 36524 45710 36576
rect 47026 36564 47032 36576
rect 46987 36536 47032 36564
rect 47026 36524 47032 36536
rect 47084 36524 47090 36576
rect 1104 36474 59340 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 59340 36474
rect 1104 36400 59340 36422
rect 8478 36320 8484 36372
rect 8536 36360 8542 36372
rect 10321 36363 10379 36369
rect 10321 36360 10333 36363
rect 8536 36332 10333 36360
rect 8536 36320 8542 36332
rect 10321 36329 10333 36332
rect 10367 36329 10379 36363
rect 18046 36360 18052 36372
rect 18007 36332 18052 36360
rect 10321 36323 10379 36329
rect 18046 36320 18052 36332
rect 18104 36320 18110 36372
rect 22462 36360 22468 36372
rect 22423 36332 22468 36360
rect 22462 36320 22468 36332
rect 22520 36320 22526 36372
rect 27617 36363 27675 36369
rect 27617 36329 27629 36363
rect 27663 36360 27675 36363
rect 27798 36360 27804 36372
rect 27663 36332 27804 36360
rect 27663 36329 27675 36332
rect 27617 36323 27675 36329
rect 27798 36320 27804 36332
rect 27856 36320 27862 36372
rect 30926 36360 30932 36372
rect 30887 36332 30932 36360
rect 30926 36320 30932 36332
rect 30984 36320 30990 36372
rect 31754 36320 31760 36372
rect 31812 36360 31818 36372
rect 33597 36363 33655 36369
rect 33597 36360 33609 36363
rect 31812 36332 33609 36360
rect 31812 36320 31818 36332
rect 33597 36329 33609 36332
rect 33643 36329 33655 36363
rect 38654 36360 38660 36372
rect 38615 36332 38660 36360
rect 33597 36323 33655 36329
rect 38654 36320 38660 36332
rect 38712 36320 38718 36372
rect 51442 36320 51448 36372
rect 51500 36360 51506 36372
rect 51537 36363 51595 36369
rect 51537 36360 51549 36363
rect 51500 36332 51549 36360
rect 51500 36320 51506 36332
rect 51537 36329 51549 36332
rect 51583 36329 51595 36363
rect 56686 36360 56692 36372
rect 56647 36332 56692 36360
rect 51537 36323 51595 36329
rect 56686 36320 56692 36332
rect 56744 36320 56750 36372
rect 8386 36184 8392 36236
rect 8444 36224 8450 36236
rect 8938 36224 8944 36236
rect 8444 36196 8944 36224
rect 8444 36184 8450 36196
rect 8938 36184 8944 36196
rect 8996 36184 9002 36236
rect 11514 36224 11520 36236
rect 11475 36196 11520 36224
rect 11514 36184 11520 36196
rect 11572 36184 11578 36236
rect 16666 36224 16672 36236
rect 16627 36196 16672 36224
rect 16666 36184 16672 36196
rect 16724 36184 16730 36236
rect 21082 36224 21088 36236
rect 21043 36196 21088 36224
rect 21082 36184 21088 36196
rect 21140 36184 21146 36236
rect 29086 36184 29092 36236
rect 29144 36224 29150 36236
rect 29549 36227 29607 36233
rect 29549 36224 29561 36227
rect 29144 36196 29561 36224
rect 29144 36184 29150 36196
rect 29549 36193 29561 36196
rect 29595 36193 29607 36227
rect 29549 36187 29607 36193
rect 6362 36116 6368 36168
rect 6420 36156 6426 36168
rect 6549 36159 6607 36165
rect 6549 36156 6561 36159
rect 6420 36128 6561 36156
rect 6420 36116 6426 36128
rect 6549 36125 6561 36128
rect 6595 36156 6607 36159
rect 6638 36156 6644 36168
rect 6595 36128 6644 36156
rect 6595 36125 6607 36128
rect 6549 36119 6607 36125
rect 6638 36116 6644 36128
rect 6696 36116 6702 36168
rect 6816 36159 6874 36165
rect 6816 36125 6828 36159
rect 6862 36156 6874 36159
rect 7926 36156 7932 36168
rect 6862 36128 7932 36156
rect 6862 36125 6874 36128
rect 6816 36119 6874 36125
rect 7926 36116 7932 36128
rect 7984 36116 7990 36168
rect 9030 36116 9036 36168
rect 9088 36156 9094 36168
rect 9197 36159 9255 36165
rect 9197 36156 9209 36159
rect 9088 36128 9209 36156
rect 9088 36116 9094 36128
rect 9197 36125 9209 36128
rect 9243 36125 9255 36159
rect 9197 36119 9255 36125
rect 11784 36159 11842 36165
rect 11784 36125 11796 36159
rect 11830 36156 11842 36159
rect 12894 36156 12900 36168
rect 11830 36128 12900 36156
rect 11830 36125 11842 36128
rect 11784 36119 11842 36125
rect 12894 36116 12900 36128
rect 12952 36116 12958 36168
rect 13998 36116 14004 36168
rect 14056 36156 14062 36168
rect 14093 36159 14151 36165
rect 14093 36156 14105 36159
rect 14056 36128 14105 36156
rect 14056 36116 14062 36128
rect 14093 36125 14105 36128
rect 14139 36156 14151 36159
rect 14734 36156 14740 36168
rect 14139 36128 14740 36156
rect 14139 36125 14151 36128
rect 14093 36119 14151 36125
rect 14734 36116 14740 36128
rect 14792 36116 14798 36168
rect 17862 36116 17868 36168
rect 17920 36156 17926 36168
rect 19245 36159 19303 36165
rect 19245 36156 19257 36159
rect 17920 36128 19257 36156
rect 17920 36116 17926 36128
rect 19245 36125 19257 36128
rect 19291 36125 19303 36159
rect 19245 36119 19303 36125
rect 21352 36159 21410 36165
rect 21352 36125 21364 36159
rect 21398 36156 21410 36159
rect 22186 36156 22192 36168
rect 21398 36128 22192 36156
rect 21398 36125 21410 36128
rect 21352 36119 21410 36125
rect 22186 36116 22192 36128
rect 22244 36116 22250 36168
rect 24394 36156 24400 36168
rect 24355 36128 24400 36156
rect 24394 36116 24400 36128
rect 24452 36116 24458 36168
rect 24664 36159 24722 36165
rect 24664 36125 24676 36159
rect 24710 36156 24722 36159
rect 25774 36156 25780 36168
rect 24710 36128 25780 36156
rect 24710 36125 24722 36128
rect 24664 36119 24722 36125
rect 25774 36116 25780 36128
rect 25832 36116 25838 36168
rect 26234 36116 26240 36168
rect 26292 36156 26298 36168
rect 27062 36156 27068 36168
rect 26292 36128 27068 36156
rect 26292 36116 26298 36128
rect 27062 36116 27068 36128
rect 27120 36116 27126 36168
rect 13814 36048 13820 36100
rect 13872 36088 13878 36100
rect 14338 36091 14396 36097
rect 14338 36088 14350 36091
rect 13872 36060 14350 36088
rect 13872 36048 13878 36060
rect 14338 36057 14350 36060
rect 14384 36057 14396 36091
rect 14338 36051 14396 36057
rect 16936 36091 16994 36097
rect 16936 36057 16948 36091
rect 16982 36088 16994 36091
rect 17770 36088 17776 36100
rect 16982 36060 17776 36088
rect 16982 36057 16994 36060
rect 16936 36051 16994 36057
rect 17770 36048 17776 36060
rect 17828 36048 17834 36100
rect 19512 36091 19570 36097
rect 19512 36057 19524 36091
rect 19558 36088 19570 36091
rect 20530 36088 20536 36100
rect 19558 36060 20536 36088
rect 19558 36057 19570 36060
rect 19512 36051 19570 36057
rect 20530 36048 20536 36060
rect 20588 36048 20594 36100
rect 26482 36091 26540 36097
rect 26482 36088 26494 36091
rect 26206 36060 26494 36088
rect 7926 36020 7932 36032
rect 7887 35992 7932 36020
rect 7926 35980 7932 35992
rect 7984 35980 7990 36032
rect 12894 36020 12900 36032
rect 12855 35992 12900 36020
rect 12894 35980 12900 35992
rect 12952 35980 12958 36032
rect 15194 35980 15200 36032
rect 15252 36020 15258 36032
rect 15473 36023 15531 36029
rect 15473 36020 15485 36023
rect 15252 35992 15485 36020
rect 15252 35980 15258 35992
rect 15473 35989 15485 35992
rect 15519 35989 15531 36023
rect 15473 35983 15531 35989
rect 20162 35980 20168 36032
rect 20220 36020 20226 36032
rect 20625 36023 20683 36029
rect 20625 36020 20637 36023
rect 20220 35992 20637 36020
rect 20220 35980 20226 35992
rect 20625 35989 20637 35992
rect 20671 35989 20683 36023
rect 20625 35983 20683 35989
rect 25777 36023 25835 36029
rect 25777 35989 25789 36023
rect 25823 36020 25835 36023
rect 26206 36020 26234 36060
rect 26482 36057 26494 36060
rect 26528 36057 26540 36091
rect 26482 36051 26540 36057
rect 25823 35992 26234 36020
rect 29564 36020 29592 36187
rect 39114 36184 39120 36236
rect 39172 36224 39178 36236
rect 39853 36227 39911 36233
rect 39853 36224 39865 36227
rect 39172 36196 39865 36224
rect 39172 36184 39178 36196
rect 39853 36193 39865 36196
rect 39899 36224 39911 36227
rect 39899 36196 39988 36224
rect 39899 36193 39911 36196
rect 39853 36187 39911 36193
rect 39960 36168 39988 36196
rect 46842 36184 46848 36236
rect 46900 36224 46906 36236
rect 48222 36224 48228 36236
rect 46900 36196 48228 36224
rect 46900 36184 46906 36196
rect 48222 36184 48228 36196
rect 48280 36184 48286 36236
rect 34606 36116 34612 36168
rect 34664 36156 34670 36168
rect 34885 36159 34943 36165
rect 34885 36156 34897 36159
rect 34664 36128 34897 36156
rect 34664 36116 34670 36128
rect 34885 36125 34897 36128
rect 34931 36156 34943 36159
rect 35434 36156 35440 36168
rect 34931 36128 35440 36156
rect 34931 36125 34943 36128
rect 34885 36119 34943 36125
rect 35434 36116 35440 36128
rect 35492 36156 35498 36168
rect 37277 36159 37335 36165
rect 37277 36156 37289 36159
rect 35492 36128 37289 36156
rect 35492 36116 35498 36128
rect 37277 36125 37289 36128
rect 37323 36125 37335 36159
rect 37277 36119 37335 36125
rect 37544 36159 37602 36165
rect 37544 36125 37556 36159
rect 37590 36156 37602 36159
rect 38746 36156 38752 36168
rect 37590 36128 38752 36156
rect 37590 36125 37602 36128
rect 37544 36119 37602 36125
rect 38746 36116 38752 36128
rect 38804 36116 38810 36168
rect 39942 36116 39948 36168
rect 40000 36116 40006 36168
rect 40120 36159 40178 36165
rect 40120 36125 40132 36159
rect 40166 36156 40178 36159
rect 40494 36156 40500 36168
rect 40166 36128 40500 36156
rect 40166 36125 40178 36128
rect 40120 36119 40178 36125
rect 40494 36116 40500 36128
rect 40552 36116 40558 36168
rect 41693 36159 41751 36165
rect 41693 36156 41705 36159
rect 40880 36128 41705 36156
rect 29816 36091 29874 36097
rect 29816 36057 29828 36091
rect 29862 36088 29874 36091
rect 31018 36088 31024 36100
rect 29862 36060 31024 36088
rect 29862 36057 29874 36060
rect 29816 36051 29874 36057
rect 31018 36048 31024 36060
rect 31076 36048 31082 36100
rect 32306 36088 32312 36100
rect 32219 36060 32312 36088
rect 32306 36048 32312 36060
rect 32364 36048 32370 36100
rect 35152 36091 35210 36097
rect 35152 36057 35164 36091
rect 35198 36088 35210 36091
rect 36078 36088 36084 36100
rect 35198 36060 36084 36088
rect 35198 36057 35210 36060
rect 35152 36051 35210 36057
rect 36078 36048 36084 36060
rect 36136 36048 36142 36100
rect 39960 36088 39988 36116
rect 40880 36088 40908 36128
rect 41693 36125 41705 36128
rect 41739 36156 41751 36159
rect 42426 36156 42432 36168
rect 41739 36128 42432 36156
rect 41739 36125 41751 36128
rect 41693 36119 41751 36125
rect 42426 36116 42432 36128
rect 42484 36116 42490 36168
rect 50154 36116 50160 36168
rect 50212 36165 50218 36168
rect 50212 36156 50222 36165
rect 51997 36159 52055 36165
rect 50212 36128 50257 36156
rect 50212 36119 50222 36128
rect 51997 36125 52009 36159
rect 52043 36156 52055 36159
rect 52730 36156 52736 36168
rect 52043 36128 52736 36156
rect 52043 36125 52055 36128
rect 51997 36119 52055 36125
rect 50212 36116 50218 36119
rect 52730 36116 52736 36128
rect 52788 36116 52794 36168
rect 55306 36156 55312 36168
rect 55267 36128 55312 36156
rect 55306 36116 55312 36128
rect 55364 36116 55370 36168
rect 41938 36091 41996 36097
rect 41938 36088 41950 36091
rect 39960 36060 40908 36088
rect 41248 36060 41950 36088
rect 29914 36020 29920 36032
rect 29564 35992 29920 36020
rect 25823 35989 25835 35992
rect 25777 35983 25835 35989
rect 29914 35980 29920 35992
rect 29972 35980 29978 36032
rect 32324 36020 32352 36048
rect 35986 36020 35992 36032
rect 32324 35992 35992 36020
rect 35986 35980 35992 35992
rect 36044 35980 36050 36032
rect 36265 36023 36323 36029
rect 36265 35989 36277 36023
rect 36311 36020 36323 36023
rect 37366 36020 37372 36032
rect 36311 35992 37372 36020
rect 36311 35989 36323 35992
rect 36265 35983 36323 35989
rect 37366 35980 37372 35992
rect 37424 35980 37430 36032
rect 41248 36029 41276 36060
rect 41938 36057 41950 36060
rect 41984 36057 41996 36091
rect 41938 36051 41996 36057
rect 46477 36091 46535 36097
rect 46477 36057 46489 36091
rect 46523 36088 46535 36091
rect 49786 36088 49792 36100
rect 46523 36060 49792 36088
rect 46523 36057 46535 36060
rect 46477 36051 46535 36057
rect 49786 36048 49792 36060
rect 49844 36048 49850 36100
rect 50062 36048 50068 36100
rect 50120 36088 50126 36100
rect 50402 36091 50460 36097
rect 50402 36088 50414 36091
rect 50120 36060 50414 36088
rect 50120 36048 50126 36060
rect 50402 36057 50414 36060
rect 50448 36057 50460 36091
rect 50402 36051 50460 36057
rect 51258 36048 51264 36100
rect 51316 36088 51322 36100
rect 52242 36091 52300 36097
rect 52242 36088 52254 36091
rect 51316 36060 52254 36088
rect 51316 36048 51322 36060
rect 52242 36057 52254 36060
rect 52288 36057 52300 36091
rect 52242 36051 52300 36057
rect 55576 36091 55634 36097
rect 55576 36057 55588 36091
rect 55622 36088 55634 36091
rect 56594 36088 56600 36100
rect 55622 36060 56600 36088
rect 55622 36057 55634 36060
rect 55576 36051 55634 36057
rect 56594 36048 56600 36060
rect 56652 36048 56658 36100
rect 41233 36023 41291 36029
rect 41233 35989 41245 36023
rect 41279 35989 41291 36023
rect 41233 35983 41291 35989
rect 41414 35980 41420 36032
rect 41472 36020 41478 36032
rect 43073 36023 43131 36029
rect 43073 36020 43085 36023
rect 41472 35992 43085 36020
rect 41472 35980 41478 35992
rect 43073 35989 43085 35992
rect 43119 35989 43131 36023
rect 43073 35983 43131 35989
rect 52546 35980 52552 36032
rect 52604 36020 52610 36032
rect 53377 36023 53435 36029
rect 53377 36020 53389 36023
rect 52604 35992 53389 36020
rect 52604 35980 52610 35992
rect 53377 35989 53389 35992
rect 53423 35989 53435 36023
rect 53377 35983 53435 35989
rect 1104 35930 59340 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 59340 35930
rect 1104 35856 59340 35878
rect 6730 35776 6736 35828
rect 6788 35816 6794 35828
rect 7745 35819 7803 35825
rect 7745 35816 7757 35819
rect 6788 35788 7757 35816
rect 6788 35776 6794 35788
rect 7745 35785 7757 35788
rect 7791 35785 7803 35819
rect 7745 35779 7803 35785
rect 23201 35819 23259 35825
rect 23201 35785 23213 35819
rect 23247 35785 23259 35819
rect 23201 35779 23259 35785
rect 6632 35751 6690 35757
rect 6632 35717 6644 35751
rect 6678 35748 6690 35751
rect 7926 35748 7932 35760
rect 6678 35720 7932 35748
rect 6678 35717 6690 35720
rect 6632 35711 6690 35717
rect 7926 35708 7932 35720
rect 7984 35708 7990 35760
rect 11784 35751 11842 35757
rect 11784 35717 11796 35751
rect 11830 35748 11842 35751
rect 12894 35748 12900 35760
rect 11830 35720 12900 35748
rect 11830 35717 11842 35720
rect 11784 35711 11842 35717
rect 12894 35708 12900 35720
rect 12952 35708 12958 35760
rect 13998 35748 14004 35760
rect 13372 35720 14004 35748
rect 3970 35680 3976 35692
rect 3931 35652 3976 35680
rect 3970 35640 3976 35652
rect 4028 35640 4034 35692
rect 11514 35680 11520 35692
rect 11427 35652 11520 35680
rect 11514 35640 11520 35652
rect 11572 35680 11578 35692
rect 11572 35652 12572 35680
rect 11572 35640 11578 35652
rect 6362 35612 6368 35624
rect 6323 35584 6368 35612
rect 6362 35572 6368 35584
rect 6420 35572 6426 35624
rect 12544 35612 12572 35652
rect 13372 35621 13400 35720
rect 13998 35708 14004 35720
rect 14056 35708 14062 35760
rect 22094 35757 22100 35760
rect 22088 35748 22100 35757
rect 22055 35720 22100 35748
rect 22088 35711 22100 35720
rect 22094 35708 22100 35711
rect 22152 35708 22158 35760
rect 23216 35748 23244 35779
rect 23658 35776 23664 35828
rect 23716 35816 23722 35828
rect 24394 35816 24400 35828
rect 23716 35788 24400 35816
rect 23716 35776 23722 35788
rect 24394 35776 24400 35788
rect 24452 35776 24458 35828
rect 25038 35816 25044 35828
rect 24999 35788 25044 35816
rect 25038 35776 25044 35788
rect 25096 35776 25102 35828
rect 28902 35776 28908 35828
rect 28960 35816 28966 35828
rect 29546 35816 29552 35828
rect 28960 35788 29552 35816
rect 28960 35776 28966 35788
rect 29546 35776 29552 35788
rect 29604 35776 29610 35828
rect 29914 35776 29920 35828
rect 29972 35816 29978 35828
rect 31754 35816 31760 35828
rect 29972 35788 31760 35816
rect 29972 35776 29978 35788
rect 31754 35776 31760 35788
rect 31812 35776 31818 35828
rect 33502 35816 33508 35828
rect 33463 35788 33508 35816
rect 33502 35776 33508 35788
rect 33560 35776 33566 35828
rect 36078 35816 36084 35828
rect 36039 35788 36084 35816
rect 36078 35776 36084 35788
rect 36136 35776 36142 35828
rect 39390 35816 39396 35828
rect 39351 35788 39396 35816
rect 39390 35776 39396 35788
rect 39448 35776 39454 35828
rect 41325 35819 41383 35825
rect 41325 35785 41337 35819
rect 41371 35816 41383 35819
rect 41371 35788 42012 35816
rect 41371 35785 41383 35788
rect 41325 35779 41383 35785
rect 23906 35751 23964 35757
rect 23906 35748 23918 35751
rect 23216 35720 23918 35748
rect 23906 35717 23918 35720
rect 23952 35717 23964 35751
rect 23906 35711 23964 35717
rect 13446 35640 13452 35692
rect 13504 35680 13510 35692
rect 13613 35683 13671 35689
rect 13613 35680 13625 35683
rect 13504 35652 13625 35680
rect 13504 35640 13510 35652
rect 13613 35649 13625 35652
rect 13659 35649 13671 35683
rect 13613 35643 13671 35649
rect 18233 35683 18291 35689
rect 18233 35649 18245 35683
rect 18279 35680 18291 35683
rect 20714 35680 20720 35692
rect 18279 35652 20720 35680
rect 18279 35649 18291 35652
rect 18233 35643 18291 35649
rect 20714 35640 20720 35652
rect 20772 35640 20778 35692
rect 21082 35640 21088 35692
rect 21140 35680 21146 35692
rect 21821 35683 21879 35689
rect 21821 35680 21833 35683
rect 21140 35652 21833 35680
rect 21140 35640 21146 35652
rect 21821 35649 21833 35652
rect 21867 35680 21879 35683
rect 23658 35680 23664 35692
rect 21867 35652 23664 35680
rect 21867 35649 21879 35652
rect 21821 35643 21879 35649
rect 23658 35640 23664 35652
rect 23716 35640 23722 35692
rect 27332 35683 27390 35689
rect 27332 35649 27344 35683
rect 27378 35680 27390 35683
rect 28350 35680 28356 35692
rect 27378 35652 28356 35680
rect 27378 35649 27390 35652
rect 27332 35643 27390 35649
rect 28350 35640 28356 35652
rect 28408 35640 28414 35692
rect 29172 35683 29230 35689
rect 29172 35649 29184 35683
rect 29218 35680 29230 35683
rect 30190 35680 30196 35692
rect 29218 35652 30196 35680
rect 29218 35649 29230 35652
rect 29172 35643 29230 35649
rect 30190 35640 30196 35652
rect 30248 35640 30254 35692
rect 31772 35680 31800 35776
rect 32392 35751 32450 35757
rect 32392 35717 32404 35751
rect 32438 35748 32450 35751
rect 36722 35748 36728 35760
rect 32438 35720 36728 35748
rect 32438 35717 32450 35720
rect 32392 35711 32450 35717
rect 36722 35708 36728 35720
rect 36780 35708 36786 35760
rect 38280 35751 38338 35757
rect 38280 35717 38292 35751
rect 38326 35748 38338 35751
rect 39482 35748 39488 35760
rect 38326 35720 39488 35748
rect 38326 35717 38338 35720
rect 38280 35711 38338 35717
rect 39482 35708 39488 35720
rect 39540 35708 39546 35760
rect 40212 35751 40270 35757
rect 40212 35717 40224 35751
rect 40258 35748 40270 35751
rect 41414 35748 41420 35760
rect 40258 35720 41420 35748
rect 40258 35717 40270 35720
rect 40212 35711 40270 35717
rect 41414 35708 41420 35720
rect 41472 35708 41478 35760
rect 41984 35748 42012 35788
rect 42674 35751 42732 35757
rect 42674 35748 42686 35751
rect 41984 35720 42686 35748
rect 42674 35717 42686 35720
rect 42720 35717 42732 35751
rect 42674 35711 42732 35717
rect 45916 35751 45974 35757
rect 45916 35717 45928 35751
rect 45962 35748 45974 35751
rect 47026 35748 47032 35760
rect 45962 35720 47032 35748
rect 45962 35717 45974 35720
rect 45916 35711 45974 35717
rect 47026 35708 47032 35720
rect 47084 35708 47090 35760
rect 55306 35748 55312 35760
rect 54588 35720 55312 35748
rect 32125 35683 32183 35689
rect 32125 35680 32137 35683
rect 31772 35652 32137 35680
rect 32125 35649 32137 35652
rect 32171 35649 32183 35683
rect 32125 35643 32183 35649
rect 34968 35683 35026 35689
rect 34968 35649 34980 35683
rect 35014 35680 35026 35683
rect 36354 35680 36360 35692
rect 35014 35652 36360 35680
rect 35014 35649 35026 35652
rect 34968 35643 35026 35649
rect 36354 35640 36360 35652
rect 36412 35640 36418 35692
rect 42429 35683 42487 35689
rect 42429 35649 42441 35683
rect 42475 35680 42487 35683
rect 42518 35680 42524 35692
rect 42475 35652 42524 35680
rect 42475 35649 42487 35652
rect 42429 35643 42487 35649
rect 42518 35640 42524 35652
rect 42576 35640 42582 35692
rect 49320 35683 49378 35689
rect 49320 35649 49332 35683
rect 49366 35680 49378 35683
rect 50798 35680 50804 35692
rect 49366 35652 50804 35680
rect 49366 35649 49378 35652
rect 49320 35643 49378 35649
rect 50798 35640 50804 35652
rect 50856 35640 50862 35692
rect 53000 35683 53058 35689
rect 53000 35649 53012 35683
rect 53046 35680 53058 35683
rect 53926 35680 53932 35692
rect 53046 35652 53932 35680
rect 53046 35649 53058 35652
rect 53000 35643 53058 35649
rect 53926 35640 53932 35652
rect 53984 35640 53990 35692
rect 54588 35689 54616 35720
rect 55306 35708 55312 35720
rect 55364 35708 55370 35760
rect 54573 35683 54631 35689
rect 54573 35649 54585 35683
rect 54619 35649 54631 35683
rect 54573 35643 54631 35649
rect 54840 35683 54898 35689
rect 54840 35649 54852 35683
rect 54886 35680 54898 35683
rect 56778 35680 56784 35692
rect 54886 35652 56784 35680
rect 54886 35649 54898 35652
rect 54840 35643 54898 35649
rect 56778 35640 56784 35652
rect 56836 35640 56842 35692
rect 13357 35615 13415 35621
rect 13357 35612 13369 35615
rect 12544 35584 13369 35612
rect 13357 35581 13369 35584
rect 13403 35581 13415 35615
rect 27062 35612 27068 35624
rect 27023 35584 27068 35612
rect 13357 35575 13415 35581
rect 27062 35572 27068 35584
rect 27120 35572 27126 35624
rect 28902 35612 28908 35624
rect 28276 35584 28908 35612
rect 4982 35436 4988 35488
rect 5040 35476 5046 35488
rect 5261 35479 5319 35485
rect 5261 35476 5273 35479
rect 5040 35448 5273 35476
rect 5040 35436 5046 35448
rect 5261 35445 5273 35448
rect 5307 35445 5319 35479
rect 12894 35476 12900 35488
rect 12855 35448 12900 35476
rect 5261 35439 5319 35445
rect 12894 35436 12900 35448
rect 12952 35436 12958 35488
rect 13630 35436 13636 35488
rect 13688 35476 13694 35488
rect 14737 35479 14795 35485
rect 14737 35476 14749 35479
rect 13688 35448 14749 35476
rect 13688 35436 13694 35448
rect 14737 35445 14749 35448
rect 14783 35445 14795 35479
rect 14737 35439 14795 35445
rect 16666 35436 16672 35488
rect 16724 35476 16730 35488
rect 17862 35476 17868 35488
rect 16724 35448 17868 35476
rect 16724 35436 16730 35448
rect 17862 35436 17868 35448
rect 17920 35476 17926 35488
rect 19242 35476 19248 35488
rect 17920 35448 19248 35476
rect 17920 35436 17926 35448
rect 19242 35436 19248 35448
rect 19300 35476 19306 35488
rect 19521 35479 19579 35485
rect 19521 35476 19533 35479
rect 19300 35448 19533 35476
rect 19300 35436 19306 35448
rect 19521 35445 19533 35448
rect 19567 35445 19579 35479
rect 19521 35439 19579 35445
rect 27062 35436 27068 35488
rect 27120 35476 27126 35488
rect 28276 35476 28304 35584
rect 28902 35572 28908 35584
rect 28960 35572 28966 35624
rect 34606 35572 34612 35624
rect 34664 35612 34670 35624
rect 34701 35615 34759 35621
rect 34701 35612 34713 35615
rect 34664 35584 34713 35612
rect 34664 35572 34670 35584
rect 34701 35581 34713 35584
rect 34747 35581 34759 35615
rect 34701 35575 34759 35581
rect 37734 35572 37740 35624
rect 37792 35612 37798 35624
rect 38013 35615 38071 35621
rect 38013 35612 38025 35615
rect 37792 35584 38025 35612
rect 37792 35572 37798 35584
rect 38013 35581 38025 35584
rect 38059 35581 38071 35615
rect 38013 35575 38071 35581
rect 39850 35572 39856 35624
rect 39908 35612 39914 35624
rect 39945 35615 40003 35621
rect 39945 35612 39957 35615
rect 39908 35584 39957 35612
rect 39908 35572 39914 35584
rect 39945 35581 39957 35584
rect 39991 35581 40003 35615
rect 39945 35575 40003 35581
rect 45554 35572 45560 35624
rect 45612 35612 45618 35624
rect 45649 35615 45707 35621
rect 45649 35612 45661 35615
rect 45612 35584 45661 35612
rect 45612 35572 45618 35584
rect 45649 35581 45661 35584
rect 45695 35581 45707 35615
rect 45649 35575 45707 35581
rect 49053 35615 49111 35621
rect 49053 35581 49065 35615
rect 49099 35581 49111 35615
rect 52730 35612 52736 35624
rect 52691 35584 52736 35612
rect 49053 35575 49111 35581
rect 28442 35476 28448 35488
rect 27120 35448 28304 35476
rect 28403 35448 28448 35476
rect 27120 35436 27126 35448
rect 28442 35436 28448 35448
rect 28500 35436 28506 35488
rect 30282 35476 30288 35488
rect 30243 35448 30288 35476
rect 30282 35436 30288 35448
rect 30340 35436 30346 35488
rect 40678 35436 40684 35488
rect 40736 35476 40742 35488
rect 43809 35479 43867 35485
rect 43809 35476 43821 35479
rect 40736 35448 43821 35476
rect 40736 35436 40742 35448
rect 43809 35445 43821 35448
rect 43855 35445 43867 35479
rect 47026 35476 47032 35488
rect 46987 35448 47032 35476
rect 43809 35439 43867 35445
rect 47026 35436 47032 35448
rect 47084 35436 47090 35488
rect 49068 35476 49096 35575
rect 52730 35572 52736 35584
rect 52788 35572 52794 35624
rect 50154 35476 50160 35488
rect 49068 35448 50160 35476
rect 50154 35436 50160 35448
rect 50212 35436 50218 35488
rect 50433 35479 50491 35485
rect 50433 35445 50445 35479
rect 50479 35476 50491 35479
rect 51166 35476 51172 35488
rect 50479 35448 51172 35476
rect 50479 35445 50491 35448
rect 50433 35439 50491 35445
rect 51166 35436 51172 35448
rect 51224 35436 51230 35488
rect 54110 35476 54116 35488
rect 54071 35448 54116 35476
rect 54110 35436 54116 35448
rect 54168 35436 54174 35488
rect 55950 35476 55956 35488
rect 55911 35448 55956 35476
rect 55950 35436 55956 35448
rect 56008 35436 56014 35488
rect 1104 35386 59340 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 59340 35386
rect 1104 35312 59340 35334
rect 12897 35275 12955 35281
rect 12897 35241 12909 35275
rect 12943 35272 12955 35275
rect 13814 35272 13820 35284
rect 12943 35244 13820 35272
rect 12943 35241 12955 35244
rect 12897 35235 12955 35241
rect 13814 35232 13820 35244
rect 13872 35232 13878 35284
rect 16666 35272 16672 35284
rect 16408 35244 16672 35272
rect 6822 35096 6828 35148
rect 6880 35136 6886 35148
rect 6917 35139 6975 35145
rect 6917 35136 6929 35139
rect 6880 35108 6929 35136
rect 6880 35096 6886 35108
rect 6917 35105 6929 35108
rect 6963 35105 6975 35139
rect 11514 35136 11520 35148
rect 11475 35108 11520 35136
rect 6917 35099 6975 35105
rect 11514 35096 11520 35108
rect 11572 35096 11578 35148
rect 16408 35145 16436 35244
rect 16666 35232 16672 35244
rect 16724 35232 16730 35284
rect 17770 35272 17776 35284
rect 17731 35244 17776 35272
rect 17770 35232 17776 35244
rect 17828 35232 17834 35284
rect 28350 35232 28356 35284
rect 28408 35272 28414 35284
rect 28445 35275 28503 35281
rect 28445 35272 28457 35275
rect 28408 35244 28457 35272
rect 28408 35232 28414 35244
rect 28445 35241 28457 35244
rect 28491 35241 28503 35275
rect 31018 35272 31024 35284
rect 30979 35244 31024 35272
rect 28445 35235 28503 35241
rect 31018 35232 31024 35244
rect 31076 35232 31082 35284
rect 31754 35272 31760 35284
rect 31496 35244 31760 35272
rect 16393 35139 16451 35145
rect 16393 35105 16405 35139
rect 16439 35105 16451 35139
rect 19242 35136 19248 35148
rect 19203 35108 19248 35136
rect 16393 35099 16451 35105
rect 19242 35096 19248 35108
rect 19300 35096 19306 35148
rect 21082 35136 21088 35148
rect 21043 35108 21088 35136
rect 21082 35096 21088 35108
rect 21140 35096 21146 35148
rect 28902 35096 28908 35148
rect 28960 35136 28966 35148
rect 31496 35145 31524 35244
rect 31754 35232 31760 35244
rect 31812 35232 31818 35284
rect 44450 35272 44456 35284
rect 44411 35244 44456 35272
rect 44450 35232 44456 35244
rect 44508 35232 44514 35284
rect 45554 35232 45560 35284
rect 45612 35272 45618 35284
rect 47029 35275 47087 35281
rect 45612 35244 46612 35272
rect 45612 35232 45618 35244
rect 29641 35139 29699 35145
rect 29641 35136 29653 35139
rect 28960 35108 29653 35136
rect 28960 35096 28966 35108
rect 29641 35105 29653 35108
rect 29687 35105 29699 35139
rect 29641 35099 29699 35105
rect 31481 35139 31539 35145
rect 31481 35105 31493 35139
rect 31527 35105 31539 35139
rect 37734 35136 37740 35148
rect 37695 35108 37740 35136
rect 31481 35099 31539 35105
rect 37734 35096 37740 35108
rect 37792 35096 37798 35148
rect 39942 35096 39948 35148
rect 40000 35136 40006 35148
rect 45664 35145 45692 35244
rect 46584 35204 46612 35244
rect 47029 35241 47041 35275
rect 47075 35272 47087 35275
rect 47118 35272 47124 35284
rect 47075 35244 47124 35272
rect 47075 35241 47087 35244
rect 47029 35235 47087 35241
rect 47118 35232 47124 35244
rect 47176 35232 47182 35284
rect 46842 35204 46848 35216
rect 46584 35176 46848 35204
rect 46842 35164 46848 35176
rect 46900 35204 46906 35216
rect 46900 35176 47716 35204
rect 46900 35164 46906 35176
rect 47688 35145 47716 35176
rect 40405 35139 40463 35145
rect 40405 35136 40417 35139
rect 40000 35108 40417 35136
rect 40000 35096 40006 35108
rect 40405 35105 40417 35108
rect 40451 35105 40463 35139
rect 45649 35139 45707 35145
rect 45649 35136 45661 35139
rect 40405 35099 40463 35105
rect 45526 35108 45661 35136
rect 11784 35071 11842 35077
rect 11784 35037 11796 35071
rect 11830 35068 11842 35071
rect 12894 35068 12900 35080
rect 11830 35040 12900 35068
rect 11830 35037 11842 35040
rect 11784 35031 11842 35037
rect 12894 35028 12900 35040
rect 12952 35028 12958 35080
rect 13998 35028 14004 35080
rect 14056 35068 14062 35080
rect 19518 35077 19524 35080
rect 14093 35071 14151 35077
rect 14093 35068 14105 35071
rect 14056 35040 14105 35068
rect 14056 35028 14062 35040
rect 14093 35037 14105 35040
rect 14139 35037 14151 35071
rect 14093 35031 14151 35037
rect 19512 35031 19524 35077
rect 19576 35068 19582 35080
rect 19576 35040 19612 35068
rect 19518 35028 19524 35031
rect 19576 35028 19582 35040
rect 24394 35028 24400 35080
rect 24452 35068 24458 35080
rect 25225 35071 25283 35077
rect 25225 35068 25237 35071
rect 24452 35040 25237 35068
rect 24452 35028 24458 35040
rect 25225 35037 25237 35040
rect 25271 35037 25283 35071
rect 25225 35031 25283 35037
rect 26234 35028 26240 35080
rect 26292 35068 26298 35080
rect 27062 35068 27068 35080
rect 26292 35040 27068 35068
rect 26292 35028 26298 35040
rect 27062 35028 27068 35040
rect 27120 35028 27126 35080
rect 29908 35071 29966 35077
rect 29908 35037 29920 35071
rect 29954 35068 29966 35071
rect 30282 35068 30288 35080
rect 29954 35040 30288 35068
rect 29954 35037 29966 35040
rect 29908 35031 29966 35037
rect 30282 35028 30288 35040
rect 30340 35028 30346 35080
rect 40678 35077 40684 35080
rect 40672 35068 40684 35077
rect 40639 35040 40684 35068
rect 40672 35031 40684 35040
rect 40678 35028 40684 35031
rect 40736 35028 40742 35080
rect 43073 35071 43131 35077
rect 43073 35037 43085 35071
rect 43119 35068 43131 35071
rect 44174 35068 44180 35080
rect 43119 35040 44180 35068
rect 43119 35037 43131 35040
rect 43073 35031 43131 35037
rect 44174 35028 44180 35040
rect 44232 35068 44238 35080
rect 45526 35068 45554 35108
rect 45649 35105 45661 35108
rect 45695 35105 45707 35139
rect 45649 35099 45707 35105
rect 47673 35139 47731 35145
rect 47673 35105 47685 35139
rect 47719 35105 47731 35139
rect 55306 35136 55312 35148
rect 55267 35108 55312 35136
rect 47673 35099 47731 35105
rect 55306 35096 55312 35108
rect 55364 35096 55370 35148
rect 44232 35040 45554 35068
rect 45916 35071 45974 35077
rect 44232 35028 44238 35040
rect 45916 35037 45928 35071
rect 45962 35068 45974 35071
rect 47026 35068 47032 35080
rect 45962 35040 47032 35068
rect 45962 35037 45974 35040
rect 45916 35031 45974 35037
rect 47026 35028 47032 35040
rect 47084 35028 47090 35080
rect 50154 35068 50160 35080
rect 50115 35040 50160 35068
rect 50154 35028 50160 35040
rect 50212 35068 50218 35080
rect 51997 35071 52055 35077
rect 51997 35068 52009 35071
rect 50212 35040 52009 35068
rect 50212 35028 50218 35040
rect 51997 35037 52009 35040
rect 52043 35037 52055 35071
rect 51997 35031 52055 35037
rect 55576 35071 55634 35077
rect 55576 35037 55588 35071
rect 55622 35068 55634 35071
rect 55950 35068 55956 35080
rect 55622 35040 55956 35068
rect 55622 35037 55634 35040
rect 55576 35031 55634 35037
rect 55950 35028 55956 35040
rect 56008 35028 56014 35080
rect 57146 35068 57152 35080
rect 57107 35040 57152 35068
rect 57146 35028 57152 35040
rect 57204 35028 57210 35080
rect 7184 35003 7242 35009
rect 7184 34969 7196 35003
rect 7230 35000 7242 35003
rect 9582 35000 9588 35012
rect 7230 34972 9588 35000
rect 7230 34969 7242 34972
rect 7184 34963 7242 34969
rect 9582 34960 9588 34972
rect 9640 34960 9646 35012
rect 14360 35003 14418 35009
rect 14360 34969 14372 35003
rect 14406 35000 14418 35003
rect 14734 35000 14740 35012
rect 14406 34972 14740 35000
rect 14406 34969 14418 34972
rect 14360 34963 14418 34969
rect 14734 34960 14740 34972
rect 14792 34960 14798 35012
rect 16660 35003 16718 35009
rect 16660 34969 16672 35003
rect 16706 35000 16718 35003
rect 18230 35000 18236 35012
rect 16706 34972 18236 35000
rect 16706 34969 16718 34972
rect 16660 34963 16718 34969
rect 18230 34960 18236 34972
rect 18288 34960 18294 35012
rect 21352 35003 21410 35009
rect 21352 34969 21364 35003
rect 21398 35000 21410 35003
rect 22830 35000 22836 35012
rect 21398 34972 22836 35000
rect 21398 34969 21410 34972
rect 21352 34963 21410 34969
rect 22830 34960 22836 34972
rect 22888 34960 22894 35012
rect 25492 35003 25550 35009
rect 25492 34969 25504 35003
rect 25538 35000 25550 35003
rect 26970 35000 26976 35012
rect 25538 34972 26976 35000
rect 25538 34969 25550 34972
rect 25492 34963 25550 34969
rect 26970 34960 26976 34972
rect 27028 34960 27034 35012
rect 27332 35003 27390 35009
rect 27332 34969 27344 35003
rect 27378 35000 27390 35003
rect 28350 35000 28356 35012
rect 27378 34972 28356 35000
rect 27378 34969 27390 34972
rect 27332 34963 27390 34969
rect 28350 34960 28356 34972
rect 28408 34960 28414 35012
rect 31748 35003 31806 35009
rect 31748 34969 31760 35003
rect 31794 35000 31806 35003
rect 31846 35000 31852 35012
rect 31794 34972 31852 35000
rect 31794 34969 31806 34972
rect 31748 34963 31806 34969
rect 31846 34960 31852 34972
rect 31904 34960 31910 35012
rect 35986 35000 35992 35012
rect 35899 34972 35992 35000
rect 35986 34960 35992 34972
rect 36044 35000 36050 35012
rect 40126 35000 40132 35012
rect 36044 34972 40132 35000
rect 36044 34960 36050 34972
rect 40126 34960 40132 34972
rect 40184 34960 40190 35012
rect 43340 35003 43398 35009
rect 43340 34969 43352 35003
rect 43386 35000 43398 35003
rect 46842 35000 46848 35012
rect 43386 34972 46848 35000
rect 43386 34969 43398 34972
rect 43340 34963 43398 34969
rect 46842 34960 46848 34972
rect 46900 34960 46906 35012
rect 47940 35003 47998 35009
rect 47940 34969 47952 35003
rect 47986 35000 47998 35003
rect 48958 35000 48964 35012
rect 47986 34972 48964 35000
rect 47986 34969 47998 34972
rect 47940 34963 47998 34969
rect 48958 34960 48964 34972
rect 49016 34960 49022 35012
rect 50424 35003 50482 35009
rect 50424 34969 50436 35003
rect 50470 35000 50482 35003
rect 51902 35000 51908 35012
rect 50470 34972 51908 35000
rect 50470 34969 50482 34972
rect 50424 34963 50482 34969
rect 51902 34960 51908 34972
rect 51960 34960 51966 35012
rect 52264 35003 52322 35009
rect 52264 34969 52276 35003
rect 52310 35000 52322 35003
rect 54018 35000 54024 35012
rect 52310 34972 54024 35000
rect 52310 34969 52322 34972
rect 52264 34963 52322 34969
rect 54018 34960 54024 34972
rect 54076 34960 54082 35012
rect 56870 34960 56876 35012
rect 56928 35000 56934 35012
rect 57394 35003 57452 35009
rect 57394 35000 57406 35003
rect 56928 34972 57406 35000
rect 56928 34960 56934 34972
rect 57394 34969 57406 34972
rect 57440 34969 57452 35003
rect 57394 34963 57452 34969
rect 8294 34932 8300 34944
rect 8255 34904 8300 34932
rect 8294 34892 8300 34904
rect 8352 34892 8358 34944
rect 15470 34932 15476 34944
rect 15431 34904 15476 34932
rect 15470 34892 15476 34904
rect 15528 34892 15534 34944
rect 20622 34932 20628 34944
rect 20583 34904 20628 34932
rect 20622 34892 20628 34904
rect 20680 34892 20686 34944
rect 22462 34932 22468 34944
rect 22423 34904 22468 34932
rect 22462 34892 22468 34904
rect 22520 34892 22526 34944
rect 26602 34932 26608 34944
rect 26563 34904 26608 34932
rect 26602 34892 26608 34904
rect 26660 34892 26666 34944
rect 30374 34892 30380 34944
rect 30432 34932 30438 34944
rect 32861 34935 32919 34941
rect 32861 34932 32873 34935
rect 30432 34904 32873 34932
rect 30432 34892 30438 34904
rect 32861 34901 32873 34904
rect 32907 34901 32919 34935
rect 41782 34932 41788 34944
rect 41743 34904 41788 34932
rect 32861 34895 32919 34901
rect 41782 34892 41788 34904
rect 41840 34892 41846 34944
rect 49053 34935 49111 34941
rect 49053 34901 49065 34935
rect 49099 34932 49111 34935
rect 49694 34932 49700 34944
rect 49099 34904 49700 34932
rect 49099 34901 49111 34904
rect 49053 34895 49111 34901
rect 49694 34892 49700 34904
rect 49752 34892 49758 34944
rect 51537 34935 51595 34941
rect 51537 34901 51549 34935
rect 51583 34932 51595 34935
rect 52086 34932 52092 34944
rect 51583 34904 52092 34932
rect 51583 34901 51595 34904
rect 51537 34895 51595 34901
rect 52086 34892 52092 34904
rect 52144 34892 52150 34944
rect 53006 34892 53012 34944
rect 53064 34932 53070 34944
rect 53377 34935 53435 34941
rect 53377 34932 53389 34935
rect 53064 34904 53389 34932
rect 53064 34892 53070 34904
rect 53377 34901 53389 34904
rect 53423 34901 53435 34935
rect 56686 34932 56692 34944
rect 56647 34904 56692 34932
rect 53377 34895 53435 34901
rect 56686 34892 56692 34904
rect 56744 34892 56750 34944
rect 58529 34935 58587 34941
rect 58529 34901 58541 34935
rect 58575 34932 58587 34935
rect 59449 34935 59507 34941
rect 59449 34932 59461 34935
rect 58575 34904 59461 34932
rect 58575 34901 58587 34904
rect 58529 34895 58587 34901
rect 59449 34901 59461 34904
rect 59495 34901 59507 34935
rect 59449 34895 59507 34901
rect 1104 34842 59340 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 59340 34842
rect 1104 34768 59340 34790
rect 10321 34731 10379 34737
rect 10321 34697 10333 34731
rect 10367 34728 10379 34731
rect 11054 34728 11060 34740
rect 10367 34700 11060 34728
rect 10367 34697 10379 34700
rect 10321 34691 10379 34697
rect 11054 34688 11060 34700
rect 11112 34688 11118 34740
rect 12897 34731 12955 34737
rect 12897 34697 12909 34731
rect 12943 34728 12955 34731
rect 13446 34728 13452 34740
rect 12943 34700 13452 34728
rect 12943 34697 12955 34700
rect 12897 34691 12955 34697
rect 13446 34688 13452 34700
rect 13504 34688 13510 34740
rect 14734 34728 14740 34740
rect 14695 34700 14740 34728
rect 14734 34688 14740 34700
rect 14792 34688 14798 34740
rect 18230 34728 18236 34740
rect 18191 34700 18236 34728
rect 18230 34688 18236 34700
rect 18288 34688 18294 34740
rect 23201 34731 23259 34737
rect 23201 34697 23213 34731
rect 23247 34728 23259 34731
rect 24486 34728 24492 34740
rect 23247 34700 24492 34728
rect 23247 34697 23259 34700
rect 23201 34691 23259 34697
rect 24486 34688 24492 34700
rect 24544 34688 24550 34740
rect 24670 34688 24676 34740
rect 24728 34728 24734 34740
rect 25133 34731 25191 34737
rect 25133 34728 25145 34731
rect 24728 34700 25145 34728
rect 24728 34688 24734 34700
rect 25133 34697 25145 34700
rect 25179 34697 25191 34731
rect 28350 34728 28356 34740
rect 28311 34700 28356 34728
rect 25133 34691 25191 34697
rect 28350 34688 28356 34700
rect 28408 34688 28414 34740
rect 30190 34728 30196 34740
rect 30151 34700 30196 34728
rect 30190 34688 30196 34700
rect 30248 34688 30254 34740
rect 36354 34728 36360 34740
rect 36315 34700 36360 34728
rect 36354 34688 36360 34700
rect 36412 34688 36418 34740
rect 38657 34731 38715 34737
rect 38657 34697 38669 34731
rect 38703 34728 38715 34731
rect 38838 34728 38844 34740
rect 38703 34700 38844 34728
rect 38703 34697 38715 34700
rect 38657 34691 38715 34697
rect 38838 34688 38844 34700
rect 38896 34688 38902 34740
rect 39114 34688 39120 34740
rect 39172 34728 39178 34740
rect 40497 34731 40555 34737
rect 40497 34728 40509 34731
rect 39172 34700 40509 34728
rect 39172 34688 39178 34700
rect 40497 34697 40509 34700
rect 40543 34697 40555 34731
rect 40497 34691 40555 34697
rect 45646 34688 45652 34740
rect 45704 34728 45710 34740
rect 46842 34728 46848 34740
rect 45704 34700 45784 34728
rect 46803 34700 46848 34728
rect 45704 34688 45710 34700
rect 3970 34620 3976 34672
rect 4028 34660 4034 34672
rect 6733 34663 6791 34669
rect 6733 34660 6745 34663
rect 4028 34632 6745 34660
rect 4028 34620 4034 34632
rect 6733 34629 6745 34632
rect 6779 34660 6791 34663
rect 11882 34660 11888 34672
rect 6779 34632 11888 34660
rect 6779 34629 6791 34632
rect 6733 34623 6791 34629
rect 11882 34620 11888 34632
rect 11940 34620 11946 34672
rect 13630 34669 13636 34672
rect 13624 34660 13636 34669
rect 13591 34632 13636 34660
rect 13624 34623 13636 34632
rect 13630 34620 13636 34623
rect 13688 34620 13694 34672
rect 19512 34663 19570 34669
rect 19512 34629 19524 34663
rect 19558 34660 19570 34663
rect 20622 34660 20628 34672
rect 19558 34632 20628 34660
rect 19558 34629 19570 34632
rect 19512 34623 19570 34629
rect 20622 34620 20628 34632
rect 20680 34620 20686 34672
rect 23750 34660 23756 34672
rect 21836 34632 23756 34660
rect 8938 34592 8944 34604
rect 8899 34564 8944 34592
rect 8938 34552 8944 34564
rect 8996 34552 9002 34604
rect 9208 34595 9266 34601
rect 9208 34561 9220 34595
rect 9254 34592 9266 34595
rect 10318 34592 10324 34604
rect 9254 34564 10324 34592
rect 9254 34561 9266 34564
rect 9208 34555 9266 34561
rect 10318 34552 10324 34564
rect 10376 34552 10382 34604
rect 11784 34595 11842 34601
rect 11784 34561 11796 34595
rect 11830 34592 11842 34595
rect 15194 34592 15200 34604
rect 11830 34564 15200 34592
rect 11830 34561 11842 34564
rect 11784 34555 11842 34561
rect 15194 34552 15200 34564
rect 15252 34552 15258 34604
rect 16666 34552 16672 34604
rect 16724 34592 16730 34604
rect 16853 34595 16911 34601
rect 16853 34592 16865 34595
rect 16724 34564 16865 34592
rect 16724 34552 16730 34564
rect 16853 34561 16865 34564
rect 16899 34561 16911 34595
rect 16853 34555 16911 34561
rect 17120 34595 17178 34601
rect 17120 34561 17132 34595
rect 17166 34592 17178 34595
rect 18506 34592 18512 34604
rect 17166 34564 18512 34592
rect 17166 34561 17178 34564
rect 17120 34555 17178 34561
rect 18506 34552 18512 34564
rect 18564 34552 18570 34604
rect 21836 34601 21864 34632
rect 23750 34620 23756 34632
rect 23808 34620 23814 34672
rect 28442 34620 28448 34672
rect 28500 34660 28506 34672
rect 29058 34663 29116 34669
rect 29058 34660 29070 34663
rect 28500 34632 29070 34660
rect 28500 34620 28506 34632
rect 29058 34629 29070 34632
rect 29104 34629 29116 34663
rect 29058 34623 29116 34629
rect 34992 34632 37320 34660
rect 21821 34595 21879 34601
rect 21821 34561 21833 34595
rect 21867 34561 21879 34595
rect 21821 34555 21879 34561
rect 22088 34595 22146 34601
rect 22088 34561 22100 34595
rect 22134 34592 22146 34595
rect 23842 34592 23848 34604
rect 22134 34564 23848 34592
rect 22134 34561 22146 34564
rect 22088 34555 22146 34561
rect 23842 34552 23848 34564
rect 23900 34552 23906 34604
rect 24020 34595 24078 34601
rect 24020 34561 24032 34595
rect 24066 34592 24078 34595
rect 25038 34592 25044 34604
rect 24066 34564 25044 34592
rect 24066 34561 24078 34564
rect 24020 34555 24078 34561
rect 25038 34552 25044 34564
rect 25096 34552 25102 34604
rect 27240 34595 27298 34601
rect 27240 34561 27252 34595
rect 27286 34592 27298 34595
rect 28350 34592 28356 34604
rect 27286 34564 28356 34592
rect 27286 34561 27298 34564
rect 27240 34555 27298 34561
rect 28350 34552 28356 34564
rect 28408 34552 28414 34604
rect 28813 34595 28871 34601
rect 28813 34561 28825 34595
rect 28859 34592 28871 34595
rect 29914 34592 29920 34604
rect 28859 34564 29920 34592
rect 28859 34561 28871 34564
rect 28813 34555 28871 34561
rect 29914 34552 29920 34564
rect 29972 34552 29978 34604
rect 31754 34552 31760 34604
rect 31812 34592 31818 34604
rect 32122 34592 32128 34604
rect 31812 34564 32128 34592
rect 31812 34552 31818 34564
rect 32122 34552 32128 34564
rect 32180 34592 32186 34604
rect 33137 34595 33195 34601
rect 33137 34592 33149 34595
rect 32180 34564 33149 34592
rect 32180 34552 32186 34564
rect 33137 34561 33149 34564
rect 33183 34561 33195 34595
rect 33137 34555 33195 34561
rect 33404 34595 33462 34601
rect 33404 34561 33416 34595
rect 33450 34592 33462 34595
rect 34698 34592 34704 34604
rect 33450 34564 34704 34592
rect 33450 34561 33462 34564
rect 33404 34555 33462 34561
rect 34698 34552 34704 34564
rect 34756 34552 34762 34604
rect 10778 34484 10784 34536
rect 10836 34524 10842 34536
rect 11517 34527 11575 34533
rect 11517 34524 11529 34527
rect 10836 34496 11529 34524
rect 10836 34484 10842 34496
rect 11517 34493 11529 34496
rect 11563 34493 11575 34527
rect 11517 34487 11575 34493
rect 13078 34484 13084 34536
rect 13136 34524 13142 34536
rect 13357 34527 13415 34533
rect 13357 34524 13369 34527
rect 13136 34496 13369 34524
rect 13136 34484 13142 34496
rect 13357 34493 13369 34496
rect 13403 34493 13415 34527
rect 19242 34524 19248 34536
rect 19203 34496 19248 34524
rect 13357 34487 13415 34493
rect 19242 34484 19248 34496
rect 19300 34484 19306 34536
rect 23750 34524 23756 34536
rect 23711 34496 23756 34524
rect 23750 34484 23756 34496
rect 23808 34484 23814 34536
rect 26878 34484 26884 34536
rect 26936 34524 26942 34536
rect 26973 34527 27031 34533
rect 26973 34524 26985 34527
rect 26936 34496 26985 34524
rect 26936 34484 26942 34496
rect 26973 34493 26985 34496
rect 27019 34493 27031 34527
rect 26973 34487 27031 34493
rect 34606 34484 34612 34536
rect 34664 34524 34670 34536
rect 34992 34533 35020 34632
rect 35244 34595 35302 34601
rect 35244 34561 35256 34595
rect 35290 34592 35302 34595
rect 36078 34592 36084 34604
rect 35290 34564 36084 34592
rect 35290 34561 35302 34564
rect 35244 34555 35302 34561
rect 36078 34552 36084 34564
rect 36136 34552 36142 34604
rect 37292 34601 37320 34632
rect 37366 34620 37372 34672
rect 37424 34660 37430 34672
rect 37522 34663 37580 34669
rect 37522 34660 37534 34663
rect 37424 34632 37534 34660
rect 37424 34620 37430 34632
rect 37522 34629 37534 34632
rect 37568 34629 37580 34663
rect 37522 34623 37580 34629
rect 37734 34620 37740 34672
rect 37792 34620 37798 34672
rect 39384 34663 39442 34669
rect 39384 34629 39396 34663
rect 39430 34660 39442 34663
rect 41782 34660 41788 34672
rect 39430 34632 41788 34660
rect 39430 34629 39442 34632
rect 39384 34623 39442 34629
rect 41782 34620 41788 34632
rect 41840 34620 41846 34672
rect 44174 34660 44180 34672
rect 43640 34632 44180 34660
rect 37277 34595 37335 34601
rect 37277 34561 37289 34595
rect 37323 34592 37335 34595
rect 37752 34592 37780 34620
rect 43640 34601 43668 34632
rect 44174 34620 44180 34632
rect 44232 34620 44238 34672
rect 45756 34669 45784 34700
rect 46842 34688 46848 34700
rect 46900 34688 46906 34740
rect 48958 34728 48964 34740
rect 48919 34700 48964 34728
rect 48958 34688 48964 34700
rect 49016 34688 49022 34740
rect 45732 34663 45790 34669
rect 45732 34629 45744 34663
rect 45778 34629 45790 34663
rect 45732 34623 45790 34629
rect 49513 34663 49571 34669
rect 49513 34629 49525 34663
rect 49559 34660 49571 34663
rect 49786 34660 49792 34672
rect 49559 34632 49792 34660
rect 49559 34629 49571 34632
rect 49513 34623 49571 34629
rect 49786 34620 49792 34632
rect 49844 34620 49850 34672
rect 52748 34632 53512 34660
rect 37323 34564 37780 34592
rect 43625 34595 43683 34601
rect 37323 34561 37335 34564
rect 37277 34555 37335 34561
rect 43625 34561 43637 34595
rect 43671 34561 43683 34595
rect 43625 34555 43683 34561
rect 43892 34595 43950 34601
rect 43892 34561 43904 34595
rect 43938 34592 43950 34595
rect 46290 34592 46296 34604
rect 43938 34564 46296 34592
rect 43938 34561 43950 34564
rect 43892 34555 43950 34561
rect 46290 34552 46296 34564
rect 46348 34552 46354 34604
rect 47848 34595 47906 34601
rect 47848 34561 47860 34595
rect 47894 34592 47906 34595
rect 48958 34592 48964 34604
rect 47894 34564 48964 34592
rect 47894 34561 47906 34564
rect 47848 34555 47906 34561
rect 48958 34552 48964 34564
rect 49016 34552 49022 34604
rect 52748 34536 52776 34632
rect 53000 34595 53058 34601
rect 53000 34561 53012 34595
rect 53046 34592 53058 34595
rect 53374 34592 53380 34604
rect 53046 34564 53380 34592
rect 53046 34561 53058 34564
rect 53000 34555 53058 34561
rect 53374 34552 53380 34564
rect 53432 34552 53438 34604
rect 53484 34592 53512 34632
rect 54110 34620 54116 34672
rect 54168 34660 54174 34672
rect 54818 34663 54876 34669
rect 54818 34660 54830 34663
rect 54168 34632 54830 34660
rect 54168 34620 54174 34632
rect 54818 34629 54830 34632
rect 54864 34629 54876 34663
rect 54818 34623 54876 34629
rect 54573 34595 54631 34601
rect 54573 34592 54585 34595
rect 53484 34564 54585 34592
rect 54573 34561 54585 34564
rect 54619 34561 54631 34595
rect 54573 34555 54631 34561
rect 34977 34527 35035 34533
rect 34977 34524 34989 34527
rect 34664 34496 34989 34524
rect 34664 34484 34670 34496
rect 34977 34493 34989 34496
rect 35023 34493 35035 34527
rect 39117 34527 39175 34533
rect 39117 34524 39129 34527
rect 34977 34487 35035 34493
rect 39040 34496 39129 34524
rect 6362 34416 6368 34468
rect 6420 34456 6426 34468
rect 6822 34456 6828 34468
rect 6420 34428 6828 34456
rect 6420 34416 6426 34428
rect 6822 34416 6828 34428
rect 6880 34456 6886 34468
rect 8021 34459 8079 34465
rect 8021 34456 8033 34459
rect 6880 34428 8033 34456
rect 6880 34416 6886 34428
rect 8021 34425 8033 34428
rect 8067 34425 8079 34459
rect 8021 34419 8079 34425
rect 20622 34388 20628 34400
rect 20583 34360 20628 34388
rect 20622 34348 20628 34360
rect 20680 34348 20686 34400
rect 34517 34391 34575 34397
rect 34517 34357 34529 34391
rect 34563 34388 34575 34391
rect 34790 34388 34796 34400
rect 34563 34360 34796 34388
rect 34563 34357 34575 34360
rect 34517 34351 34575 34357
rect 34790 34348 34796 34360
rect 34848 34348 34854 34400
rect 37918 34348 37924 34400
rect 37976 34388 37982 34400
rect 39040 34388 39068 34496
rect 39117 34493 39129 34496
rect 39163 34493 39175 34527
rect 39117 34487 39175 34493
rect 44910 34484 44916 34536
rect 44968 34524 44974 34536
rect 45462 34524 45468 34536
rect 44968 34496 45468 34524
rect 44968 34484 44974 34496
rect 45462 34484 45468 34496
rect 45520 34484 45526 34536
rect 47578 34524 47584 34536
rect 47539 34496 47584 34524
rect 47578 34484 47584 34496
rect 47636 34484 47642 34536
rect 52730 34524 52736 34536
rect 52691 34496 52736 34524
rect 52730 34484 52736 34496
rect 52788 34484 52794 34536
rect 54018 34484 54024 34536
rect 54076 34524 54082 34536
rect 54076 34496 54156 34524
rect 54076 34484 54082 34496
rect 54128 34465 54156 34496
rect 54113 34459 54171 34465
rect 54113 34425 54125 34459
rect 54159 34425 54171 34459
rect 54113 34419 54171 34425
rect 39850 34388 39856 34400
rect 37976 34360 39856 34388
rect 37976 34348 37982 34360
rect 39850 34348 39856 34360
rect 39908 34348 39914 34400
rect 45002 34388 45008 34400
rect 44963 34360 45008 34388
rect 45002 34348 45008 34360
rect 45060 34348 45066 34400
rect 50154 34348 50160 34400
rect 50212 34388 50218 34400
rect 50801 34391 50859 34397
rect 50801 34388 50813 34391
rect 50212 34360 50813 34388
rect 50212 34348 50218 34360
rect 50801 34357 50813 34360
rect 50847 34357 50859 34391
rect 55950 34388 55956 34400
rect 55911 34360 55956 34388
rect 50801 34351 50859 34357
rect 55950 34348 55956 34360
rect 56008 34348 56014 34400
rect 1104 34298 59340 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 59340 34298
rect 1104 34224 59340 34246
rect 10318 34184 10324 34196
rect 10279 34156 10324 34184
rect 10318 34144 10324 34156
rect 10376 34144 10382 34196
rect 15286 34144 15292 34196
rect 15344 34184 15350 34196
rect 15473 34187 15531 34193
rect 15473 34184 15485 34187
rect 15344 34156 15485 34184
rect 15344 34144 15350 34156
rect 15473 34153 15485 34156
rect 15519 34153 15531 34187
rect 18506 34184 18512 34196
rect 18467 34156 18512 34184
rect 15473 34147 15531 34153
rect 18506 34144 18512 34156
rect 18564 34144 18570 34196
rect 21082 34144 21088 34196
rect 21140 34184 21146 34196
rect 21818 34184 21824 34196
rect 21140 34156 21824 34184
rect 21140 34144 21146 34156
rect 21818 34144 21824 34156
rect 21876 34184 21882 34196
rect 22373 34187 22431 34193
rect 22373 34184 22385 34187
rect 21876 34156 22385 34184
rect 21876 34144 21882 34156
rect 22373 34153 22385 34156
rect 22419 34153 22431 34187
rect 22373 34147 22431 34153
rect 26970 34144 26976 34196
rect 27028 34184 27034 34196
rect 27617 34187 27675 34193
rect 27617 34184 27629 34187
rect 27028 34156 27629 34184
rect 27028 34144 27034 34156
rect 27617 34153 27629 34156
rect 27663 34153 27675 34187
rect 27617 34147 27675 34153
rect 30929 34187 30987 34193
rect 30929 34153 30941 34187
rect 30975 34184 30987 34187
rect 31846 34184 31852 34196
rect 30975 34156 31852 34184
rect 30975 34153 30987 34156
rect 30929 34147 30987 34153
rect 31846 34144 31852 34156
rect 31904 34144 31910 34196
rect 36078 34184 36084 34196
rect 36039 34156 36084 34184
rect 36078 34144 36084 34156
rect 36136 34144 36142 34196
rect 50798 34144 50804 34196
rect 50856 34184 50862 34196
rect 51537 34187 51595 34193
rect 51537 34184 51549 34187
rect 50856 34156 51549 34184
rect 50856 34144 50862 34156
rect 51537 34153 51549 34156
rect 51583 34153 51595 34187
rect 53374 34184 53380 34196
rect 53335 34156 53380 34184
rect 51537 34147 51595 34153
rect 53374 34144 53380 34156
rect 53432 34144 53438 34196
rect 56594 34144 56600 34196
rect 56652 34184 56658 34196
rect 56689 34187 56747 34193
rect 56689 34184 56701 34187
rect 56652 34156 56701 34184
rect 56652 34144 56658 34156
rect 56689 34153 56701 34156
rect 56735 34153 56747 34187
rect 56689 34147 56747 34153
rect 8938 34048 8944 34060
rect 8899 34020 8944 34048
rect 8938 34008 8944 34020
rect 8996 34008 9002 34060
rect 16666 34008 16672 34060
rect 16724 34048 16730 34060
rect 17129 34051 17187 34057
rect 17129 34048 17141 34051
rect 16724 34020 17141 34048
rect 16724 34008 16730 34020
rect 17129 34017 17141 34020
rect 17175 34017 17187 34051
rect 17129 34011 17187 34017
rect 26234 34008 26240 34060
rect 26292 34048 26298 34060
rect 26292 34020 26337 34048
rect 26292 34008 26298 34020
rect 28902 34008 28908 34060
rect 28960 34048 28966 34060
rect 29549 34051 29607 34057
rect 29549 34048 29561 34051
rect 28960 34020 29561 34048
rect 28960 34008 28966 34020
rect 29549 34017 29561 34020
rect 29595 34017 29607 34051
rect 39850 34048 39856 34060
rect 39811 34020 39856 34048
rect 29549 34011 29607 34017
rect 39850 34008 39856 34020
rect 39908 34008 39914 34060
rect 57146 34048 57152 34060
rect 57107 34020 57152 34048
rect 57146 34008 57152 34020
rect 57204 34008 57210 34060
rect 3786 33940 3792 33992
rect 3844 33980 3850 33992
rect 4893 33983 4951 33989
rect 4893 33980 4905 33983
rect 3844 33952 4905 33980
rect 3844 33940 3850 33952
rect 4893 33949 4905 33952
rect 4939 33980 4951 33983
rect 6362 33980 6368 33992
rect 4939 33952 6368 33980
rect 4939 33949 4951 33952
rect 4893 33943 4951 33949
rect 6362 33940 6368 33952
rect 6420 33980 6426 33992
rect 6733 33983 6791 33989
rect 6733 33980 6745 33983
rect 6420 33952 6745 33980
rect 6420 33940 6426 33952
rect 6733 33949 6745 33952
rect 6779 33949 6791 33983
rect 8956 33980 8984 34008
rect 10778 33980 10784 33992
rect 8956 33952 10784 33980
rect 6733 33943 6791 33949
rect 10778 33940 10784 33952
rect 10836 33940 10842 33992
rect 13998 33940 14004 33992
rect 14056 33980 14062 33992
rect 14093 33983 14151 33989
rect 14093 33980 14105 33983
rect 14056 33952 14105 33980
rect 14056 33940 14062 33952
rect 14093 33949 14105 33952
rect 14139 33949 14151 33983
rect 14093 33943 14151 33949
rect 14360 33983 14418 33989
rect 14360 33949 14372 33983
rect 14406 33980 14418 33983
rect 15470 33980 15476 33992
rect 14406 33952 15476 33980
rect 14406 33949 14418 33952
rect 14360 33943 14418 33949
rect 15470 33940 15476 33952
rect 15528 33940 15534 33992
rect 19242 33980 19248 33992
rect 19203 33952 19248 33980
rect 19242 33940 19248 33952
rect 19300 33940 19306 33992
rect 19512 33983 19570 33989
rect 19512 33949 19524 33983
rect 19558 33980 19570 33983
rect 20622 33980 20628 33992
rect 19558 33952 20628 33980
rect 19558 33949 19570 33952
rect 19512 33943 19570 33949
rect 20622 33940 20628 33952
rect 20680 33940 20686 33992
rect 24394 33980 24400 33992
rect 24355 33952 24400 33980
rect 24394 33940 24400 33952
rect 24452 33940 24458 33992
rect 29822 33989 29828 33992
rect 29816 33943 29828 33989
rect 29880 33980 29886 33992
rect 31662 33980 31668 33992
rect 29880 33952 29916 33980
rect 31623 33952 31668 33980
rect 29822 33940 29828 33943
rect 29880 33940 29886 33952
rect 31662 33940 31668 33952
rect 31720 33940 31726 33992
rect 34606 33940 34612 33992
rect 34664 33980 34670 33992
rect 34701 33983 34759 33989
rect 34701 33980 34713 33983
rect 34664 33952 34713 33980
rect 34664 33940 34670 33952
rect 34701 33949 34713 33952
rect 34747 33949 34759 33983
rect 34701 33943 34759 33949
rect 34790 33940 34796 33992
rect 34848 33980 34854 33992
rect 34957 33983 35015 33989
rect 34957 33980 34969 33983
rect 34848 33952 34969 33980
rect 34848 33940 34854 33952
rect 34957 33949 34969 33952
rect 35003 33949 35015 33983
rect 37918 33980 37924 33992
rect 37879 33952 37924 33980
rect 34957 33943 35015 33949
rect 37918 33940 37924 33952
rect 37976 33940 37982 33992
rect 38188 33983 38246 33989
rect 38188 33949 38200 33983
rect 38234 33980 38246 33983
rect 39114 33980 39120 33992
rect 38234 33952 39120 33980
rect 38234 33949 38246 33952
rect 38188 33943 38246 33949
rect 39114 33940 39120 33952
rect 39172 33940 39178 33992
rect 42521 33983 42579 33989
rect 42521 33949 42533 33983
rect 42567 33980 42579 33983
rect 42610 33980 42616 33992
rect 42567 33952 42616 33980
rect 42567 33949 42579 33952
rect 42521 33943 42579 33949
rect 42610 33940 42616 33952
rect 42668 33940 42674 33992
rect 44910 33940 44916 33992
rect 44968 33980 44974 33992
rect 45005 33983 45063 33989
rect 45005 33980 45017 33983
rect 44968 33952 45017 33980
rect 44968 33940 44974 33952
rect 45005 33949 45017 33952
rect 45051 33949 45063 33983
rect 45005 33943 45063 33949
rect 46845 33983 46903 33989
rect 46845 33949 46857 33983
rect 46891 33980 46903 33983
rect 47578 33980 47584 33992
rect 46891 33952 47584 33980
rect 46891 33949 46903 33952
rect 46845 33943 46903 33949
rect 47578 33940 47584 33952
rect 47636 33980 47642 33992
rect 50154 33980 50160 33992
rect 47636 33952 50160 33980
rect 47636 33940 47642 33952
rect 50154 33940 50160 33952
rect 50212 33940 50218 33992
rect 51997 33983 52055 33989
rect 51997 33980 52009 33983
rect 51092 33952 52009 33980
rect 51092 33924 51120 33952
rect 51997 33949 52009 33952
rect 52043 33949 52055 33983
rect 51997 33943 52055 33949
rect 52086 33940 52092 33992
rect 52144 33980 52150 33992
rect 52253 33983 52311 33989
rect 52253 33980 52265 33983
rect 52144 33952 52265 33980
rect 52144 33940 52150 33952
rect 52253 33949 52265 33952
rect 52299 33949 52311 33983
rect 52253 33943 52311 33949
rect 55309 33983 55367 33989
rect 55309 33949 55321 33983
rect 55355 33949 55367 33983
rect 55309 33943 55367 33949
rect 55576 33983 55634 33989
rect 55576 33949 55588 33983
rect 55622 33980 55634 33983
rect 56686 33980 56692 33992
rect 55622 33952 56692 33980
rect 55622 33949 55634 33952
rect 55576 33943 55634 33949
rect 5160 33915 5218 33921
rect 5160 33881 5172 33915
rect 5206 33912 5218 33915
rect 5994 33912 6000 33924
rect 5206 33884 6000 33912
rect 5206 33881 5218 33884
rect 5160 33875 5218 33881
rect 5994 33872 6000 33884
rect 6052 33872 6058 33924
rect 7000 33915 7058 33921
rect 7000 33881 7012 33915
rect 7046 33912 7058 33915
rect 7742 33912 7748 33924
rect 7046 33884 7748 33912
rect 7046 33881 7058 33884
rect 7000 33875 7058 33881
rect 7742 33872 7748 33884
rect 7800 33872 7806 33924
rect 9208 33915 9266 33921
rect 9208 33881 9220 33915
rect 9254 33912 9266 33915
rect 10318 33912 10324 33924
rect 9254 33884 10324 33912
rect 9254 33881 9266 33884
rect 9208 33875 9266 33881
rect 10318 33872 10324 33884
rect 10376 33872 10382 33924
rect 11048 33915 11106 33921
rect 11048 33881 11060 33915
rect 11094 33912 11106 33915
rect 12066 33912 12072 33924
rect 11094 33884 12072 33912
rect 11094 33881 11106 33884
rect 11048 33875 11106 33881
rect 12066 33872 12072 33884
rect 12124 33872 12130 33924
rect 17396 33915 17454 33921
rect 17396 33881 17408 33915
rect 17442 33912 17454 33915
rect 18414 33912 18420 33924
rect 17442 33884 18420 33912
rect 17442 33881 17454 33884
rect 17396 33875 17454 33881
rect 18414 33872 18420 33884
rect 18472 33872 18478 33924
rect 20714 33872 20720 33924
rect 20772 33912 20778 33924
rect 21085 33915 21143 33921
rect 21085 33912 21097 33915
rect 20772 33884 21097 33912
rect 20772 33872 20778 33884
rect 21085 33881 21097 33884
rect 21131 33912 21143 33915
rect 24664 33915 24722 33921
rect 21131 33884 22508 33912
rect 21131 33881 21143 33884
rect 21085 33875 21143 33881
rect 6270 33844 6276 33856
rect 6231 33816 6276 33844
rect 6270 33804 6276 33816
rect 6328 33804 6334 33856
rect 8110 33844 8116 33856
rect 8071 33816 8116 33844
rect 8110 33804 8116 33816
rect 8168 33804 8174 33856
rect 12161 33847 12219 33853
rect 12161 33813 12173 33847
rect 12207 33844 12219 33847
rect 12526 33844 12532 33856
rect 12207 33816 12532 33844
rect 12207 33813 12219 33816
rect 12161 33807 12219 33813
rect 12526 33804 12532 33816
rect 12584 33804 12590 33856
rect 20622 33844 20628 33856
rect 20583 33816 20628 33844
rect 20622 33804 20628 33816
rect 20680 33804 20686 33856
rect 22480 33844 22508 33884
rect 24664 33881 24676 33915
rect 24710 33912 24722 33915
rect 25682 33912 25688 33924
rect 24710 33884 25688 33912
rect 24710 33881 24722 33884
rect 24664 33875 24722 33881
rect 25682 33872 25688 33884
rect 25740 33872 25746 33924
rect 26326 33872 26332 33924
rect 26384 33912 26390 33924
rect 26482 33915 26540 33921
rect 26482 33912 26494 33915
rect 26384 33884 26494 33912
rect 26384 33872 26390 33884
rect 26482 33881 26494 33884
rect 26528 33881 26540 33915
rect 26482 33875 26540 33881
rect 31932 33915 31990 33921
rect 31932 33881 31944 33915
rect 31978 33912 31990 33915
rect 33502 33912 33508 33924
rect 31978 33884 33508 33912
rect 31978 33881 31990 33884
rect 31932 33875 31990 33881
rect 33502 33872 33508 33884
rect 33560 33872 33566 33924
rect 39666 33872 39672 33924
rect 39724 33912 39730 33924
rect 40098 33915 40156 33921
rect 40098 33912 40110 33915
rect 39724 33884 40110 33912
rect 39724 33872 39730 33884
rect 40098 33881 40110 33884
rect 40144 33881 40156 33915
rect 40098 33875 40156 33881
rect 42788 33915 42846 33921
rect 42788 33881 42800 33915
rect 42834 33912 42846 33915
rect 43806 33912 43812 33924
rect 42834 33884 43812 33912
rect 42834 33881 42846 33884
rect 42788 33875 42846 33881
rect 43806 33872 43812 33884
rect 43864 33872 43870 33924
rect 45272 33915 45330 33921
rect 45272 33881 45284 33915
rect 45318 33912 45330 33915
rect 45554 33912 45560 33924
rect 45318 33884 45560 33912
rect 45318 33881 45330 33884
rect 45272 33875 45330 33881
rect 45554 33872 45560 33884
rect 45612 33872 45618 33924
rect 47112 33915 47170 33921
rect 47112 33881 47124 33915
rect 47158 33912 47170 33915
rect 48866 33912 48872 33924
rect 47158 33884 48872 33912
rect 47158 33881 47170 33884
rect 47112 33875 47170 33881
rect 48866 33872 48872 33884
rect 48924 33872 48930 33924
rect 50424 33915 50482 33921
rect 50424 33881 50436 33915
rect 50470 33912 50482 33915
rect 50798 33912 50804 33924
rect 50470 33884 50804 33912
rect 50470 33881 50482 33884
rect 50424 33875 50482 33881
rect 50798 33872 50804 33884
rect 50856 33872 50862 33924
rect 51074 33872 51080 33924
rect 51132 33872 51138 33924
rect 52730 33872 52736 33924
rect 52788 33912 52794 33924
rect 55324 33912 55352 33943
rect 56686 33940 56692 33952
rect 56744 33940 56750 33992
rect 57146 33912 57152 33924
rect 52788 33884 57152 33912
rect 52788 33872 52794 33884
rect 57146 33872 57152 33884
rect 57204 33872 57210 33924
rect 57416 33915 57474 33921
rect 57416 33881 57428 33915
rect 57462 33912 57474 33915
rect 58434 33912 58440 33924
rect 57462 33884 58440 33912
rect 57462 33881 57474 33884
rect 57416 33875 57474 33881
rect 58434 33872 58440 33884
rect 58492 33872 58498 33924
rect 24854 33844 24860 33856
rect 22480 33816 24860 33844
rect 24854 33804 24860 33816
rect 24912 33804 24918 33856
rect 25774 33844 25780 33856
rect 25735 33816 25780 33844
rect 25774 33804 25780 33816
rect 25832 33804 25838 33856
rect 33042 33844 33048 33856
rect 33003 33816 33048 33844
rect 33042 33804 33048 33816
rect 33100 33804 33106 33856
rect 39298 33844 39304 33856
rect 39259 33816 39304 33844
rect 39298 33804 39304 33816
rect 39356 33804 39362 33856
rect 40586 33804 40592 33856
rect 40644 33844 40650 33856
rect 41233 33847 41291 33853
rect 41233 33844 41245 33847
rect 40644 33816 41245 33844
rect 40644 33804 40650 33816
rect 41233 33813 41245 33816
rect 41279 33813 41291 33847
rect 43898 33844 43904 33856
rect 43859 33816 43904 33844
rect 41233 33807 41291 33813
rect 43898 33804 43904 33816
rect 43956 33804 43962 33856
rect 46382 33844 46388 33856
rect 46343 33816 46388 33844
rect 46382 33804 46388 33816
rect 46440 33804 46446 33856
rect 48222 33844 48228 33856
rect 48183 33816 48228 33844
rect 48222 33804 48228 33816
rect 48280 33804 48286 33856
rect 58526 33844 58532 33856
rect 58487 33816 58532 33844
rect 58526 33804 58532 33816
rect 58584 33804 58590 33856
rect 1104 33754 59340 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 59340 33754
rect 1104 33680 59340 33702
rect 7742 33640 7748 33652
rect 7703 33612 7748 33640
rect 7742 33600 7748 33612
rect 7800 33600 7806 33652
rect 9582 33640 9588 33652
rect 9543 33612 9588 33640
rect 9582 33600 9588 33612
rect 9640 33600 9646 33652
rect 18414 33640 18420 33652
rect 18375 33612 18420 33640
rect 18414 33600 18420 33612
rect 18472 33600 18478 33652
rect 25038 33640 25044 33652
rect 24999 33612 25044 33640
rect 25038 33600 25044 33612
rect 25096 33600 25102 33652
rect 28350 33640 28356 33652
rect 28311 33612 28356 33640
rect 28350 33600 28356 33612
rect 28408 33600 28414 33652
rect 33502 33640 33508 33652
rect 33463 33612 33508 33640
rect 33502 33600 33508 33612
rect 33560 33600 33566 33652
rect 34698 33600 34704 33652
rect 34756 33640 34762 33652
rect 35345 33643 35403 33649
rect 35345 33640 35357 33643
rect 34756 33612 35357 33640
rect 34756 33600 34762 33612
rect 35345 33609 35357 33612
rect 35391 33609 35403 33643
rect 39666 33640 39672 33652
rect 39627 33612 39672 33640
rect 35345 33603 35403 33609
rect 39666 33600 39672 33612
rect 39724 33600 39730 33652
rect 43806 33640 43812 33652
rect 43767 33612 43812 33640
rect 43806 33600 43812 33612
rect 43864 33600 43870 33652
rect 48958 33640 48964 33652
rect 48919 33612 48964 33640
rect 48958 33600 48964 33612
rect 49016 33600 49022 33652
rect 50798 33640 50804 33652
rect 50759 33612 50804 33640
rect 50798 33600 50804 33612
rect 50856 33600 50862 33652
rect 53926 33600 53932 33652
rect 53984 33640 53990 33652
rect 54113 33643 54171 33649
rect 54113 33640 54125 33643
rect 53984 33612 54125 33640
rect 53984 33600 53990 33612
rect 54113 33609 54125 33612
rect 54159 33609 54171 33643
rect 54113 33603 54171 33609
rect 6270 33532 6276 33584
rect 6328 33572 6334 33584
rect 6610 33575 6668 33581
rect 6610 33572 6622 33575
rect 6328 33544 6622 33572
rect 6328 33532 6334 33544
rect 6610 33541 6622 33544
rect 6656 33541 6668 33575
rect 6610 33535 6668 33541
rect 8472 33575 8530 33581
rect 8472 33541 8484 33575
rect 8518 33572 8530 33575
rect 8570 33572 8576 33584
rect 8518 33544 8576 33572
rect 8518 33541 8530 33544
rect 8472 33535 8530 33541
rect 8570 33532 8576 33544
rect 8628 33532 8634 33584
rect 11882 33572 11888 33584
rect 11795 33544 11888 33572
rect 11882 33532 11888 33544
rect 11940 33572 11946 33584
rect 13354 33572 13360 33584
rect 11940 33544 13360 33572
rect 11940 33532 11946 33544
rect 13354 33532 13360 33544
rect 13412 33532 13418 33584
rect 19242 33572 19248 33584
rect 17052 33544 19248 33572
rect 4332 33507 4390 33513
rect 4332 33473 4344 33507
rect 4378 33504 4390 33507
rect 5166 33504 5172 33516
rect 4378 33476 5172 33504
rect 4378 33473 4390 33476
rect 4332 33467 4390 33473
rect 5166 33464 5172 33476
rect 5224 33464 5230 33516
rect 6362 33504 6368 33516
rect 6323 33476 6368 33504
rect 6362 33464 6368 33476
rect 6420 33504 6426 33516
rect 6914 33504 6920 33516
rect 6420 33476 6920 33504
rect 6420 33464 6426 33476
rect 6914 33464 6920 33476
rect 6972 33464 6978 33516
rect 8205 33507 8263 33513
rect 8205 33473 8217 33507
rect 8251 33504 8263 33507
rect 8938 33504 8944 33516
rect 8251 33476 8944 33504
rect 8251 33473 8263 33476
rect 8205 33467 8263 33473
rect 8938 33464 8944 33476
rect 8996 33464 9002 33516
rect 14360 33507 14418 33513
rect 14360 33473 14372 33507
rect 14406 33504 14418 33507
rect 14734 33504 14740 33516
rect 14406 33476 14740 33504
rect 14406 33473 14418 33476
rect 14360 33467 14418 33473
rect 14734 33464 14740 33476
rect 14792 33464 14798 33516
rect 17052 33513 17080 33544
rect 19242 33532 19248 33544
rect 19300 33532 19306 33584
rect 19512 33575 19570 33581
rect 19512 33541 19524 33575
rect 19558 33572 19570 33575
rect 20622 33572 20628 33584
rect 19558 33544 20628 33572
rect 19558 33541 19570 33544
rect 19512 33535 19570 33541
rect 20622 33532 20628 33544
rect 20680 33532 20686 33584
rect 23928 33575 23986 33581
rect 23928 33541 23940 33575
rect 23974 33572 23986 33575
rect 25774 33572 25780 33584
rect 23974 33544 25780 33572
rect 23974 33541 23986 33544
rect 23928 33535 23986 33541
rect 25774 33532 25780 33544
rect 25832 33532 25838 33584
rect 26602 33532 26608 33584
rect 26660 33572 26666 33584
rect 27218 33575 27276 33581
rect 27218 33572 27230 33575
rect 26660 33544 27230 33572
rect 26660 33532 26666 33544
rect 27218 33541 27230 33544
rect 27264 33541 27276 33575
rect 27218 33535 27276 33541
rect 30092 33575 30150 33581
rect 30092 33541 30104 33575
rect 30138 33572 30150 33575
rect 30374 33572 30380 33584
rect 30138 33544 30380 33572
rect 30138 33541 30150 33544
rect 30092 33535 30150 33541
rect 30374 33532 30380 33544
rect 30432 33532 30438 33584
rect 38556 33575 38614 33581
rect 38556 33541 38568 33575
rect 38602 33572 38614 33575
rect 39298 33572 39304 33584
rect 38602 33544 39304 33572
rect 38602 33541 38614 33544
rect 38556 33535 38614 33541
rect 39298 33532 39304 33544
rect 39356 33532 39362 33584
rect 40126 33572 40132 33584
rect 40087 33544 40132 33572
rect 40126 33532 40132 33544
rect 40184 33532 40190 33584
rect 43898 33532 43904 33584
rect 43956 33572 43962 33584
rect 44514 33575 44572 33581
rect 44514 33572 44526 33575
rect 43956 33544 44526 33572
rect 43956 33532 43962 33544
rect 44514 33541 44526 33544
rect 44560 33541 44572 33575
rect 44514 33535 44572 33541
rect 47848 33575 47906 33581
rect 47848 33541 47860 33575
rect 47894 33572 47906 33575
rect 48222 33572 48228 33584
rect 47894 33544 48228 33572
rect 47894 33541 47906 33544
rect 47848 33535 47906 33541
rect 48222 33532 48228 33544
rect 48280 33532 48286 33584
rect 49694 33581 49700 33584
rect 49688 33572 49700 33581
rect 49655 33544 49700 33572
rect 49688 33535 49700 33544
rect 49694 33532 49700 33535
rect 49752 33532 49758 33584
rect 53006 33581 53012 33584
rect 53000 33572 53012 33581
rect 52967 33544 53012 33572
rect 53000 33535 53012 33544
rect 53006 33532 53012 33535
rect 53064 33532 53070 33584
rect 54662 33532 54668 33584
rect 54720 33572 54726 33584
rect 54757 33575 54815 33581
rect 54757 33572 54769 33575
rect 54720 33544 54769 33572
rect 54720 33532 54726 33544
rect 54757 33541 54769 33544
rect 54803 33541 54815 33575
rect 54757 33535 54815 33541
rect 56505 33575 56563 33581
rect 56505 33541 56517 33575
rect 56551 33572 56563 33575
rect 57146 33572 57152 33584
rect 56551 33544 57152 33572
rect 56551 33541 56563 33544
rect 56505 33535 56563 33541
rect 57146 33532 57152 33544
rect 57204 33532 57210 33584
rect 17037 33507 17095 33513
rect 17037 33473 17049 33507
rect 17083 33473 17095 33507
rect 17037 33467 17095 33473
rect 17304 33507 17362 33513
rect 17304 33473 17316 33507
rect 17350 33504 17362 33507
rect 18874 33504 18880 33516
rect 17350 33476 18880 33504
rect 17350 33473 17362 33476
rect 17304 33467 17362 33473
rect 18874 33464 18880 33476
rect 18932 33464 18938 33516
rect 21818 33504 21824 33516
rect 21779 33476 21824 33504
rect 21818 33464 21824 33476
rect 21876 33464 21882 33516
rect 22094 33513 22100 33516
rect 22088 33467 22100 33513
rect 22152 33504 22158 33516
rect 23661 33507 23719 33513
rect 22152 33476 22188 33504
rect 22094 33464 22100 33467
rect 22152 33464 22158 33476
rect 23661 33473 23673 33507
rect 23707 33504 23719 33507
rect 23750 33504 23756 33516
rect 23707 33476 23756 33504
rect 23707 33473 23719 33476
rect 23661 33467 23719 33473
rect 23750 33464 23756 33476
rect 23808 33504 23814 33516
rect 24394 33504 24400 33516
rect 23808 33476 24400 33504
rect 23808 33464 23814 33476
rect 24394 33464 24400 33476
rect 24452 33464 24458 33516
rect 29825 33507 29883 33513
rect 29825 33473 29837 33507
rect 29871 33504 29883 33507
rect 29914 33504 29920 33516
rect 29871 33476 29920 33504
rect 29871 33473 29883 33476
rect 29825 33467 29883 33473
rect 29914 33464 29920 33476
rect 29972 33464 29978 33516
rect 31754 33464 31760 33516
rect 31812 33504 31818 33516
rect 32381 33507 32439 33513
rect 32381 33504 32393 33507
rect 31812 33476 32393 33504
rect 31812 33464 31818 33476
rect 32381 33473 32393 33476
rect 32427 33473 32439 33507
rect 32381 33467 32439 33473
rect 33870 33464 33876 33516
rect 33928 33504 33934 33516
rect 34221 33507 34279 33513
rect 34221 33504 34233 33507
rect 33928 33476 34233 33504
rect 33928 33464 33934 33476
rect 34221 33473 34233 33476
rect 34267 33473 34279 33507
rect 34221 33467 34279 33473
rect 42696 33507 42754 33513
rect 42696 33473 42708 33507
rect 42742 33504 42754 33507
rect 43806 33504 43812 33516
rect 42742 33476 43812 33504
rect 42742 33473 42754 33476
rect 42696 33467 42754 33473
rect 43806 33464 43812 33476
rect 43864 33464 43870 33516
rect 49421 33507 49479 33513
rect 49421 33504 49433 33507
rect 47596 33476 49433 33504
rect 47596 33448 47624 33476
rect 49421 33473 49433 33476
rect 49467 33473 49479 33507
rect 49421 33467 49479 33473
rect 3786 33396 3792 33448
rect 3844 33436 3850 33448
rect 4065 33439 4123 33445
rect 4065 33436 4077 33439
rect 3844 33408 4077 33436
rect 3844 33396 3850 33408
rect 4065 33405 4077 33408
rect 4111 33405 4123 33439
rect 4065 33399 4123 33405
rect 13998 33396 14004 33448
rect 14056 33436 14062 33448
rect 14093 33439 14151 33445
rect 14093 33436 14105 33439
rect 14056 33408 14105 33436
rect 14056 33396 14062 33408
rect 14093 33405 14105 33408
rect 14139 33405 14151 33439
rect 19242 33436 19248 33448
rect 19203 33408 19248 33436
rect 14093 33399 14151 33405
rect 19242 33396 19248 33408
rect 19300 33396 19306 33448
rect 26970 33436 26976 33448
rect 26931 33408 26976 33436
rect 26970 33396 26976 33408
rect 27028 33396 27034 33448
rect 32122 33436 32128 33448
rect 32083 33408 32128 33436
rect 32122 33396 32128 33408
rect 32180 33396 32186 33448
rect 33965 33439 34023 33445
rect 33965 33405 33977 33439
rect 34011 33405 34023 33439
rect 33965 33399 34023 33405
rect 20530 33328 20536 33380
rect 20588 33368 20594 33380
rect 20625 33371 20683 33377
rect 20625 33368 20637 33371
rect 20588 33340 20637 33368
rect 20588 33328 20594 33340
rect 20625 33337 20637 33340
rect 20671 33337 20683 33371
rect 20625 33331 20683 33337
rect 5445 33303 5503 33309
rect 5445 33269 5457 33303
rect 5491 33300 5503 33303
rect 5902 33300 5908 33312
rect 5491 33272 5908 33300
rect 5491 33269 5503 33272
rect 5445 33263 5503 33269
rect 5902 33260 5908 33272
rect 5960 33260 5966 33312
rect 13078 33260 13084 33312
rect 13136 33300 13142 33312
rect 13173 33303 13231 33309
rect 13173 33300 13185 33303
rect 13136 33272 13185 33300
rect 13136 33260 13142 33272
rect 13173 33269 13185 33272
rect 13219 33269 13231 33303
rect 15470 33300 15476 33312
rect 15431 33272 15476 33300
rect 13173 33263 13231 33269
rect 15470 33260 15476 33272
rect 15528 33260 15534 33312
rect 23198 33300 23204 33312
rect 23159 33272 23204 33300
rect 23198 33260 23204 33272
rect 23256 33260 23262 33312
rect 31202 33300 31208 33312
rect 31163 33272 31208 33300
rect 31202 33260 31208 33272
rect 31260 33260 31266 33312
rect 31662 33260 31668 33312
rect 31720 33300 31726 33312
rect 33980 33300 34008 33399
rect 37918 33396 37924 33448
rect 37976 33436 37982 33448
rect 38289 33439 38347 33445
rect 38289 33436 38301 33439
rect 37976 33408 38301 33436
rect 37976 33396 37982 33408
rect 38289 33405 38301 33408
rect 38335 33405 38347 33439
rect 42150 33436 42156 33448
rect 38289 33399 38347 33405
rect 41432 33408 42156 33436
rect 34698 33300 34704 33312
rect 31720 33272 34704 33300
rect 31720 33260 31726 33272
rect 34698 33260 34704 33272
rect 34756 33260 34762 33312
rect 39850 33260 39856 33312
rect 39908 33300 39914 33312
rect 41432 33309 41460 33408
rect 42150 33396 42156 33408
rect 42208 33436 42214 33448
rect 42429 33439 42487 33445
rect 42429 33436 42441 33439
rect 42208 33408 42441 33436
rect 42208 33396 42214 33408
rect 42429 33405 42441 33408
rect 42475 33405 42487 33439
rect 42429 33399 42487 33405
rect 44174 33396 44180 33448
rect 44232 33436 44238 33448
rect 44269 33439 44327 33445
rect 44269 33436 44281 33439
rect 44232 33408 44281 33436
rect 44232 33396 44238 33408
rect 44269 33405 44281 33408
rect 44315 33405 44327 33439
rect 47578 33436 47584 33448
rect 47539 33408 47584 33436
rect 44269 33399 44327 33405
rect 47578 33396 47584 33408
rect 47636 33396 47642 33448
rect 51074 33396 51080 33448
rect 51132 33436 51138 33448
rect 52730 33436 52736 33448
rect 51132 33408 52736 33436
rect 51132 33396 51138 33408
rect 52730 33396 52736 33408
rect 52788 33396 52794 33448
rect 41417 33303 41475 33309
rect 41417 33300 41429 33303
rect 39908 33272 41429 33300
rect 39908 33260 39914 33272
rect 41417 33269 41429 33272
rect 41463 33269 41475 33303
rect 45646 33300 45652 33312
rect 45607 33272 45652 33300
rect 41417 33263 41475 33269
rect 45646 33260 45652 33272
rect 45704 33260 45710 33312
rect 1104 33210 59340 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 59340 33210
rect 1104 33136 59340 33158
rect 5166 33096 5172 33108
rect 5127 33068 5172 33096
rect 5166 33056 5172 33068
rect 5224 33056 5230 33108
rect 5994 33056 6000 33108
rect 6052 33096 6058 33108
rect 7009 33099 7067 33105
rect 7009 33096 7021 33099
rect 6052 33068 7021 33096
rect 6052 33056 6058 33068
rect 7009 33065 7021 33068
rect 7055 33065 7067 33099
rect 10318 33096 10324 33108
rect 10279 33068 10324 33096
rect 7009 33059 7067 33065
rect 10318 33056 10324 33068
rect 10376 33056 10382 33108
rect 12066 33056 12072 33108
rect 12124 33096 12130 33108
rect 12161 33099 12219 33105
rect 12161 33096 12173 33099
rect 12124 33068 12173 33096
rect 12124 33056 12130 33068
rect 12161 33065 12173 33068
rect 12207 33065 12219 33099
rect 12161 33059 12219 33065
rect 20993 33099 21051 33105
rect 20993 33065 21005 33099
rect 21039 33096 21051 33099
rect 22094 33096 22100 33108
rect 21039 33068 22100 33096
rect 21039 33065 21051 33068
rect 20993 33059 21051 33065
rect 22094 33056 22100 33068
rect 22152 33056 22158 33108
rect 22830 33096 22836 33108
rect 22791 33068 22836 33096
rect 22830 33056 22836 33068
rect 22888 33056 22894 33108
rect 25777 33099 25835 33105
rect 25777 33065 25789 33099
rect 25823 33096 25835 33099
rect 26326 33096 26332 33108
rect 25823 33068 26332 33096
rect 25823 33065 25835 33068
rect 25777 33059 25835 33065
rect 26326 33056 26332 33068
rect 26384 33056 26390 33108
rect 36173 33099 36231 33105
rect 36173 33065 36185 33099
rect 36219 33096 36231 33099
rect 36998 33096 37004 33108
rect 36219 33068 37004 33096
rect 36219 33065 36231 33068
rect 36173 33059 36231 33065
rect 36998 33056 37004 33068
rect 37056 33056 37062 33108
rect 46290 33056 46296 33108
rect 46348 33096 46354 33108
rect 46385 33099 46443 33105
rect 46385 33096 46397 33099
rect 46348 33068 46397 33096
rect 46348 33056 46354 33068
rect 46385 33065 46397 33068
rect 46431 33065 46443 33099
rect 46385 33059 46443 33065
rect 51902 33056 51908 33108
rect 51960 33096 51966 33108
rect 52273 33099 52331 33105
rect 52273 33096 52285 33099
rect 51960 33068 52285 33096
rect 51960 33056 51966 33068
rect 52273 33065 52285 33068
rect 52319 33065 52331 33099
rect 52273 33059 52331 33065
rect 56689 33099 56747 33105
rect 56689 33065 56701 33099
rect 56735 33096 56747 33099
rect 56778 33096 56784 33108
rect 56735 33068 56784 33096
rect 56735 33065 56747 33068
rect 56689 33059 56747 33065
rect 56778 33056 56784 33068
rect 56836 33056 56842 33108
rect 58434 33056 58440 33108
rect 58492 33096 58498 33108
rect 58529 33099 58587 33105
rect 58529 33096 58541 33099
rect 58492 33068 58541 33096
rect 58492 33056 58498 33068
rect 58529 33065 58541 33068
rect 58575 33065 58587 33099
rect 58529 33059 58587 33065
rect 8938 32960 8944 32972
rect 8899 32932 8944 32960
rect 8938 32920 8944 32932
rect 8996 32920 9002 32972
rect 13998 32920 14004 32972
rect 14056 32960 14062 32972
rect 14829 32963 14887 32969
rect 14829 32960 14841 32963
rect 14056 32932 14841 32960
rect 14056 32920 14062 32932
rect 14829 32929 14841 32932
rect 14875 32929 14887 32963
rect 16666 32960 16672 32972
rect 16627 32932 16672 32960
rect 14829 32923 14887 32929
rect 16666 32920 16672 32932
rect 16724 32920 16730 32972
rect 29914 32960 29920 32972
rect 29875 32932 29920 32960
rect 29914 32920 29920 32932
rect 29972 32920 29978 32972
rect 39850 32920 39856 32972
rect 39908 32960 39914 32972
rect 40313 32963 40371 32969
rect 40313 32960 40325 32963
rect 39908 32932 40325 32960
rect 39908 32920 39914 32932
rect 40313 32929 40325 32932
rect 40359 32929 40371 32963
rect 42150 32960 42156 32972
rect 42111 32932 42156 32960
rect 40313 32923 40371 32929
rect 42150 32920 42156 32932
rect 42208 32920 42214 32972
rect 52730 32920 52736 32972
rect 52788 32960 52794 32972
rect 53377 32963 53435 32969
rect 53377 32960 53389 32963
rect 52788 32932 53389 32960
rect 52788 32920 52794 32932
rect 53377 32929 53389 32932
rect 53423 32929 53435 32963
rect 57146 32960 57152 32972
rect 57107 32932 57152 32960
rect 53377 32923 53435 32929
rect 3326 32852 3332 32904
rect 3384 32892 3390 32904
rect 3786 32892 3792 32904
rect 3384 32864 3792 32892
rect 3384 32852 3390 32864
rect 3786 32852 3792 32864
rect 3844 32852 3850 32904
rect 5629 32895 5687 32901
rect 5629 32861 5641 32895
rect 5675 32892 5687 32895
rect 8956 32892 8984 32920
rect 10226 32892 10232 32904
rect 5675 32864 6316 32892
rect 8956 32864 10232 32892
rect 5675 32861 5687 32864
rect 5629 32855 5687 32861
rect 4056 32827 4114 32833
rect 4056 32793 4068 32827
rect 4102 32824 4114 32827
rect 4706 32824 4712 32836
rect 4102 32796 4712 32824
rect 4102 32793 4114 32796
rect 4056 32787 4114 32793
rect 4706 32784 4712 32796
rect 4764 32784 4770 32836
rect 5902 32833 5908 32836
rect 5896 32824 5908 32833
rect 5863 32796 5908 32824
rect 5896 32787 5908 32796
rect 5902 32784 5908 32787
rect 5960 32784 5966 32836
rect 6288 32824 6316 32864
rect 10226 32852 10232 32864
rect 10284 32892 10290 32904
rect 11054 32901 11060 32904
rect 10781 32895 10839 32901
rect 10781 32892 10793 32895
rect 10284 32864 10793 32892
rect 10284 32852 10290 32864
rect 10781 32861 10793 32864
rect 10827 32861 10839 32895
rect 11048 32892 11060 32901
rect 11015 32864 11060 32892
rect 10781 32855 10839 32861
rect 11048 32855 11060 32864
rect 11054 32852 11060 32855
rect 11112 32852 11118 32904
rect 19242 32852 19248 32904
rect 19300 32892 19306 32904
rect 19613 32895 19671 32901
rect 19613 32892 19625 32895
rect 19300 32864 19625 32892
rect 19300 32852 19306 32864
rect 19613 32861 19625 32864
rect 19659 32861 19671 32895
rect 19613 32855 19671 32861
rect 19880 32895 19938 32901
rect 19880 32861 19892 32895
rect 19926 32892 19938 32895
rect 20162 32892 20168 32904
rect 19926 32864 20168 32892
rect 19926 32861 19938 32864
rect 19880 32855 19938 32861
rect 6914 32824 6920 32836
rect 6288 32796 6920 32824
rect 6914 32784 6920 32796
rect 6972 32784 6978 32836
rect 9208 32827 9266 32833
rect 9208 32793 9220 32827
rect 9254 32824 9266 32827
rect 9582 32824 9588 32836
rect 9254 32796 9588 32824
rect 9254 32793 9266 32796
rect 9208 32787 9266 32793
rect 9582 32784 9588 32796
rect 9640 32784 9646 32836
rect 15096 32827 15154 32833
rect 15096 32793 15108 32827
rect 15142 32824 15154 32827
rect 16574 32824 16580 32836
rect 15142 32796 16580 32824
rect 15142 32793 15154 32796
rect 15096 32787 15154 32793
rect 16574 32784 16580 32796
rect 16632 32784 16638 32836
rect 16936 32827 16994 32833
rect 16936 32793 16948 32827
rect 16982 32824 16994 32827
rect 17954 32824 17960 32836
rect 16982 32796 17960 32824
rect 16982 32793 16994 32796
rect 16936 32787 16994 32793
rect 17954 32784 17960 32796
rect 18012 32784 18018 32836
rect 19628 32824 19656 32855
rect 20162 32852 20168 32864
rect 20220 32852 20226 32904
rect 21453 32895 21511 32901
rect 21453 32861 21465 32895
rect 21499 32861 21511 32895
rect 21453 32855 21511 32861
rect 21720 32895 21778 32901
rect 21720 32861 21732 32895
rect 21766 32892 21778 32895
rect 23198 32892 23204 32904
rect 21766 32864 23204 32892
rect 21766 32861 21778 32864
rect 21720 32855 21778 32861
rect 21468 32824 21496 32855
rect 23198 32852 23204 32864
rect 23256 32852 23262 32904
rect 24394 32892 24400 32904
rect 24307 32864 24400 32892
rect 24394 32852 24400 32864
rect 24452 32852 24458 32904
rect 24670 32901 24676 32904
rect 24664 32892 24676 32901
rect 24631 32864 24676 32892
rect 24664 32855 24676 32864
rect 24670 32852 24676 32855
rect 24728 32852 24734 32904
rect 26970 32892 26976 32904
rect 26883 32864 26976 32892
rect 26970 32852 26976 32864
rect 27028 32892 27034 32904
rect 27522 32892 27528 32904
rect 27028 32864 27528 32892
rect 27028 32852 27034 32864
rect 27522 32852 27528 32864
rect 27580 32852 27586 32904
rect 30184 32895 30242 32901
rect 30184 32861 30196 32895
rect 30230 32892 30242 32895
rect 31202 32892 31208 32904
rect 30230 32864 31208 32892
rect 30230 32861 30242 32864
rect 30184 32855 30242 32861
rect 31202 32852 31208 32864
rect 31260 32852 31266 32904
rect 31941 32895 31999 32901
rect 31941 32861 31953 32895
rect 31987 32861 31999 32895
rect 31941 32855 31999 32861
rect 32208 32895 32266 32901
rect 32208 32861 32220 32895
rect 32254 32892 32266 32895
rect 33042 32892 33048 32904
rect 32254 32864 33048 32892
rect 32254 32861 32266 32864
rect 32208 32855 32266 32861
rect 21818 32824 21824 32836
rect 19628 32796 21824 32824
rect 21818 32784 21824 32796
rect 21876 32784 21882 32836
rect 23290 32784 23296 32836
rect 23348 32824 23354 32836
rect 24412 32824 24440 32852
rect 25038 32824 25044 32836
rect 23348 32796 25044 32824
rect 23348 32784 23354 32796
rect 25038 32784 25044 32796
rect 25096 32824 25102 32836
rect 26988 32824 27016 32852
rect 25096 32796 27016 32824
rect 27240 32827 27298 32833
rect 25096 32784 25102 32796
rect 27240 32793 27252 32827
rect 27286 32824 27298 32827
rect 28626 32824 28632 32836
rect 27286 32796 28632 32824
rect 27286 32793 27298 32796
rect 27240 32787 27298 32793
rect 28626 32784 28632 32796
rect 28684 32784 28690 32836
rect 31956 32824 31984 32855
rect 33042 32852 33048 32864
rect 33100 32852 33106 32904
rect 34793 32895 34851 32901
rect 34793 32861 34805 32895
rect 34839 32892 34851 32895
rect 35894 32892 35900 32904
rect 34839 32864 35900 32892
rect 34839 32861 34851 32864
rect 34793 32855 34851 32861
rect 35894 32852 35900 32864
rect 35952 32892 35958 32904
rect 40586 32901 40592 32904
rect 36633 32895 36691 32901
rect 36633 32892 36645 32895
rect 35952 32864 36645 32892
rect 35952 32852 35958 32864
rect 36633 32861 36645 32864
rect 36679 32861 36691 32895
rect 40580 32892 40592 32901
rect 40547 32864 40592 32892
rect 36633 32855 36691 32861
rect 40580 32855 40592 32864
rect 40586 32852 40592 32855
rect 40644 32852 40650 32904
rect 45005 32895 45063 32901
rect 45005 32861 45017 32895
rect 45051 32861 45063 32895
rect 45005 32855 45063 32861
rect 45272 32895 45330 32901
rect 45272 32861 45284 32895
rect 45318 32892 45330 32895
rect 45646 32892 45652 32904
rect 45318 32864 45652 32892
rect 45318 32861 45330 32864
rect 45272 32855 45330 32861
rect 32122 32824 32128 32836
rect 31956 32796 32128 32824
rect 32122 32784 32128 32796
rect 32180 32784 32186 32836
rect 34606 32784 34612 32836
rect 34664 32824 34670 32836
rect 35038 32827 35096 32833
rect 35038 32824 35050 32827
rect 34664 32796 35050 32824
rect 34664 32784 34670 32796
rect 35038 32793 35050 32796
rect 35084 32793 35096 32827
rect 35038 32787 35096 32793
rect 36900 32827 36958 32833
rect 36900 32793 36912 32827
rect 36946 32824 36958 32827
rect 38654 32824 38660 32836
rect 36946 32796 38660 32824
rect 36946 32793 36958 32796
rect 36900 32787 36958 32793
rect 38654 32784 38660 32796
rect 38712 32784 38718 32836
rect 41782 32784 41788 32836
rect 41840 32824 41846 32836
rect 42398 32827 42456 32833
rect 42398 32824 42410 32827
rect 41840 32796 42410 32824
rect 41840 32784 41846 32796
rect 42398 32793 42410 32796
rect 42444 32793 42456 32827
rect 45020 32824 45048 32855
rect 45646 32852 45652 32864
rect 45704 32852 45710 32904
rect 46845 32895 46903 32901
rect 46845 32892 46857 32895
rect 46400 32864 46857 32892
rect 46400 32824 46428 32864
rect 46845 32861 46857 32864
rect 46891 32892 46903 32895
rect 47578 32892 47584 32904
rect 46891 32864 47584 32892
rect 46891 32861 46903 32864
rect 46845 32855 46903 32861
rect 47578 32852 47584 32864
rect 47636 32852 47642 32904
rect 50798 32852 50804 32904
rect 50856 32892 50862 32904
rect 50893 32895 50951 32901
rect 50893 32892 50905 32895
rect 50856 32864 50905 32892
rect 50856 32852 50862 32864
rect 50893 32861 50905 32864
rect 50939 32892 50951 32895
rect 50982 32892 50988 32904
rect 50939 32864 50988 32892
rect 50939 32861 50951 32864
rect 50893 32855 50951 32861
rect 50982 32852 50988 32864
rect 51040 32852 51046 32904
rect 51166 32901 51172 32904
rect 51160 32892 51172 32901
rect 51127 32864 51172 32892
rect 51160 32855 51172 32864
rect 51166 32852 51172 32855
rect 51224 32852 51230 32904
rect 53392 32892 53420 32923
rect 57146 32920 57152 32932
rect 57204 32920 57210 32972
rect 55309 32895 55367 32901
rect 55309 32892 55321 32895
rect 53392 32864 55321 32892
rect 55309 32861 55321 32864
rect 55355 32861 55367 32895
rect 55309 32855 55367 32861
rect 55576 32895 55634 32901
rect 55576 32861 55588 32895
rect 55622 32892 55634 32895
rect 55950 32892 55956 32904
rect 55622 32864 55956 32892
rect 55622 32861 55634 32864
rect 55576 32855 55634 32861
rect 55950 32852 55956 32864
rect 56008 32852 56014 32904
rect 59449 32895 59507 32901
rect 59449 32892 59461 32895
rect 56888 32864 59461 32892
rect 45020 32796 46428 32824
rect 42398 32787 42456 32793
rect 16206 32756 16212 32768
rect 16167 32728 16212 32756
rect 16206 32716 16212 32728
rect 16264 32716 16270 32768
rect 18046 32756 18052 32768
rect 18007 32728 18052 32756
rect 18046 32716 18052 32728
rect 18104 32716 18110 32768
rect 28350 32756 28356 32768
rect 28311 32728 28356 32756
rect 28350 32716 28356 32728
rect 28408 32716 28414 32768
rect 31294 32756 31300 32768
rect 31255 32728 31300 32756
rect 31294 32716 31300 32728
rect 31352 32716 31358 32768
rect 33318 32756 33324 32768
rect 33279 32728 33324 32756
rect 33318 32716 33324 32728
rect 33376 32716 33382 32768
rect 36446 32716 36452 32768
rect 36504 32756 36510 32768
rect 38013 32759 38071 32765
rect 38013 32756 38025 32759
rect 36504 32728 38025 32756
rect 36504 32716 36510 32728
rect 38013 32725 38025 32728
rect 38059 32725 38071 32759
rect 41690 32756 41696 32768
rect 41651 32728 41696 32756
rect 38013 32719 38071 32725
rect 41690 32716 41696 32728
rect 41748 32716 41754 32768
rect 43530 32756 43536 32768
rect 43491 32728 43536 32756
rect 43530 32716 43536 32728
rect 43588 32716 43594 32768
rect 45526 32756 45554 32796
rect 46474 32784 46480 32836
rect 46532 32824 46538 32836
rect 47090 32827 47148 32833
rect 47090 32824 47102 32827
rect 46532 32796 47102 32824
rect 46532 32784 46538 32796
rect 47090 32793 47102 32796
rect 47136 32793 47148 32827
rect 47090 32787 47148 32793
rect 53644 32827 53702 32833
rect 53644 32793 53656 32827
rect 53690 32824 53702 32827
rect 56888 32824 56916 32864
rect 59449 32861 59461 32864
rect 59495 32861 59507 32895
rect 59449 32855 59507 32861
rect 57422 32833 57428 32836
rect 53690 32796 56916 32824
rect 53690 32793 53702 32796
rect 53644 32787 53702 32793
rect 57416 32787 57428 32833
rect 57480 32824 57486 32836
rect 57480 32796 57516 32824
rect 57422 32784 57428 32787
rect 57480 32784 57486 32796
rect 45646 32756 45652 32768
rect 45526 32728 45652 32756
rect 45646 32716 45652 32728
rect 45704 32716 45710 32768
rect 48222 32756 48228 32768
rect 48183 32728 48228 32756
rect 48222 32716 48228 32728
rect 48280 32716 48286 32768
rect 52362 32716 52368 32768
rect 52420 32756 52426 32768
rect 54757 32759 54815 32765
rect 54757 32756 54769 32759
rect 52420 32728 54769 32756
rect 52420 32716 52426 32728
rect 54757 32725 54769 32728
rect 54803 32725 54815 32759
rect 54757 32719 54815 32725
rect 1104 32666 59340 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 59340 32666
rect 1104 32592 59340 32614
rect 4706 32552 4712 32564
rect 4667 32524 4712 32552
rect 4706 32512 4712 32524
rect 4764 32512 4770 32564
rect 7745 32555 7803 32561
rect 7745 32521 7757 32555
rect 7791 32552 7803 32555
rect 8570 32552 8576 32564
rect 7791 32524 8576 32552
rect 7791 32521 7803 32524
rect 7745 32515 7803 32521
rect 8570 32512 8576 32524
rect 8628 32512 8634 32564
rect 9582 32552 9588 32564
rect 9543 32524 9588 32552
rect 9582 32512 9588 32524
rect 9640 32512 9646 32564
rect 18874 32512 18880 32564
rect 18932 32552 18938 32564
rect 19889 32555 19947 32561
rect 19889 32552 19901 32555
rect 18932 32524 19901 32552
rect 18932 32512 18938 32524
rect 19889 32521 19901 32524
rect 19935 32521 19947 32555
rect 19889 32515 19947 32521
rect 23842 32512 23848 32564
rect 23900 32552 23906 32564
rect 23937 32555 23995 32561
rect 23937 32552 23949 32555
rect 23900 32524 23949 32552
rect 23900 32512 23906 32524
rect 23937 32521 23949 32524
rect 23983 32521 23995 32555
rect 23937 32515 23995 32521
rect 25682 32512 25688 32564
rect 25740 32552 25746 32564
rect 25777 32555 25835 32561
rect 25777 32552 25789 32555
rect 25740 32524 25789 32552
rect 25740 32512 25746 32524
rect 25777 32521 25789 32524
rect 25823 32521 25835 32555
rect 25777 32515 25835 32521
rect 31481 32555 31539 32561
rect 31481 32521 31493 32555
rect 31527 32552 31539 32555
rect 31754 32552 31760 32564
rect 31527 32524 31760 32552
rect 31527 32521 31539 32524
rect 31481 32515 31539 32521
rect 31754 32512 31760 32524
rect 31812 32512 31818 32564
rect 38654 32552 38660 32564
rect 38615 32524 38660 32552
rect 38654 32512 38660 32524
rect 38712 32512 38718 32564
rect 43806 32552 43812 32564
rect 43767 32524 43812 32552
rect 43806 32512 43812 32524
rect 43864 32512 43870 32564
rect 45554 32512 45560 32564
rect 45612 32552 45618 32564
rect 45649 32555 45707 32561
rect 45649 32552 45661 32555
rect 45612 32524 45661 32552
rect 45612 32512 45618 32524
rect 45649 32521 45661 32524
rect 45695 32521 45707 32555
rect 45649 32515 45707 32521
rect 48866 32512 48872 32564
rect 48924 32552 48930 32564
rect 48961 32555 49019 32561
rect 48961 32552 48973 32555
rect 48924 32524 48973 32552
rect 48924 32512 48930 32524
rect 48961 32521 48973 32524
rect 49007 32521 49019 32555
rect 48961 32515 49019 32521
rect 57333 32555 57391 32561
rect 57333 32521 57345 32555
rect 57379 32552 57391 32555
rect 57422 32552 57428 32564
rect 57379 32524 57428 32552
rect 57379 32521 57391 32524
rect 57333 32515 57391 32521
rect 57422 32512 57428 32524
rect 57480 32512 57486 32564
rect 6632 32487 6690 32493
rect 6632 32453 6644 32487
rect 6678 32484 6690 32487
rect 8110 32484 8116 32496
rect 6678 32456 8116 32484
rect 6678 32453 6690 32456
rect 6632 32447 6690 32453
rect 8110 32444 8116 32456
rect 8168 32444 8174 32496
rect 8294 32444 8300 32496
rect 8352 32484 8358 32496
rect 12526 32493 12532 32496
rect 8450 32487 8508 32493
rect 8450 32484 8462 32487
rect 8352 32456 8462 32484
rect 8352 32444 8358 32456
rect 8450 32453 8462 32456
rect 8496 32453 8508 32487
rect 12520 32484 12532 32493
rect 12487 32456 12532 32484
rect 8450 32447 8508 32453
rect 12520 32447 12532 32456
rect 12526 32444 12532 32447
rect 12584 32444 12590 32496
rect 18046 32444 18052 32496
rect 18104 32484 18110 32496
rect 18754 32487 18812 32493
rect 18754 32484 18766 32487
rect 18104 32456 18766 32484
rect 18104 32444 18110 32456
rect 18754 32453 18766 32456
rect 18800 32453 18812 32487
rect 18754 32447 18812 32453
rect 22462 32444 22468 32496
rect 22520 32484 22526 32496
rect 22802 32487 22860 32493
rect 22802 32484 22814 32487
rect 22520 32456 22814 32484
rect 22520 32444 22526 32456
rect 22802 32453 22814 32456
rect 22848 32453 22860 32487
rect 22802 32447 22860 32453
rect 30368 32487 30426 32493
rect 30368 32453 30380 32487
rect 30414 32484 30426 32487
rect 31294 32484 31300 32496
rect 30414 32456 31300 32484
rect 30414 32453 30426 32456
rect 30368 32447 30426 32453
rect 31294 32444 31300 32456
rect 31352 32444 31358 32496
rect 32392 32487 32450 32493
rect 32392 32453 32404 32487
rect 32438 32484 32450 32487
rect 33318 32484 33324 32496
rect 32438 32456 33324 32484
rect 32438 32453 32450 32456
rect 32392 32447 32450 32453
rect 33318 32444 33324 32456
rect 33376 32444 33382 32496
rect 37918 32444 37924 32496
rect 37976 32484 37982 32496
rect 40120 32487 40178 32493
rect 37976 32456 39896 32484
rect 37976 32444 37982 32456
rect 3326 32416 3332 32428
rect 3287 32388 3332 32416
rect 3326 32376 3332 32388
rect 3384 32376 3390 32428
rect 3596 32419 3654 32425
rect 3596 32385 3608 32419
rect 3642 32416 3654 32419
rect 5166 32416 5172 32428
rect 3642 32388 5172 32416
rect 3642 32385 3654 32388
rect 3596 32379 3654 32385
rect 5166 32376 5172 32388
rect 5224 32376 5230 32428
rect 6365 32419 6423 32425
rect 6365 32385 6377 32419
rect 6411 32416 6423 32419
rect 6914 32416 6920 32428
rect 6411 32388 6920 32416
rect 6411 32385 6423 32388
rect 6365 32379 6423 32385
rect 6914 32376 6920 32388
rect 6972 32416 6978 32428
rect 8205 32419 8263 32425
rect 8205 32416 8217 32419
rect 6972 32388 8217 32416
rect 6972 32376 6978 32388
rect 8205 32385 8217 32388
rect 8251 32385 8263 32419
rect 13078 32416 13084 32428
rect 8205 32379 8263 32385
rect 12268 32388 13084 32416
rect 12066 32308 12072 32360
rect 12124 32348 12130 32360
rect 12268 32357 12296 32388
rect 13078 32376 13084 32388
rect 13136 32416 13142 32428
rect 13136 32388 13308 32416
rect 13136 32376 13142 32388
rect 12253 32351 12311 32357
rect 12253 32348 12265 32351
rect 12124 32320 12265 32348
rect 12124 32308 12130 32320
rect 12253 32317 12265 32320
rect 12299 32317 12311 32351
rect 13280 32348 13308 32388
rect 13814 32376 13820 32428
rect 13872 32416 13878 32428
rect 14349 32419 14407 32425
rect 14349 32416 14361 32419
rect 13872 32388 14361 32416
rect 13872 32376 13878 32388
rect 14349 32385 14361 32388
rect 14395 32385 14407 32419
rect 16666 32416 16672 32428
rect 16627 32388 16672 32416
rect 14349 32379 14407 32385
rect 16666 32376 16672 32388
rect 16724 32376 16730 32428
rect 16936 32419 16994 32425
rect 16936 32385 16948 32419
rect 16982 32416 16994 32419
rect 17310 32416 17316 32428
rect 16982 32388 17316 32416
rect 16982 32385 16994 32388
rect 16936 32379 16994 32385
rect 17310 32376 17316 32388
rect 17368 32376 17374 32428
rect 18509 32419 18567 32425
rect 18509 32385 18521 32419
rect 18555 32416 18567 32419
rect 19242 32416 19248 32428
rect 18555 32388 19248 32416
rect 18555 32385 18567 32388
rect 18509 32379 18567 32385
rect 19242 32376 19248 32388
rect 19300 32376 19306 32428
rect 21818 32376 21824 32428
rect 21876 32416 21882 32428
rect 22557 32419 22615 32425
rect 22557 32416 22569 32419
rect 21876 32388 22569 32416
rect 21876 32376 21882 32388
rect 22557 32385 22569 32388
rect 22603 32416 22615 32419
rect 24397 32419 24455 32425
rect 24397 32416 24409 32419
rect 22603 32388 24409 32416
rect 22603 32385 22615 32388
rect 22557 32379 22615 32385
rect 24397 32385 24409 32388
rect 24443 32385 24455 32419
rect 24397 32379 24455 32385
rect 24486 32376 24492 32428
rect 24544 32416 24550 32428
rect 24653 32419 24711 32425
rect 24653 32416 24665 32419
rect 24544 32388 24665 32416
rect 24544 32376 24550 32388
rect 24653 32385 24665 32388
rect 24699 32385 24711 32419
rect 24653 32379 24711 32385
rect 28160 32419 28218 32425
rect 28160 32385 28172 32419
rect 28206 32416 28218 32419
rect 29086 32416 29092 32428
rect 28206 32388 29092 32416
rect 28206 32385 28218 32388
rect 28160 32379 28218 32385
rect 29086 32376 29092 32388
rect 29144 32376 29150 32428
rect 29914 32376 29920 32428
rect 29972 32416 29978 32428
rect 30101 32419 30159 32425
rect 30101 32416 30113 32419
rect 29972 32388 30113 32416
rect 29972 32376 29978 32388
rect 30101 32385 30113 32388
rect 30147 32385 30159 32419
rect 30101 32379 30159 32385
rect 31662 32376 31668 32428
rect 31720 32416 31726 32428
rect 32125 32419 32183 32425
rect 32125 32416 32137 32419
rect 31720 32388 32137 32416
rect 31720 32376 31726 32388
rect 32125 32385 32137 32388
rect 32171 32385 32183 32419
rect 32125 32379 32183 32385
rect 34609 32419 34667 32425
rect 34609 32385 34621 32419
rect 34655 32416 34667 32419
rect 34698 32416 34704 32428
rect 34655 32388 34704 32416
rect 34655 32385 34667 32388
rect 34609 32379 34667 32385
rect 34698 32376 34704 32388
rect 34756 32376 34762 32428
rect 34876 32419 34934 32425
rect 34876 32385 34888 32419
rect 34922 32416 34934 32419
rect 36354 32416 36360 32428
rect 34922 32388 36360 32416
rect 34922 32385 34934 32388
rect 34876 32379 34934 32385
rect 36354 32376 36360 32388
rect 36412 32376 36418 32428
rect 37544 32419 37602 32425
rect 37544 32385 37556 32419
rect 37590 32416 37602 32419
rect 39298 32416 39304 32428
rect 37590 32388 39304 32416
rect 37590 32385 37602 32388
rect 37544 32379 37602 32385
rect 39298 32376 39304 32388
rect 39356 32376 39362 32428
rect 39868 32425 39896 32456
rect 40120 32453 40132 32487
rect 40166 32484 40178 32487
rect 41690 32484 41696 32496
rect 40166 32456 41696 32484
rect 40166 32453 40178 32456
rect 40120 32447 40178 32453
rect 41690 32444 41696 32456
rect 41748 32444 41754 32496
rect 44174 32484 44180 32496
rect 42444 32456 44180 32484
rect 39853 32419 39911 32425
rect 39853 32385 39865 32419
rect 39899 32416 39911 32419
rect 40402 32416 40408 32428
rect 39899 32388 40408 32416
rect 39899 32385 39911 32388
rect 39853 32379 39911 32385
rect 40402 32376 40408 32388
rect 40460 32376 40466 32428
rect 42150 32376 42156 32428
rect 42208 32416 42214 32428
rect 42444 32425 42472 32456
rect 44174 32444 44180 32456
rect 44232 32484 44238 32496
rect 44536 32487 44594 32493
rect 44232 32456 44312 32484
rect 44232 32444 44238 32456
rect 42429 32419 42487 32425
rect 42429 32416 42441 32419
rect 42208 32388 42441 32416
rect 42208 32376 42214 32388
rect 42429 32385 42441 32388
rect 42475 32385 42487 32419
rect 42429 32379 42487 32385
rect 42696 32419 42754 32425
rect 42696 32385 42708 32419
rect 42742 32416 42754 32419
rect 43622 32416 43628 32428
rect 42742 32388 43628 32416
rect 42742 32385 42754 32388
rect 42696 32379 42754 32385
rect 43622 32376 43628 32388
rect 43680 32376 43686 32428
rect 44284 32425 44312 32456
rect 44536 32453 44548 32487
rect 44582 32484 44594 32487
rect 45002 32484 45008 32496
rect 44582 32456 45008 32484
rect 44582 32453 44594 32456
rect 44536 32447 44594 32453
rect 45002 32444 45008 32456
rect 45060 32444 45066 32496
rect 47848 32487 47906 32493
rect 47848 32453 47860 32487
rect 47894 32484 47906 32487
rect 48222 32484 48228 32496
rect 47894 32456 48228 32484
rect 47894 32453 47906 32456
rect 47848 32447 47906 32453
rect 48222 32444 48228 32456
rect 48280 32444 48286 32496
rect 54380 32487 54438 32493
rect 54380 32453 54392 32487
rect 54426 32484 54438 32487
rect 58526 32484 58532 32496
rect 54426 32456 58532 32484
rect 54426 32453 54438 32456
rect 54380 32447 54438 32453
rect 58526 32444 58532 32456
rect 58584 32444 58590 32496
rect 44269 32419 44327 32425
rect 44269 32385 44281 32419
rect 44315 32385 44327 32419
rect 47578 32416 47584 32428
rect 47539 32388 47584 32416
rect 44269 32379 44327 32385
rect 47578 32376 47584 32388
rect 47636 32376 47642 32428
rect 51068 32419 51126 32425
rect 51068 32385 51080 32419
rect 51114 32416 51126 32419
rect 52270 32416 52276 32428
rect 51114 32388 52276 32416
rect 51114 32385 51126 32388
rect 51068 32379 51126 32385
rect 52270 32376 52276 32388
rect 52328 32376 52334 32428
rect 52730 32376 52736 32428
rect 52788 32416 52794 32428
rect 54113 32419 54171 32425
rect 54113 32416 54125 32419
rect 52788 32388 54125 32416
rect 52788 32376 52794 32388
rect 54113 32385 54125 32388
rect 54159 32416 54171 32419
rect 55953 32419 56011 32425
rect 55953 32416 55965 32419
rect 54159 32388 55965 32416
rect 54159 32385 54171 32388
rect 54113 32379 54171 32385
rect 55953 32385 55965 32388
rect 55999 32385 56011 32419
rect 55953 32379 56011 32385
rect 56220 32419 56278 32425
rect 56220 32385 56232 32419
rect 56266 32416 56278 32419
rect 57882 32416 57888 32428
rect 56266 32388 57888 32416
rect 56266 32385 56278 32388
rect 56220 32379 56278 32385
rect 57882 32376 57888 32388
rect 57940 32376 57946 32428
rect 14093 32351 14151 32357
rect 14093 32348 14105 32351
rect 13280 32320 14105 32348
rect 12253 32311 12311 32317
rect 14093 32317 14105 32320
rect 14139 32317 14151 32351
rect 14093 32311 14151 32317
rect 27522 32308 27528 32360
rect 27580 32348 27586 32360
rect 27893 32351 27951 32357
rect 27893 32348 27905 32351
rect 27580 32320 27905 32348
rect 27580 32308 27586 32320
rect 27893 32317 27905 32320
rect 27939 32317 27951 32351
rect 27893 32311 27951 32317
rect 35894 32308 35900 32360
rect 35952 32348 35958 32360
rect 37274 32348 37280 32360
rect 35952 32320 37280 32348
rect 35952 32308 35958 32320
rect 37274 32308 37280 32320
rect 37332 32308 37338 32360
rect 50798 32348 50804 32360
rect 50759 32320 50804 32348
rect 50798 32308 50804 32320
rect 50856 32308 50862 32360
rect 17954 32240 17960 32292
rect 18012 32280 18018 32292
rect 18049 32283 18107 32289
rect 18049 32280 18061 32283
rect 18012 32252 18061 32280
rect 18012 32240 18018 32252
rect 18049 32249 18061 32252
rect 18095 32249 18107 32283
rect 18049 32243 18107 32249
rect 10502 32172 10508 32224
rect 10560 32212 10566 32224
rect 13633 32215 13691 32221
rect 13633 32212 13645 32215
rect 10560 32184 13645 32212
rect 10560 32172 10566 32184
rect 13633 32181 13645 32184
rect 13679 32181 13691 32215
rect 13633 32175 13691 32181
rect 13906 32172 13912 32224
rect 13964 32212 13970 32224
rect 15473 32215 15531 32221
rect 15473 32212 15485 32215
rect 13964 32184 15485 32212
rect 13964 32172 13970 32184
rect 15473 32181 15485 32184
rect 15519 32181 15531 32215
rect 29270 32212 29276 32224
rect 29231 32184 29276 32212
rect 15473 32175 15531 32181
rect 29270 32172 29276 32184
rect 29328 32172 29334 32224
rect 33502 32212 33508 32224
rect 33463 32184 33508 32212
rect 33502 32172 33508 32184
rect 33560 32172 33566 32224
rect 35986 32212 35992 32224
rect 35947 32184 35992 32212
rect 35986 32172 35992 32184
rect 36044 32172 36050 32224
rect 41230 32212 41236 32224
rect 41191 32184 41236 32212
rect 41230 32172 41236 32184
rect 41288 32172 41294 32224
rect 51074 32172 51080 32224
rect 51132 32212 51138 32224
rect 52181 32215 52239 32221
rect 52181 32212 52193 32215
rect 51132 32184 52193 32212
rect 51132 32172 51138 32184
rect 52181 32181 52193 32184
rect 52227 32181 52239 32215
rect 55490 32212 55496 32224
rect 55451 32184 55496 32212
rect 52181 32175 52239 32181
rect 55490 32172 55496 32184
rect 55548 32172 55554 32224
rect 1104 32122 59340 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 59340 32122
rect 1104 32048 59340 32070
rect 4982 32008 4988 32020
rect 3804 31980 4988 32008
rect 2866 31764 2872 31816
rect 2924 31804 2930 31816
rect 3804 31813 3832 31980
rect 4982 31968 4988 31980
rect 5040 31968 5046 32020
rect 5166 32008 5172 32020
rect 5127 31980 5172 32008
rect 5166 31968 5172 31980
rect 5224 31968 5230 32020
rect 16574 31968 16580 32020
rect 16632 32008 16638 32020
rect 17313 32011 17371 32017
rect 17313 32008 17325 32011
rect 16632 31980 17325 32008
rect 16632 31968 16638 31980
rect 17313 31977 17325 31980
rect 17359 31977 17371 32011
rect 27522 32008 27528 32020
rect 27483 31980 27528 32008
rect 17313 31971 17371 31977
rect 27522 31968 27528 31980
rect 27580 31968 27586 32020
rect 33505 32011 33563 32017
rect 33505 31977 33517 32011
rect 33551 32008 33563 32011
rect 33870 32008 33876 32020
rect 33551 31980 33876 32008
rect 33551 31977 33563 31980
rect 33505 31971 33563 31977
rect 33870 31968 33876 31980
rect 33928 31968 33934 32020
rect 39298 32008 39304 32020
rect 39259 31980 39304 32008
rect 39298 31968 39304 31980
rect 39356 31968 39362 32020
rect 41782 32008 41788 32020
rect 41743 31980 41788 32008
rect 41782 31968 41788 31980
rect 41840 31968 41846 32020
rect 43622 32008 43628 32020
rect 43583 31980 43628 32008
rect 43622 31968 43628 31980
rect 43680 31968 43686 32020
rect 46385 32011 46443 32017
rect 46385 31977 46397 32011
rect 46431 32008 46443 32011
rect 46474 32008 46480 32020
rect 46431 31980 46480 32008
rect 46431 31977 46443 31980
rect 46385 31971 46443 31977
rect 46474 31968 46480 31980
rect 46532 31968 46538 32020
rect 50798 32008 50804 32020
rect 48240 31980 50804 32008
rect 11609 31943 11667 31949
rect 11609 31909 11621 31943
rect 11655 31909 11667 31943
rect 11609 31903 11667 31909
rect 10226 31872 10232 31884
rect 10187 31844 10232 31872
rect 10226 31832 10232 31844
rect 10284 31832 10290 31884
rect 11624 31872 11652 31903
rect 31202 31900 31208 31952
rect 31260 31940 31266 31952
rect 31573 31943 31631 31949
rect 31573 31940 31585 31943
rect 31260 31912 31585 31940
rect 31260 31900 31266 31912
rect 31573 31909 31585 31912
rect 31619 31909 31631 31943
rect 31573 31903 31631 31909
rect 11624 31844 12204 31872
rect 3789 31807 3847 31813
rect 3789 31804 3801 31807
rect 2924 31776 3801 31804
rect 2924 31764 2930 31776
rect 3789 31773 3801 31776
rect 3835 31773 3847 31807
rect 3789 31767 3847 31773
rect 4056 31807 4114 31813
rect 4056 31773 4068 31807
rect 4102 31804 4114 31807
rect 10244 31804 10272 31832
rect 10502 31813 10508 31816
rect 10496 31804 10508 31813
rect 4102 31776 4200 31804
rect 10244 31776 10364 31804
rect 10463 31776 10508 31804
rect 4102 31773 4114 31776
rect 4056 31767 4114 31773
rect 4172 31736 4200 31776
rect 4246 31736 4252 31748
rect 4172 31708 4252 31736
rect 4246 31696 4252 31708
rect 4304 31696 4310 31748
rect 10336 31736 10364 31776
rect 10496 31767 10508 31776
rect 10502 31764 10508 31767
rect 10560 31764 10566 31816
rect 11514 31804 11520 31816
rect 10612 31776 11520 31804
rect 10612 31736 10640 31776
rect 11514 31764 11520 31776
rect 11572 31804 11578 31816
rect 12066 31804 12072 31816
rect 11572 31776 12072 31804
rect 11572 31764 11578 31776
rect 12066 31764 12072 31776
rect 12124 31764 12130 31816
rect 12176 31804 12204 31844
rect 13078 31832 13084 31884
rect 13136 31872 13142 31884
rect 14093 31875 14151 31881
rect 14093 31872 14105 31875
rect 13136 31844 14105 31872
rect 13136 31832 13142 31844
rect 14093 31841 14105 31844
rect 14139 31841 14151 31875
rect 14093 31835 14151 31841
rect 19242 31832 19248 31884
rect 19300 31872 19306 31884
rect 19613 31875 19671 31881
rect 19613 31872 19625 31875
rect 19300 31844 19625 31872
rect 19300 31832 19306 31844
rect 19613 31841 19625 31844
rect 19659 31841 19671 31875
rect 19613 31835 19671 31841
rect 35894 31832 35900 31884
rect 35952 31872 35958 31884
rect 35952 31844 35997 31872
rect 35952 31832 35958 31844
rect 37274 31832 37280 31884
rect 37332 31872 37338 31884
rect 37918 31872 37924 31884
rect 37332 31844 37924 31872
rect 37332 31832 37338 31844
rect 37918 31832 37924 31844
rect 37976 31832 37982 31884
rect 40402 31872 40408 31884
rect 40363 31844 40408 31872
rect 40402 31832 40408 31844
rect 40460 31832 40466 31884
rect 42150 31832 42156 31884
rect 42208 31872 42214 31884
rect 42245 31875 42303 31881
rect 42245 31872 42257 31875
rect 42208 31844 42257 31872
rect 42208 31832 42214 31844
rect 42245 31841 42257 31844
rect 42291 31841 42303 31875
rect 42245 31835 42303 31841
rect 44910 31832 44916 31884
rect 44968 31872 44974 31884
rect 48240 31881 48268 31980
rect 50798 31968 50804 31980
rect 50856 31968 50862 32020
rect 54757 32011 54815 32017
rect 54757 31977 54769 32011
rect 54803 32008 54815 32011
rect 56870 32008 56876 32020
rect 54803 31980 56876 32008
rect 54803 31977 54815 31980
rect 54757 31971 54815 31977
rect 56870 31968 56876 31980
rect 56928 31968 56934 32020
rect 57882 32008 57888 32020
rect 57843 31980 57888 32008
rect 57882 31968 57888 31980
rect 57940 31968 57946 32020
rect 45005 31875 45063 31881
rect 45005 31872 45017 31875
rect 44968 31844 45017 31872
rect 44968 31832 44974 31844
rect 45005 31841 45017 31844
rect 45051 31841 45063 31875
rect 45005 31835 45063 31841
rect 48225 31875 48283 31881
rect 48225 31841 48237 31875
rect 48271 31841 48283 31875
rect 48225 31835 48283 31841
rect 50798 31832 50804 31884
rect 50856 31872 50862 31884
rect 51537 31875 51595 31881
rect 51537 31872 51549 31875
rect 50856 31844 51549 31872
rect 50856 31832 50862 31844
rect 51537 31841 51549 31844
rect 51583 31841 51595 31875
rect 51537 31835 51595 31841
rect 52730 31832 52736 31884
rect 52788 31872 52794 31884
rect 53377 31875 53435 31881
rect 53377 31872 53389 31875
rect 52788 31844 53389 31872
rect 52788 31832 52794 31844
rect 53377 31841 53389 31844
rect 53423 31841 53435 31875
rect 53377 31835 53435 31841
rect 12325 31807 12383 31813
rect 12325 31804 12337 31807
rect 12176 31776 12337 31804
rect 12325 31773 12337 31776
rect 12371 31773 12383 31807
rect 12325 31767 12383 31773
rect 14360 31807 14418 31813
rect 14360 31773 14372 31807
rect 14406 31804 14418 31807
rect 15470 31804 15476 31816
rect 14406 31776 15476 31804
rect 14406 31773 14418 31776
rect 14360 31767 14418 31773
rect 15470 31764 15476 31776
rect 15528 31764 15534 31816
rect 15933 31807 15991 31813
rect 15933 31773 15945 31807
rect 15979 31804 15991 31807
rect 16666 31804 16672 31816
rect 15979 31776 16672 31804
rect 15979 31773 15991 31776
rect 15933 31767 15991 31773
rect 16666 31764 16672 31776
rect 16724 31764 16730 31816
rect 19880 31807 19938 31813
rect 19880 31773 19892 31807
rect 19926 31804 19938 31807
rect 21266 31804 21272 31816
rect 19926 31776 21272 31804
rect 19926 31773 19938 31776
rect 19880 31767 19938 31773
rect 21266 31764 21272 31776
rect 21324 31764 21330 31816
rect 22373 31807 22431 31813
rect 22373 31773 22385 31807
rect 22419 31804 22431 31807
rect 22462 31804 22468 31816
rect 22419 31776 22468 31804
rect 22419 31773 22431 31776
rect 22373 31767 22431 31773
rect 22462 31764 22468 31776
rect 22520 31764 22526 31816
rect 22640 31807 22698 31813
rect 22640 31773 22652 31807
rect 22686 31804 22698 31807
rect 23658 31804 23664 31816
rect 22686 31776 23664 31804
rect 22686 31773 22698 31776
rect 22640 31767 22698 31773
rect 23658 31764 23664 31776
rect 23716 31764 23722 31816
rect 24854 31764 24860 31816
rect 24912 31804 24918 31816
rect 26053 31807 26111 31813
rect 26053 31804 26065 31807
rect 24912 31776 26065 31804
rect 24912 31764 24918 31776
rect 26053 31773 26065 31776
rect 26099 31773 26111 31807
rect 26053 31767 26111 31773
rect 30193 31807 30251 31813
rect 30193 31773 30205 31807
rect 30239 31804 30251 31807
rect 30460 31807 30518 31813
rect 30239 31776 30420 31804
rect 30239 31773 30251 31776
rect 30193 31767 30251 31773
rect 10336 31708 10640 31736
rect 15562 31696 15568 31748
rect 15620 31736 15626 31748
rect 16178 31739 16236 31745
rect 16178 31736 16190 31739
rect 15620 31708 16190 31736
rect 15620 31696 15626 31708
rect 16178 31705 16190 31708
rect 16224 31705 16236 31739
rect 30392 31736 30420 31776
rect 30460 31773 30472 31807
rect 30506 31804 30518 31807
rect 31478 31804 31484 31816
rect 30506 31776 31484 31804
rect 30506 31773 30518 31776
rect 30460 31767 30518 31773
rect 31478 31764 31484 31776
rect 31536 31764 31542 31816
rect 32122 31804 32128 31816
rect 32083 31776 32128 31804
rect 32122 31764 32128 31776
rect 32180 31764 32186 31816
rect 32392 31807 32450 31813
rect 32392 31773 32404 31807
rect 32438 31804 32450 31807
rect 33502 31804 33508 31816
rect 32438 31776 33508 31804
rect 32438 31773 32450 31776
rect 32392 31767 32450 31773
rect 33502 31764 33508 31776
rect 33560 31764 33566 31816
rect 36164 31807 36222 31813
rect 36164 31773 36176 31807
rect 36210 31804 36222 31807
rect 36446 31804 36452 31816
rect 36210 31776 36452 31804
rect 36210 31773 36222 31776
rect 36164 31767 36222 31773
rect 36446 31764 36452 31776
rect 36504 31764 36510 31816
rect 38188 31807 38246 31813
rect 38188 31773 38200 31807
rect 38234 31804 38246 31807
rect 39298 31804 39304 31816
rect 38234 31776 39304 31804
rect 38234 31773 38246 31776
rect 38188 31767 38246 31773
rect 39298 31764 39304 31776
rect 39356 31764 39362 31816
rect 40672 31807 40730 31813
rect 40672 31773 40684 31807
rect 40718 31804 40730 31807
rect 41230 31804 41236 31816
rect 40718 31776 41236 31804
rect 40718 31773 40730 31776
rect 40672 31767 40730 31773
rect 41230 31764 41236 31776
rect 41288 31764 41294 31816
rect 42512 31807 42570 31813
rect 42512 31773 42524 31807
rect 42558 31804 42570 31807
rect 43530 31804 43536 31816
rect 42558 31776 43536 31804
rect 42558 31773 42570 31776
rect 42512 31767 42570 31773
rect 43530 31764 43536 31776
rect 43588 31764 43594 31816
rect 45272 31807 45330 31813
rect 45272 31773 45284 31807
rect 45318 31804 45330 31807
rect 46382 31804 46388 31816
rect 45318 31776 46388 31804
rect 45318 31773 45330 31776
rect 45272 31767 45330 31773
rect 46382 31764 46388 31776
rect 46440 31764 46446 31816
rect 48492 31807 48550 31813
rect 48492 31773 48504 31807
rect 48538 31804 48550 31807
rect 50154 31804 50160 31816
rect 48538 31776 50160 31804
rect 48538 31773 48550 31776
rect 48492 31767 48550 31773
rect 50154 31764 50160 31776
rect 50212 31764 50218 31816
rect 51804 31807 51862 31813
rect 51804 31773 51816 31807
rect 51850 31804 51862 31807
rect 52362 31804 52368 31816
rect 51850 31776 52368 31804
rect 51850 31773 51862 31776
rect 51804 31767 51862 31773
rect 52362 31764 52368 31776
rect 52420 31764 52426 31816
rect 53644 31807 53702 31813
rect 53644 31773 53656 31807
rect 53690 31804 53702 31807
rect 55490 31804 55496 31816
rect 53690 31776 55496 31804
rect 53690 31773 53702 31776
rect 53644 31767 53702 31773
rect 55490 31764 55496 31776
rect 55548 31764 55554 31816
rect 56505 31807 56563 31813
rect 56505 31773 56517 31807
rect 56551 31804 56563 31807
rect 56772 31807 56830 31813
rect 56551 31776 56640 31804
rect 56551 31773 56563 31776
rect 56505 31767 56563 31773
rect 32140 31736 32168 31764
rect 30392 31708 32168 31736
rect 56612 31736 56640 31776
rect 56772 31773 56784 31807
rect 56818 31804 56830 31807
rect 58526 31804 58532 31816
rect 56818 31776 58532 31804
rect 56818 31773 56830 31776
rect 56772 31767 56830 31773
rect 58526 31764 58532 31776
rect 58584 31764 58590 31816
rect 57054 31736 57060 31748
rect 56612 31708 57060 31736
rect 16178 31699 16236 31705
rect 57054 31696 57060 31708
rect 57112 31696 57118 31748
rect 13446 31668 13452 31680
rect 13407 31640 13452 31668
rect 13446 31628 13452 31640
rect 13504 31628 13510 31680
rect 15470 31668 15476 31680
rect 15431 31640 15476 31668
rect 15470 31628 15476 31640
rect 15528 31628 15534 31680
rect 20990 31668 20996 31680
rect 20951 31640 20996 31668
rect 20990 31628 20996 31640
rect 21048 31628 21054 31680
rect 23750 31668 23756 31680
rect 23711 31640 23756 31668
rect 23750 31628 23756 31640
rect 23808 31628 23814 31680
rect 37274 31668 37280 31680
rect 37235 31640 37280 31668
rect 37274 31628 37280 31640
rect 37332 31628 37338 31680
rect 49602 31668 49608 31680
rect 49563 31640 49608 31668
rect 49602 31628 49608 31640
rect 49660 31628 49666 31680
rect 52454 31628 52460 31680
rect 52512 31668 52518 31680
rect 52917 31671 52975 31677
rect 52917 31668 52929 31671
rect 52512 31640 52929 31668
rect 52512 31628 52518 31640
rect 52917 31637 52929 31640
rect 52963 31637 52975 31671
rect 52917 31631 52975 31637
rect 1104 31578 59340 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 59340 31578
rect 1104 31504 59340 31526
rect 4246 31464 4252 31476
rect 4207 31436 4252 31464
rect 4246 31424 4252 31436
rect 4304 31424 4310 31476
rect 14734 31464 14740 31476
rect 14695 31436 14740 31464
rect 14734 31424 14740 31436
rect 14792 31424 14798 31476
rect 21266 31464 21272 31476
rect 21227 31436 21272 31464
rect 21266 31424 21272 31436
rect 21324 31424 21330 31476
rect 30834 31424 30840 31476
rect 30892 31464 30898 31476
rect 31110 31464 31116 31476
rect 30892 31436 31116 31464
rect 30892 31424 30898 31436
rect 31110 31424 31116 31436
rect 31168 31464 31174 31476
rect 34606 31464 34612 31476
rect 31168 31436 34468 31464
rect 34567 31436 34612 31464
rect 31168 31424 31174 31436
rect 3694 31356 3700 31408
rect 3752 31396 3758 31408
rect 29825 31399 29883 31405
rect 29825 31396 29837 31399
rect 3752 31368 29837 31396
rect 3752 31356 3758 31368
rect 29825 31365 29837 31368
rect 29871 31365 29883 31399
rect 29825 31359 29883 31365
rect 33496 31399 33554 31405
rect 33496 31365 33508 31399
rect 33542 31396 33554 31399
rect 33594 31396 33600 31408
rect 33542 31368 33600 31396
rect 33542 31365 33554 31368
rect 33496 31359 33554 31365
rect 33594 31356 33600 31368
rect 33652 31356 33658 31408
rect 34440 31396 34468 31436
rect 34606 31424 34612 31436
rect 34664 31424 34670 31476
rect 36354 31424 36360 31476
rect 36412 31464 36418 31476
rect 36449 31467 36507 31473
rect 36449 31464 36461 31467
rect 36412 31436 36461 31464
rect 36412 31424 36418 31436
rect 36449 31433 36461 31436
rect 36495 31433 36507 31467
rect 43990 31464 43996 31476
rect 43951 31436 43996 31464
rect 36449 31427 36507 31433
rect 43990 31424 43996 31436
rect 44048 31424 44054 31476
rect 50341 31467 50399 31473
rect 50341 31433 50353 31467
rect 50387 31464 50399 31467
rect 51258 31464 51264 31476
rect 50387 31436 51264 31464
rect 50387 31433 50399 31436
rect 50341 31427 50399 31433
rect 51258 31424 51264 31436
rect 51316 31424 51322 31476
rect 52181 31467 52239 31473
rect 52181 31433 52193 31467
rect 52227 31433 52239 31467
rect 52181 31427 52239 31433
rect 35336 31399 35394 31405
rect 34440 31368 35195 31396
rect 2866 31328 2872 31340
rect 2827 31300 2872 31328
rect 2866 31288 2872 31300
rect 2924 31288 2930 31340
rect 3136 31331 3194 31337
rect 3136 31297 3148 31331
rect 3182 31328 3194 31331
rect 3970 31328 3976 31340
rect 3182 31300 3976 31328
rect 3182 31297 3194 31300
rect 3136 31291 3194 31297
rect 3970 31288 3976 31300
rect 4028 31288 4034 31340
rect 11514 31328 11520 31340
rect 11475 31300 11520 31328
rect 11514 31288 11520 31300
rect 11572 31288 11578 31340
rect 11784 31331 11842 31337
rect 11784 31297 11796 31331
rect 11830 31328 11842 31331
rect 13446 31328 13452 31340
rect 11830 31300 13452 31328
rect 11830 31297 11842 31300
rect 11784 31291 11842 31297
rect 13446 31288 13452 31300
rect 13504 31288 13510 31340
rect 13624 31331 13682 31337
rect 13624 31297 13636 31331
rect 13670 31328 13682 31331
rect 13906 31328 13912 31340
rect 13670 31300 13912 31328
rect 13670 31297 13682 31300
rect 13624 31291 13682 31297
rect 13906 31288 13912 31300
rect 13964 31288 13970 31340
rect 16666 31288 16672 31340
rect 16724 31328 16730 31340
rect 18049 31331 18107 31337
rect 18049 31328 18061 31331
rect 16724 31300 18061 31328
rect 16724 31288 16730 31300
rect 18049 31297 18061 31300
rect 18095 31297 18107 31331
rect 18049 31291 18107 31297
rect 18316 31331 18374 31337
rect 18316 31297 18328 31331
rect 18362 31328 18374 31331
rect 19334 31328 19340 31340
rect 18362 31300 19340 31328
rect 18362 31297 18374 31300
rect 18316 31291 18374 31297
rect 19334 31288 19340 31300
rect 19392 31288 19398 31340
rect 20156 31331 20214 31337
rect 20156 31297 20168 31331
rect 20202 31328 20214 31331
rect 21266 31328 21272 31340
rect 20202 31300 21272 31328
rect 20202 31297 20214 31300
rect 20156 31291 20214 31297
rect 21266 31288 21272 31300
rect 21324 31288 21330 31340
rect 22462 31288 22468 31340
rect 22520 31328 22526 31340
rect 23201 31331 23259 31337
rect 23201 31328 23213 31331
rect 22520 31300 23213 31328
rect 22520 31288 22526 31300
rect 23201 31297 23213 31300
rect 23247 31328 23259 31331
rect 23290 31328 23296 31340
rect 23247 31300 23296 31328
rect 23247 31297 23259 31300
rect 23201 31291 23259 31297
rect 23290 31288 23296 31300
rect 23348 31288 23354 31340
rect 23468 31331 23526 31337
rect 23468 31297 23480 31331
rect 23514 31328 23526 31331
rect 25308 31331 25366 31337
rect 23514 31300 24900 31328
rect 23514 31297 23526 31300
rect 23468 31291 23526 31297
rect 13078 31220 13084 31272
rect 13136 31260 13142 31272
rect 13357 31263 13415 31269
rect 13357 31260 13369 31263
rect 13136 31232 13369 31260
rect 13136 31220 13142 31232
rect 13357 31229 13369 31232
rect 13403 31229 13415 31263
rect 13357 31223 13415 31229
rect 19242 31220 19248 31272
rect 19300 31260 19306 31272
rect 19889 31263 19947 31269
rect 19889 31260 19901 31263
rect 19300 31232 19901 31260
rect 19300 31220 19306 31232
rect 19889 31229 19901 31232
rect 19935 31229 19947 31263
rect 19889 31223 19947 31229
rect 12894 31124 12900 31136
rect 12855 31096 12900 31124
rect 12894 31084 12900 31096
rect 12952 31084 12958 31136
rect 19426 31124 19432 31136
rect 19387 31096 19432 31124
rect 19426 31084 19432 31096
rect 19484 31084 19490 31136
rect 24578 31124 24584 31136
rect 24539 31096 24584 31124
rect 24578 31084 24584 31096
rect 24636 31084 24642 31136
rect 24872 31124 24900 31300
rect 25308 31297 25320 31331
rect 25354 31328 25366 31331
rect 27062 31328 27068 31340
rect 25354 31300 27068 31328
rect 25354 31297 25366 31300
rect 25308 31291 25366 31297
rect 27062 31288 27068 31300
rect 27120 31288 27126 31340
rect 28252 31331 28310 31337
rect 28252 31297 28264 31331
rect 28298 31328 28310 31331
rect 29730 31328 29736 31340
rect 28298 31300 29736 31328
rect 28298 31297 28310 31300
rect 28252 31291 28310 31297
rect 29730 31288 29736 31300
rect 29788 31288 29794 31340
rect 34698 31288 34704 31340
rect 34756 31328 34762 31340
rect 35069 31331 35127 31337
rect 35069 31328 35081 31331
rect 34756 31300 35081 31328
rect 34756 31288 34762 31300
rect 35069 31297 35081 31300
rect 35115 31297 35127 31331
rect 35167 31328 35195 31368
rect 35336 31365 35348 31399
rect 35382 31396 35394 31399
rect 37274 31396 37280 31408
rect 35382 31368 37280 31396
rect 35382 31365 35394 31368
rect 35336 31359 35394 31365
rect 37274 31356 37280 31368
rect 37332 31356 37338 31408
rect 40494 31396 40500 31408
rect 37844 31368 40500 31396
rect 37844 31328 37872 31368
rect 40494 31356 40500 31368
rect 40552 31356 40558 31408
rect 42880 31399 42938 31405
rect 42880 31365 42892 31399
rect 42926 31396 42938 31399
rect 44266 31396 44272 31408
rect 42926 31368 44272 31396
rect 42926 31365 42938 31368
rect 42880 31359 42938 31365
rect 44266 31356 44272 31368
rect 44324 31356 44330 31408
rect 49228 31399 49286 31405
rect 49228 31365 49240 31399
rect 49274 31396 49286 31399
rect 52196 31396 52224 31427
rect 49274 31368 52224 31396
rect 49274 31365 49286 31368
rect 49228 31359 49286 31365
rect 35167 31300 37872 31328
rect 35069 31291 35127 31297
rect 37918 31288 37924 31340
rect 37976 31328 37982 31340
rect 38289 31331 38347 31337
rect 38289 31328 38301 31331
rect 37976 31300 38301 31328
rect 37976 31288 37982 31300
rect 38289 31297 38301 31300
rect 38335 31297 38347 31331
rect 38289 31291 38347 31297
rect 38556 31331 38614 31337
rect 38556 31297 38568 31331
rect 38602 31328 38614 31331
rect 40586 31328 40592 31340
rect 38602 31300 40592 31328
rect 38602 31297 38614 31300
rect 38556 31291 38614 31297
rect 40586 31288 40592 31300
rect 40644 31288 40650 31340
rect 40764 31331 40822 31337
rect 40764 31297 40776 31331
rect 40810 31328 40822 31331
rect 42426 31328 42432 31340
rect 40810 31300 42432 31328
rect 40810 31297 40822 31300
rect 40764 31291 40822 31297
rect 42426 31288 42432 31300
rect 42484 31288 42490 31340
rect 42610 31328 42616 31340
rect 42571 31300 42616 31328
rect 42610 31288 42616 31300
rect 42668 31288 42674 31340
rect 45646 31328 45652 31340
rect 45607 31300 45652 31328
rect 45646 31288 45652 31300
rect 45704 31288 45710 31340
rect 45916 31331 45974 31337
rect 45916 31297 45928 31331
rect 45962 31328 45974 31331
rect 46934 31328 46940 31340
rect 45962 31300 46940 31328
rect 45962 31297 45974 31300
rect 45916 31291 45974 31297
rect 46934 31288 46940 31300
rect 46992 31288 46998 31340
rect 47578 31288 47584 31340
rect 47636 31328 47642 31340
rect 48961 31331 49019 31337
rect 48961 31328 48973 31331
rect 47636 31300 48973 31328
rect 47636 31288 47642 31300
rect 48961 31297 48973 31300
rect 49007 31297 49019 31331
rect 50798 31328 50804 31340
rect 50759 31300 50804 31328
rect 48961 31291 49019 31297
rect 50798 31288 50804 31300
rect 50856 31288 50862 31340
rect 51068 31331 51126 31337
rect 51068 31297 51080 31331
rect 51114 31328 51126 31331
rect 52178 31328 52184 31340
rect 51114 31300 52184 31328
rect 51114 31297 51126 31300
rect 51068 31291 51126 31297
rect 52178 31288 52184 31300
rect 52236 31288 52242 31340
rect 54472 31331 54530 31337
rect 54472 31297 54484 31331
rect 54518 31328 54530 31331
rect 56686 31328 56692 31340
rect 54518 31300 56692 31328
rect 54518 31297 54530 31300
rect 54472 31291 54530 31297
rect 56686 31288 56692 31300
rect 56744 31288 56750 31340
rect 25038 31260 25044 31272
rect 24999 31232 25044 31260
rect 25038 31220 25044 31232
rect 25096 31220 25102 31272
rect 27522 31220 27528 31272
rect 27580 31260 27586 31272
rect 27985 31263 28043 31269
rect 27985 31260 27997 31263
rect 27580 31232 27997 31260
rect 27580 31220 27586 31232
rect 27985 31229 27997 31232
rect 28031 31229 28043 31263
rect 33226 31260 33232 31272
rect 33187 31232 33232 31260
rect 27985 31223 28043 31229
rect 33226 31220 33232 31232
rect 33284 31220 33290 31272
rect 39574 31220 39580 31272
rect 39632 31260 39638 31272
rect 40497 31263 40555 31269
rect 40497 31260 40509 31263
rect 39632 31232 40509 31260
rect 39632 31220 39638 31232
rect 40497 31229 40509 31232
rect 40543 31229 40555 31263
rect 40497 31223 40555 31229
rect 52730 31220 52736 31272
rect 52788 31260 52794 31272
rect 54205 31263 54263 31269
rect 54205 31260 54217 31263
rect 52788 31232 54217 31260
rect 52788 31220 52794 31232
rect 54205 31229 54217 31232
rect 54251 31229 54263 31263
rect 54205 31223 54263 31229
rect 26234 31124 26240 31136
rect 24872 31096 26240 31124
rect 26234 31084 26240 31096
rect 26292 31084 26298 31136
rect 26418 31124 26424 31136
rect 26379 31096 26424 31124
rect 26418 31084 26424 31096
rect 26476 31084 26482 31136
rect 29362 31124 29368 31136
rect 29323 31096 29368 31124
rect 29362 31084 29368 31096
rect 29420 31084 29426 31136
rect 39666 31124 39672 31136
rect 39627 31096 39672 31124
rect 39666 31084 39672 31096
rect 39724 31084 39730 31136
rect 41690 31084 41696 31136
rect 41748 31124 41754 31136
rect 41877 31127 41935 31133
rect 41877 31124 41889 31127
rect 41748 31096 41889 31124
rect 41748 31084 41754 31096
rect 41877 31093 41889 31096
rect 41923 31093 41935 31127
rect 47026 31124 47032 31136
rect 46987 31096 47032 31124
rect 41877 31087 41935 31093
rect 47026 31084 47032 31096
rect 47084 31084 47090 31136
rect 55582 31124 55588 31136
rect 55543 31096 55588 31124
rect 55582 31084 55588 31096
rect 55640 31084 55646 31136
rect 1104 31034 59340 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 59340 31034
rect 1104 30960 59340 30982
rect 13449 30923 13507 30929
rect 13449 30889 13461 30923
rect 13495 30920 13507 30923
rect 13814 30920 13820 30932
rect 13495 30892 13820 30920
rect 13495 30889 13507 30892
rect 13449 30883 13507 30889
rect 13814 30880 13820 30892
rect 13872 30880 13878 30932
rect 15473 30923 15531 30929
rect 15473 30889 15485 30923
rect 15519 30920 15531 30923
rect 15562 30920 15568 30932
rect 15519 30892 15568 30920
rect 15519 30889 15531 30892
rect 15473 30883 15531 30889
rect 15562 30880 15568 30892
rect 15620 30880 15626 30932
rect 17310 30920 17316 30932
rect 17271 30892 17316 30920
rect 17310 30880 17316 30892
rect 17368 30880 17374 30932
rect 33226 30880 33232 30932
rect 33284 30920 33290 30932
rect 39298 30920 39304 30932
rect 33284 30892 39160 30920
rect 39259 30892 39304 30920
rect 33284 30880 33290 30892
rect 39132 30852 39160 30892
rect 39298 30880 39304 30892
rect 39356 30880 39362 30932
rect 52270 30920 52276 30932
rect 52231 30892 52276 30920
rect 52270 30880 52276 30892
rect 52328 30880 52334 30932
rect 58526 30920 58532 30932
rect 58487 30892 58532 30920
rect 58526 30880 58532 30892
rect 58584 30880 58590 30932
rect 41230 30852 41236 30864
rect 39132 30824 41236 30852
rect 41230 30812 41236 30824
rect 41288 30812 41294 30864
rect 11514 30744 11520 30796
rect 11572 30784 11578 30796
rect 12069 30787 12127 30793
rect 12069 30784 12081 30787
rect 11572 30756 12081 30784
rect 11572 30744 11578 30756
rect 12069 30753 12081 30756
rect 12115 30753 12127 30787
rect 22462 30784 22468 30796
rect 22423 30756 22468 30784
rect 12069 30747 12127 30753
rect 22462 30744 22468 30756
rect 22520 30744 22526 30796
rect 42794 30744 42800 30796
rect 42852 30784 42858 30796
rect 43073 30787 43131 30793
rect 43073 30784 43085 30787
rect 42852 30756 43085 30784
rect 42852 30744 42858 30756
rect 43073 30753 43085 30756
rect 43119 30753 43131 30787
rect 43073 30747 43131 30753
rect 47578 30744 47584 30796
rect 47636 30784 47642 30796
rect 48225 30787 48283 30793
rect 48225 30784 48237 30787
rect 47636 30756 48237 30784
rect 47636 30744 47642 30756
rect 48225 30753 48237 30756
rect 48271 30753 48283 30787
rect 48225 30747 48283 30753
rect 3881 30719 3939 30725
rect 3881 30685 3893 30719
rect 3927 30716 3939 30719
rect 4522 30716 4528 30728
rect 3927 30688 4528 30716
rect 3927 30685 3939 30688
rect 3881 30679 3939 30685
rect 4522 30676 4528 30688
rect 4580 30676 4586 30728
rect 6457 30719 6515 30725
rect 6457 30685 6469 30719
rect 6503 30716 6515 30719
rect 7006 30716 7012 30728
rect 6503 30688 7012 30716
rect 6503 30685 6515 30688
rect 6457 30679 6515 30685
rect 7006 30676 7012 30688
rect 7064 30676 7070 30728
rect 9306 30716 9312 30728
rect 9267 30688 9312 30716
rect 9306 30676 9312 30688
rect 9364 30676 9370 30728
rect 12336 30719 12394 30725
rect 12336 30685 12348 30719
rect 12382 30716 12394 30719
rect 12894 30716 12900 30728
rect 12382 30688 12900 30716
rect 12382 30685 12394 30688
rect 12336 30679 12394 30685
rect 12894 30676 12900 30688
rect 12952 30676 12958 30728
rect 14090 30716 14096 30728
rect 14051 30688 14096 30716
rect 14090 30676 14096 30688
rect 14148 30676 14154 30728
rect 14360 30719 14418 30725
rect 14360 30685 14372 30719
rect 14406 30716 14418 30719
rect 15470 30716 15476 30728
rect 14406 30688 15476 30716
rect 14406 30685 14418 30688
rect 14360 30679 14418 30685
rect 15470 30676 15476 30688
rect 15528 30676 15534 30728
rect 15930 30716 15936 30728
rect 15891 30688 15936 30716
rect 15930 30676 15936 30688
rect 15988 30676 15994 30728
rect 16206 30725 16212 30728
rect 16200 30716 16212 30725
rect 16167 30688 16212 30716
rect 16200 30679 16212 30688
rect 16206 30676 16212 30679
rect 16264 30676 16270 30728
rect 20622 30716 20628 30728
rect 20583 30688 20628 30716
rect 20622 30676 20628 30688
rect 20680 30676 20686 30728
rect 23750 30716 23756 30728
rect 22572 30688 23756 30716
rect 4148 30651 4206 30657
rect 4148 30617 4160 30651
rect 4194 30648 4206 30651
rect 5810 30648 5816 30660
rect 4194 30620 5816 30648
rect 4194 30617 4206 30620
rect 4148 30611 4206 30617
rect 5810 30608 5816 30620
rect 5868 30608 5874 30660
rect 6724 30651 6782 30657
rect 6724 30617 6736 30651
rect 6770 30648 6782 30651
rect 8202 30648 8208 30660
rect 6770 30620 8208 30648
rect 6770 30617 6782 30620
rect 6724 30611 6782 30617
rect 8202 30608 8208 30620
rect 8260 30608 8266 30660
rect 9576 30651 9634 30657
rect 9576 30617 9588 30651
rect 9622 30648 9634 30651
rect 10962 30648 10968 30660
rect 9622 30620 10968 30648
rect 9622 30617 9634 30620
rect 9576 30611 9634 30617
rect 10962 30608 10968 30620
rect 11020 30608 11026 30660
rect 20892 30651 20950 30657
rect 20892 30617 20904 30651
rect 20938 30648 20950 30651
rect 22572 30648 22600 30688
rect 23750 30676 23756 30688
rect 23808 30676 23814 30728
rect 24946 30676 24952 30728
rect 25004 30716 25010 30728
rect 25777 30719 25835 30725
rect 25777 30716 25789 30719
rect 25004 30688 25789 30716
rect 25004 30676 25010 30688
rect 25777 30685 25789 30688
rect 25823 30685 25835 30719
rect 25777 30679 25835 30685
rect 27522 30676 27528 30728
rect 27580 30716 27586 30728
rect 27617 30719 27675 30725
rect 27617 30716 27629 30719
rect 27580 30688 27629 30716
rect 27580 30676 27586 30688
rect 27617 30685 27629 30688
rect 27663 30685 27675 30719
rect 27617 30679 27675 30685
rect 27884 30719 27942 30725
rect 27884 30685 27896 30719
rect 27930 30716 27942 30719
rect 29362 30716 29368 30728
rect 27930 30688 29368 30716
rect 27930 30685 27942 30688
rect 27884 30679 27942 30685
rect 29362 30676 29368 30688
rect 29420 30676 29426 30728
rect 31113 30719 31171 30725
rect 31113 30685 31125 30719
rect 31159 30716 31171 30719
rect 32122 30716 32128 30728
rect 31159 30688 32128 30716
rect 31159 30685 31171 30688
rect 31113 30679 31171 30685
rect 32122 30676 32128 30688
rect 32180 30676 32186 30728
rect 34698 30716 34704 30728
rect 34659 30688 34704 30716
rect 34698 30676 34704 30688
rect 34756 30676 34762 30728
rect 34968 30719 35026 30725
rect 34968 30685 34980 30719
rect 35014 30716 35026 30719
rect 35986 30716 35992 30728
rect 35014 30688 35992 30716
rect 35014 30685 35026 30688
rect 34968 30679 35026 30685
rect 35986 30676 35992 30688
rect 36044 30676 36050 30728
rect 37921 30719 37979 30725
rect 37921 30685 37933 30719
rect 37967 30685 37979 30719
rect 37921 30679 37979 30685
rect 38188 30719 38246 30725
rect 38188 30685 38200 30719
rect 38234 30716 38246 30719
rect 39666 30716 39672 30728
rect 38234 30688 39672 30716
rect 38234 30685 38246 30688
rect 38188 30679 38246 30685
rect 20938 30620 22600 30648
rect 22732 30651 22790 30657
rect 20938 30617 20950 30620
rect 20892 30611 20950 30617
rect 22732 30617 22744 30651
rect 22778 30648 22790 30651
rect 24486 30648 24492 30660
rect 22778 30620 24492 30648
rect 22778 30617 22790 30620
rect 22732 30611 22790 30617
rect 24486 30608 24492 30620
rect 24544 30608 24550 30660
rect 26044 30651 26102 30657
rect 26044 30617 26056 30651
rect 26090 30648 26102 30651
rect 29270 30648 29276 30660
rect 26090 30620 29276 30648
rect 26090 30617 26102 30620
rect 26044 30611 26102 30617
rect 29270 30608 29276 30620
rect 29328 30608 29334 30660
rect 31380 30651 31438 30657
rect 31380 30617 31392 30651
rect 31426 30648 31438 30651
rect 33502 30648 33508 30660
rect 31426 30620 33508 30648
rect 31426 30617 31438 30620
rect 31380 30611 31438 30617
rect 33502 30608 33508 30620
rect 33560 30608 33566 30660
rect 37734 30608 37740 30660
rect 37792 30648 37798 30660
rect 37936 30648 37964 30679
rect 39666 30676 39672 30688
rect 39724 30676 39730 30728
rect 41233 30719 41291 30725
rect 41233 30685 41245 30719
rect 41279 30716 41291 30719
rect 42978 30716 42984 30728
rect 41279 30688 42984 30716
rect 41279 30685 41291 30688
rect 41233 30679 41291 30685
rect 42978 30676 42984 30688
rect 43036 30676 43042 30728
rect 44266 30716 44272 30728
rect 43272 30688 44272 30716
rect 39574 30648 39580 30660
rect 37792 30620 39580 30648
rect 37792 30608 37798 30620
rect 39574 30608 39580 30620
rect 39632 30608 39638 30660
rect 41500 30651 41558 30657
rect 41500 30617 41512 30651
rect 41546 30648 41558 30651
rect 43272 30648 43300 30688
rect 44266 30676 44272 30688
rect 44324 30676 44330 30728
rect 45646 30676 45652 30728
rect 45704 30716 45710 30728
rect 46385 30719 46443 30725
rect 46385 30716 46397 30719
rect 45704 30688 46397 30716
rect 45704 30676 45710 30688
rect 46385 30685 46397 30688
rect 46431 30685 46443 30719
rect 46385 30679 46443 30685
rect 48492 30719 48550 30725
rect 48492 30685 48504 30719
rect 48538 30716 48550 30719
rect 49602 30716 49608 30728
rect 48538 30688 49608 30716
rect 48538 30685 48550 30688
rect 48492 30679 48550 30685
rect 49602 30676 49608 30688
rect 49660 30676 49666 30728
rect 50798 30676 50804 30728
rect 50856 30716 50862 30728
rect 50893 30719 50951 30725
rect 50893 30716 50905 30719
rect 50856 30688 50905 30716
rect 50856 30676 50862 30688
rect 50893 30685 50905 30688
rect 50939 30685 50951 30719
rect 50893 30679 50951 30685
rect 51160 30719 51218 30725
rect 51160 30685 51172 30719
rect 51206 30716 51218 30719
rect 52454 30716 52460 30728
rect 51206 30688 52460 30716
rect 51206 30685 51218 30688
rect 51160 30679 51218 30685
rect 52454 30676 52460 30688
rect 52512 30676 52518 30728
rect 52730 30716 52736 30728
rect 52691 30688 52736 30716
rect 52730 30676 52736 30688
rect 52788 30716 52794 30728
rect 55582 30725 55588 30728
rect 55309 30719 55367 30725
rect 55309 30716 55321 30719
rect 52788 30688 55321 30716
rect 52788 30676 52794 30688
rect 55309 30685 55321 30688
rect 55355 30685 55367 30719
rect 55576 30716 55588 30725
rect 55543 30688 55588 30716
rect 55309 30679 55367 30685
rect 55576 30679 55588 30688
rect 55582 30676 55588 30679
rect 55640 30676 55646 30728
rect 57054 30676 57060 30728
rect 57112 30716 57118 30728
rect 57149 30719 57207 30725
rect 57149 30716 57161 30719
rect 57112 30688 57161 30716
rect 57112 30676 57118 30688
rect 57149 30685 57161 30688
rect 57195 30685 57207 30719
rect 57149 30679 57207 30685
rect 41546 30620 43300 30648
rect 43340 30651 43398 30657
rect 41546 30617 41558 30620
rect 41500 30611 41558 30617
rect 43340 30617 43352 30651
rect 43386 30648 43398 30651
rect 44358 30648 44364 30660
rect 43386 30620 44364 30648
rect 43386 30617 43398 30620
rect 43340 30611 43398 30617
rect 44358 30608 44364 30620
rect 44416 30608 44422 30660
rect 46652 30651 46710 30657
rect 46652 30617 46664 30651
rect 46698 30648 46710 30651
rect 47118 30648 47124 30660
rect 46698 30620 47124 30648
rect 46698 30617 46710 30620
rect 46652 30611 46710 30617
rect 47118 30608 47124 30620
rect 47176 30608 47182 30660
rect 53000 30651 53058 30657
rect 53000 30617 53012 30651
rect 53046 30648 53058 30651
rect 56594 30648 56600 30660
rect 53046 30620 56600 30648
rect 53046 30617 53058 30620
rect 53000 30611 53058 30617
rect 56594 30608 56600 30620
rect 56652 30608 56658 30660
rect 56778 30608 56784 30660
rect 56836 30648 56842 30660
rect 57394 30651 57452 30657
rect 57394 30648 57406 30651
rect 56836 30620 57406 30648
rect 56836 30608 56842 30620
rect 57394 30617 57406 30620
rect 57440 30617 57452 30651
rect 57394 30611 57452 30617
rect 5258 30580 5264 30592
rect 5219 30552 5264 30580
rect 5258 30540 5264 30552
rect 5316 30540 5322 30592
rect 6178 30540 6184 30592
rect 6236 30580 6242 30592
rect 7837 30583 7895 30589
rect 7837 30580 7849 30583
rect 6236 30552 7849 30580
rect 6236 30540 6242 30552
rect 7837 30549 7849 30552
rect 7883 30549 7895 30583
rect 7837 30543 7895 30549
rect 9674 30540 9680 30592
rect 9732 30580 9738 30592
rect 10689 30583 10747 30589
rect 10689 30580 10701 30583
rect 9732 30552 10701 30580
rect 9732 30540 9738 30552
rect 10689 30549 10701 30552
rect 10735 30549 10747 30583
rect 22002 30580 22008 30592
rect 21963 30552 22008 30580
rect 10689 30543 10747 30549
rect 22002 30540 22008 30552
rect 22060 30540 22066 30592
rect 23842 30580 23848 30592
rect 23803 30552 23848 30580
rect 23842 30540 23848 30552
rect 23900 30540 23906 30592
rect 27154 30580 27160 30592
rect 27115 30552 27160 30580
rect 27154 30540 27160 30552
rect 27212 30540 27218 30592
rect 28994 30580 29000 30592
rect 28955 30552 29000 30580
rect 28994 30540 29000 30552
rect 29052 30540 29058 30592
rect 31754 30540 31760 30592
rect 31812 30580 31818 30592
rect 32493 30583 32551 30589
rect 32493 30580 32505 30583
rect 31812 30552 32505 30580
rect 31812 30540 31818 30552
rect 32493 30549 32505 30552
rect 32539 30549 32551 30583
rect 36078 30580 36084 30592
rect 36039 30552 36084 30580
rect 32493 30543 32551 30549
rect 36078 30540 36084 30552
rect 36136 30540 36142 30592
rect 42610 30580 42616 30592
rect 42571 30552 42616 30580
rect 42610 30540 42616 30552
rect 42668 30540 42674 30592
rect 44174 30540 44180 30592
rect 44232 30580 44238 30592
rect 44453 30583 44511 30589
rect 44453 30580 44465 30583
rect 44232 30552 44465 30580
rect 44232 30540 44238 30552
rect 44453 30549 44465 30552
rect 44499 30549 44511 30583
rect 47762 30580 47768 30592
rect 47723 30552 47768 30580
rect 44453 30543 44511 30549
rect 47762 30540 47768 30552
rect 47820 30540 47826 30592
rect 49602 30580 49608 30592
rect 49563 30552 49608 30580
rect 49602 30540 49608 30552
rect 49660 30540 49666 30592
rect 54113 30583 54171 30589
rect 54113 30549 54125 30583
rect 54159 30580 54171 30583
rect 55398 30580 55404 30592
rect 54159 30552 55404 30580
rect 54159 30549 54171 30552
rect 54113 30543 54171 30549
rect 55398 30540 55404 30552
rect 55456 30540 55462 30592
rect 56689 30583 56747 30589
rect 56689 30549 56701 30583
rect 56735 30580 56747 30583
rect 57238 30580 57244 30592
rect 56735 30552 57244 30580
rect 56735 30549 56747 30552
rect 56689 30543 56747 30549
rect 57238 30540 57244 30552
rect 57296 30540 57302 30592
rect 1104 30490 59340 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 59340 30490
rect 1104 30416 59340 30438
rect 3970 30376 3976 30388
rect 3931 30348 3976 30376
rect 3970 30336 3976 30348
rect 4028 30336 4034 30388
rect 5810 30376 5816 30388
rect 5771 30348 5816 30376
rect 5810 30336 5816 30348
rect 5868 30336 5874 30388
rect 10962 30376 10968 30388
rect 10923 30348 10968 30376
rect 10962 30336 10968 30348
rect 11020 30336 11026 30388
rect 19334 30336 19340 30388
rect 19392 30376 19398 30388
rect 19429 30379 19487 30385
rect 19429 30376 19441 30379
rect 19392 30348 19441 30376
rect 19392 30336 19398 30348
rect 19429 30345 19441 30348
rect 19475 30345 19487 30379
rect 21266 30376 21272 30388
rect 21227 30348 21272 30376
rect 19429 30339 19487 30345
rect 21266 30336 21272 30348
rect 21324 30336 21330 30388
rect 24486 30336 24492 30388
rect 24544 30376 24550 30388
rect 24581 30379 24639 30385
rect 24581 30376 24593 30379
rect 24544 30348 24593 30376
rect 24544 30336 24550 30348
rect 24581 30345 24593 30348
rect 24627 30345 24639 30379
rect 29730 30376 29736 30388
rect 29691 30348 29736 30376
rect 24581 30339 24639 30345
rect 29730 30336 29736 30348
rect 29788 30336 29794 30388
rect 33502 30376 33508 30388
rect 33463 30348 33508 30376
rect 33502 30336 33508 30348
rect 33560 30336 33566 30388
rect 40586 30336 40592 30388
rect 40644 30376 40650 30388
rect 40957 30379 41015 30385
rect 40957 30376 40969 30379
rect 40644 30348 40969 30376
rect 40644 30336 40650 30348
rect 40957 30345 40969 30348
rect 41003 30345 41015 30379
rect 52178 30376 52184 30388
rect 52139 30348 52184 30376
rect 40957 30339 41015 30345
rect 52178 30336 52184 30348
rect 52236 30336 52242 30388
rect 56686 30376 56692 30388
rect 56647 30348 56692 30376
rect 56686 30336 56692 30348
rect 56744 30336 56750 30388
rect 14360 30311 14418 30317
rect 2608 30280 4476 30308
rect 2608 30249 2636 30280
rect 2593 30243 2651 30249
rect 2593 30209 2605 30243
rect 2639 30209 2651 30243
rect 2593 30203 2651 30209
rect 2860 30243 2918 30249
rect 2860 30209 2872 30243
rect 2906 30240 2918 30243
rect 3970 30240 3976 30252
rect 2906 30212 3976 30240
rect 2906 30209 2918 30212
rect 2860 30203 2918 30209
rect 3970 30200 3976 30212
rect 4028 30200 4034 30252
rect 4448 30249 4476 30280
rect 9600 30280 11560 30308
rect 4433 30243 4491 30249
rect 4433 30209 4445 30243
rect 4479 30240 4491 30243
rect 4522 30240 4528 30252
rect 4479 30212 4528 30240
rect 4479 30209 4491 30212
rect 4433 30203 4491 30209
rect 4522 30200 4528 30212
rect 4580 30200 4586 30252
rect 4700 30243 4758 30249
rect 4700 30209 4712 30243
rect 4746 30240 4758 30243
rect 5810 30240 5816 30252
rect 4746 30212 5816 30240
rect 4746 30209 4758 30212
rect 4700 30203 4758 30209
rect 5810 30200 5816 30212
rect 5868 30200 5874 30252
rect 8012 30243 8070 30249
rect 8012 30209 8024 30243
rect 8058 30240 8070 30243
rect 8386 30240 8392 30252
rect 8058 30212 8392 30240
rect 8058 30209 8070 30212
rect 8012 30203 8070 30209
rect 8386 30200 8392 30212
rect 8444 30200 8450 30252
rect 9600 30184 9628 30280
rect 11532 30252 11560 30280
rect 14360 30277 14372 30311
rect 14406 30308 14418 30311
rect 15654 30308 15660 30320
rect 14406 30280 15660 30308
rect 14406 30277 14418 30280
rect 14360 30271 14418 30277
rect 15654 30268 15660 30280
rect 15712 30268 15718 30320
rect 25308 30311 25366 30317
rect 25308 30277 25320 30311
rect 25354 30308 25366 30311
rect 26418 30308 26424 30320
rect 25354 30280 26424 30308
rect 25354 30277 25366 30280
rect 25308 30271 25366 30277
rect 26418 30268 26424 30280
rect 26476 30268 26482 30320
rect 28620 30311 28678 30317
rect 28620 30277 28632 30311
rect 28666 30308 28678 30311
rect 31202 30308 31208 30320
rect 28666 30280 31208 30308
rect 28666 30277 28678 30280
rect 28620 30271 28678 30277
rect 31202 30268 31208 30280
rect 31260 30268 31266 30320
rect 41230 30268 41236 30320
rect 41288 30308 41294 30320
rect 42518 30308 42524 30320
rect 41288 30280 42524 30308
rect 41288 30268 41294 30280
rect 42518 30268 42524 30280
rect 42576 30308 42582 30320
rect 42794 30308 42800 30320
rect 42576 30280 42800 30308
rect 42576 30268 42582 30280
rect 42794 30268 42800 30280
rect 42852 30268 42858 30320
rect 45916 30311 45974 30317
rect 45916 30277 45928 30311
rect 45962 30308 45974 30311
rect 47762 30308 47768 30320
rect 45962 30280 47768 30308
rect 45962 30277 45974 30280
rect 45916 30271 45974 30277
rect 47762 30268 47768 30280
rect 47820 30268 47826 30320
rect 51074 30317 51080 30320
rect 51068 30308 51080 30317
rect 51035 30280 51080 30308
rect 51068 30271 51080 30280
rect 51074 30268 51080 30271
rect 51132 30268 51138 30320
rect 9852 30243 9910 30249
rect 9852 30209 9864 30243
rect 9898 30240 9910 30243
rect 10870 30240 10876 30252
rect 9898 30212 10876 30240
rect 9898 30209 9910 30212
rect 9852 30203 9910 30209
rect 10870 30200 10876 30212
rect 10928 30200 10934 30252
rect 11514 30240 11520 30252
rect 11427 30212 11520 30240
rect 11514 30200 11520 30212
rect 11572 30200 11578 30252
rect 11784 30243 11842 30249
rect 11784 30209 11796 30243
rect 11830 30240 11842 30243
rect 13262 30240 13268 30252
rect 11830 30212 13268 30240
rect 11830 30209 11842 30212
rect 11784 30203 11842 30209
rect 13262 30200 13268 30212
rect 13320 30200 13326 30252
rect 13998 30200 14004 30252
rect 14056 30240 14062 30252
rect 14093 30243 14151 30249
rect 14093 30240 14105 30243
rect 14056 30212 14105 30240
rect 14056 30200 14062 30212
rect 14093 30209 14105 30212
rect 14139 30209 14151 30243
rect 14093 30203 14151 30209
rect 18316 30243 18374 30249
rect 18316 30209 18328 30243
rect 18362 30240 18374 30243
rect 19978 30240 19984 30252
rect 18362 30212 19984 30240
rect 18362 30209 18374 30212
rect 18316 30203 18374 30209
rect 19978 30200 19984 30212
rect 20036 30200 20042 30252
rect 20156 30243 20214 30249
rect 20156 30209 20168 30243
rect 20202 30240 20214 30243
rect 21910 30240 21916 30252
rect 20202 30212 21916 30240
rect 20202 30209 20214 30212
rect 20156 30203 20214 30209
rect 21910 30200 21916 30212
rect 21968 30200 21974 30252
rect 23468 30243 23526 30249
rect 23468 30209 23480 30243
rect 23514 30240 23526 30243
rect 25866 30240 25872 30252
rect 23514 30212 25872 30240
rect 23514 30209 23526 30212
rect 23468 30203 23526 30209
rect 25866 30200 25872 30212
rect 25924 30200 25930 30252
rect 28353 30243 28411 30249
rect 28353 30209 28365 30243
rect 28399 30240 28411 30243
rect 28902 30240 28908 30252
rect 28399 30212 28908 30240
rect 28399 30209 28411 30212
rect 28353 30203 28411 30209
rect 28902 30200 28908 30212
rect 28960 30240 28966 30252
rect 30193 30243 30251 30249
rect 30193 30240 30205 30243
rect 28960 30212 30205 30240
rect 28960 30200 28966 30212
rect 30193 30209 30205 30212
rect 30239 30209 30251 30243
rect 30193 30203 30251 30209
rect 30460 30243 30518 30249
rect 30460 30209 30472 30243
rect 30506 30240 30518 30243
rect 31386 30240 31392 30252
rect 30506 30212 31392 30240
rect 30506 30209 30518 30212
rect 30460 30203 30518 30209
rect 31386 30200 31392 30212
rect 31444 30200 31450 30252
rect 31570 30200 31576 30252
rect 31628 30240 31634 30252
rect 32381 30243 32439 30249
rect 32381 30240 32393 30243
rect 31628 30212 32393 30240
rect 31628 30200 31634 30212
rect 32381 30209 32393 30212
rect 32427 30209 32439 30243
rect 32381 30203 32439 30209
rect 34241 30243 34299 30249
rect 34241 30209 34253 30243
rect 34287 30240 34299 30243
rect 37734 30240 37740 30252
rect 34287 30212 35894 30240
rect 37695 30212 37740 30240
rect 34287 30209 34299 30212
rect 34241 30203 34299 30209
rect 6914 30132 6920 30184
rect 6972 30172 6978 30184
rect 7745 30175 7803 30181
rect 7745 30172 7757 30175
rect 6972 30144 7757 30172
rect 6972 30132 6978 30144
rect 7745 30141 7757 30144
rect 7791 30141 7803 30175
rect 7745 30135 7803 30141
rect 9306 30132 9312 30184
rect 9364 30172 9370 30184
rect 9582 30172 9588 30184
rect 9364 30144 9588 30172
rect 9364 30132 9370 30144
rect 9582 30132 9588 30144
rect 9640 30132 9646 30184
rect 15930 30132 15936 30184
rect 15988 30172 15994 30184
rect 18046 30172 18052 30184
rect 15988 30144 18052 30172
rect 15988 30132 15994 30144
rect 18046 30132 18052 30144
rect 18104 30132 18110 30184
rect 19889 30175 19947 30181
rect 19889 30141 19901 30175
rect 19935 30141 19947 30175
rect 23198 30172 23204 30184
rect 23159 30144 23204 30172
rect 19889 30135 19947 30141
rect 15378 30064 15384 30116
rect 15436 30104 15442 30116
rect 15473 30107 15531 30113
rect 15473 30104 15485 30107
rect 15436 30076 15485 30104
rect 15436 30064 15442 30076
rect 15473 30073 15485 30076
rect 15519 30073 15531 30107
rect 15473 30067 15531 30073
rect 9122 30036 9128 30048
rect 9083 30008 9128 30036
rect 9122 29996 9128 30008
rect 9180 29996 9186 30048
rect 12434 29996 12440 30048
rect 12492 30036 12498 30048
rect 12897 30039 12955 30045
rect 12897 30036 12909 30039
rect 12492 30008 12909 30036
rect 12492 29996 12498 30008
rect 12897 30005 12909 30008
rect 12943 30005 12955 30039
rect 12897 29999 12955 30005
rect 18046 29996 18052 30048
rect 18104 30036 18110 30048
rect 19242 30036 19248 30048
rect 18104 30008 19248 30036
rect 18104 29996 18110 30008
rect 19242 29996 19248 30008
rect 19300 30036 19306 30048
rect 19904 30036 19932 30135
rect 23198 30132 23204 30144
rect 23256 30132 23262 30184
rect 24946 30132 24952 30184
rect 25004 30172 25010 30184
rect 25041 30175 25099 30181
rect 25041 30172 25053 30175
rect 25004 30144 25053 30172
rect 25004 30132 25010 30144
rect 25041 30141 25053 30144
rect 25087 30141 25099 30175
rect 32122 30172 32128 30184
rect 32083 30144 32128 30172
rect 25041 30135 25099 30141
rect 32122 30132 32128 30144
rect 32180 30132 32186 30184
rect 26234 30064 26240 30116
rect 26292 30104 26298 30116
rect 26421 30107 26479 30113
rect 26421 30104 26433 30107
rect 26292 30076 26433 30104
rect 26292 30064 26298 30076
rect 26421 30073 26433 30076
rect 26467 30073 26479 30107
rect 26421 30067 26479 30073
rect 31478 30064 31484 30116
rect 31536 30104 31542 30116
rect 31573 30107 31631 30113
rect 31573 30104 31585 30107
rect 31536 30076 31585 30104
rect 31536 30064 31542 30076
rect 31573 30073 31585 30076
rect 31619 30073 31631 30107
rect 31573 30067 31631 30073
rect 19300 30008 19932 30036
rect 19300 29996 19306 30008
rect 34698 29996 34704 30048
rect 34756 30036 34762 30048
rect 35529 30039 35587 30045
rect 35529 30036 35541 30039
rect 34756 30008 35541 30036
rect 34756 29996 34762 30008
rect 35529 30005 35541 30008
rect 35575 30005 35587 30039
rect 35866 30036 35894 30212
rect 37734 30200 37740 30212
rect 37792 30200 37798 30252
rect 38004 30243 38062 30249
rect 38004 30209 38016 30243
rect 38050 30240 38062 30243
rect 38838 30240 38844 30252
rect 38050 30212 38844 30240
rect 38050 30209 38062 30212
rect 38004 30203 38062 30209
rect 38838 30200 38844 30212
rect 38896 30200 38902 30252
rect 39833 30243 39891 30249
rect 39833 30240 39845 30243
rect 39132 30212 39845 30240
rect 39132 30113 39160 30212
rect 39833 30209 39845 30212
rect 39879 30209 39891 30243
rect 39833 30203 39891 30209
rect 44076 30243 44134 30249
rect 44076 30209 44088 30243
rect 44122 30240 44134 30243
rect 47026 30240 47032 30252
rect 44122 30212 47032 30240
rect 44122 30209 44134 30212
rect 44076 30203 44134 30209
rect 47026 30200 47032 30212
rect 47084 30200 47090 30252
rect 49228 30243 49286 30249
rect 49228 30209 49240 30243
rect 49274 30240 49286 30243
rect 52546 30240 52552 30252
rect 49274 30212 52552 30240
rect 49274 30209 49286 30212
rect 49228 30203 49286 30209
rect 52546 30200 52552 30212
rect 52604 30200 52610 30252
rect 53006 30249 53012 30252
rect 53000 30203 53012 30249
rect 53064 30240 53070 30252
rect 55576 30243 55634 30249
rect 53064 30212 53100 30240
rect 53006 30200 53012 30203
rect 53064 30200 53070 30212
rect 55576 30209 55588 30243
rect 55622 30240 55634 30243
rect 56686 30240 56692 30252
rect 55622 30212 56692 30240
rect 55622 30209 55634 30212
rect 55576 30203 55634 30209
rect 56686 30200 56692 30212
rect 56744 30200 56750 30252
rect 39574 30172 39580 30184
rect 39535 30144 39580 30172
rect 39574 30132 39580 30144
rect 39632 30132 39638 30184
rect 42978 30132 42984 30184
rect 43036 30172 43042 30184
rect 43809 30175 43867 30181
rect 43809 30172 43821 30175
rect 43036 30144 43821 30172
rect 43036 30132 43042 30144
rect 43809 30141 43821 30144
rect 43855 30141 43867 30175
rect 45646 30172 45652 30184
rect 45607 30144 45652 30172
rect 43809 30135 43867 30141
rect 45646 30132 45652 30144
rect 45704 30132 45710 30184
rect 46842 30132 46848 30184
rect 46900 30172 46906 30184
rect 48961 30175 49019 30181
rect 48961 30172 48973 30175
rect 46900 30144 48973 30172
rect 46900 30132 46906 30144
rect 48961 30141 48973 30144
rect 49007 30141 49019 30175
rect 50798 30172 50804 30184
rect 50711 30144 50804 30172
rect 48961 30135 49019 30141
rect 39117 30107 39175 30113
rect 39117 30073 39129 30107
rect 39163 30073 39175 30107
rect 39117 30067 39175 30073
rect 38654 30036 38660 30048
rect 35866 30008 38660 30036
rect 35529 29999 35587 30005
rect 38654 29996 38660 30008
rect 38712 29996 38718 30048
rect 45189 30039 45247 30045
rect 45189 30005 45201 30039
rect 45235 30036 45247 30039
rect 45830 30036 45836 30048
rect 45235 30008 45836 30036
rect 45235 30005 45247 30008
rect 45189 29999 45247 30005
rect 45830 29996 45836 30008
rect 45888 29996 45894 30048
rect 47026 30036 47032 30048
rect 46987 30008 47032 30036
rect 47026 29996 47032 30008
rect 47084 29996 47090 30048
rect 48976 30036 49004 30135
rect 50798 30132 50804 30144
rect 50856 30132 50862 30184
rect 52730 30172 52736 30184
rect 52643 30144 52736 30172
rect 52730 30132 52736 30144
rect 52788 30132 52794 30184
rect 55309 30175 55367 30181
rect 55309 30141 55321 30175
rect 55355 30141 55367 30175
rect 55309 30135 55367 30141
rect 50154 30064 50160 30116
rect 50212 30104 50218 30116
rect 50341 30107 50399 30113
rect 50341 30104 50353 30107
rect 50212 30076 50353 30104
rect 50212 30064 50218 30076
rect 50341 30073 50353 30076
rect 50387 30073 50399 30107
rect 50341 30067 50399 30073
rect 50816 30036 50844 30132
rect 52748 30036 52776 30132
rect 54110 30036 54116 30048
rect 48976 30008 52776 30036
rect 54071 30008 54116 30036
rect 54110 29996 54116 30008
rect 54168 29996 54174 30048
rect 55324 30036 55352 30135
rect 57054 30036 57060 30048
rect 55324 30008 57060 30036
rect 57054 29996 57060 30008
rect 57112 29996 57118 30048
rect 1104 29946 59340 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 59340 29946
rect 1104 29872 59340 29894
rect 13262 29832 13268 29844
rect 13223 29804 13268 29832
rect 13262 29792 13268 29804
rect 13320 29792 13326 29844
rect 21910 29792 21916 29844
rect 21968 29832 21974 29844
rect 22005 29835 22063 29841
rect 22005 29832 22017 29835
rect 21968 29804 22017 29832
rect 21968 29792 21974 29804
rect 22005 29801 22017 29804
rect 22051 29801 22063 29835
rect 22005 29795 22063 29801
rect 27062 29792 27068 29844
rect 27120 29832 27126 29844
rect 27157 29835 27215 29841
rect 27157 29832 27169 29835
rect 27120 29804 27169 29832
rect 27120 29792 27126 29804
rect 27157 29801 27169 29804
rect 27203 29801 27215 29835
rect 27157 29795 27215 29801
rect 28997 29835 29055 29841
rect 28997 29801 29009 29835
rect 29043 29832 29055 29835
rect 29086 29832 29092 29844
rect 29043 29804 29092 29832
rect 29043 29801 29055 29804
rect 28997 29795 29055 29801
rect 29086 29792 29092 29804
rect 29144 29792 29150 29844
rect 31386 29832 31392 29844
rect 31347 29804 31392 29832
rect 31386 29792 31392 29804
rect 31444 29792 31450 29844
rect 37734 29832 37740 29844
rect 37476 29804 37740 29832
rect 11514 29656 11520 29708
rect 11572 29696 11578 29708
rect 11885 29699 11943 29705
rect 11885 29696 11897 29699
rect 11572 29668 11897 29696
rect 11572 29656 11578 29668
rect 11885 29665 11897 29668
rect 11931 29665 11943 29699
rect 11885 29659 11943 29665
rect 19242 29656 19248 29708
rect 19300 29696 19306 29708
rect 20622 29696 20628 29708
rect 19300 29668 20628 29696
rect 19300 29656 19306 29668
rect 20622 29656 20628 29668
rect 20680 29656 20686 29708
rect 28810 29656 28816 29708
rect 28868 29696 28874 29708
rect 37476 29705 37504 29804
rect 37734 29792 37740 29804
rect 37792 29792 37798 29844
rect 38838 29832 38844 29844
rect 38799 29804 38844 29832
rect 38838 29792 38844 29804
rect 38896 29792 38902 29844
rect 42426 29792 42432 29844
rect 42484 29832 42490 29844
rect 42613 29835 42671 29841
rect 42613 29832 42625 29835
rect 42484 29804 42625 29832
rect 42484 29792 42490 29804
rect 42613 29801 42625 29804
rect 42659 29801 42671 29835
rect 46842 29832 46848 29844
rect 42613 29795 42671 29801
rect 45756 29804 46848 29832
rect 30009 29699 30067 29705
rect 30009 29696 30021 29699
rect 28868 29668 30021 29696
rect 28868 29656 28874 29668
rect 30009 29665 30021 29668
rect 30055 29665 30067 29699
rect 30009 29659 30067 29665
rect 37461 29699 37519 29705
rect 37461 29665 37473 29699
rect 37507 29665 37519 29699
rect 41230 29696 41236 29708
rect 41191 29668 41236 29696
rect 37461 29659 37519 29665
rect 41230 29656 41236 29668
rect 41288 29656 41294 29708
rect 42978 29656 42984 29708
rect 43036 29696 43042 29708
rect 45756 29705 45784 29804
rect 46842 29792 46848 29804
rect 46900 29792 46906 29844
rect 47118 29832 47124 29844
rect 47079 29804 47124 29832
rect 47118 29792 47124 29804
rect 47176 29792 47182 29844
rect 53006 29792 53012 29844
rect 53064 29832 53070 29844
rect 53101 29835 53159 29841
rect 53101 29832 53113 29835
rect 53064 29804 53113 29832
rect 53064 29792 53070 29804
rect 53101 29801 53113 29804
rect 53147 29801 53159 29835
rect 56686 29832 56692 29844
rect 56647 29804 56692 29832
rect 53101 29795 53159 29801
rect 56686 29792 56692 29804
rect 56744 29792 56750 29844
rect 43073 29699 43131 29705
rect 43073 29696 43085 29699
rect 43036 29668 43085 29696
rect 43036 29656 43042 29668
rect 43073 29665 43085 29668
rect 43119 29665 43131 29699
rect 43073 29659 43131 29665
rect 45741 29699 45799 29705
rect 45741 29665 45753 29699
rect 45787 29665 45799 29699
rect 45741 29659 45799 29665
rect 50798 29656 50804 29708
rect 50856 29696 50862 29708
rect 51721 29699 51779 29705
rect 51721 29696 51733 29699
rect 50856 29668 51733 29696
rect 50856 29656 50862 29668
rect 51721 29665 51733 29668
rect 51767 29665 51779 29699
rect 51721 29659 51779 29665
rect 52730 29656 52736 29708
rect 52788 29696 52794 29708
rect 55309 29699 55367 29705
rect 55309 29696 55321 29699
rect 52788 29668 55321 29696
rect 52788 29656 52794 29668
rect 55309 29665 55321 29668
rect 55355 29665 55367 29699
rect 55309 29659 55367 29665
rect 5169 29631 5227 29637
rect 5169 29597 5181 29631
rect 5215 29597 5227 29631
rect 5169 29591 5227 29597
rect 5436 29631 5494 29637
rect 5436 29597 5448 29631
rect 5482 29628 5494 29631
rect 6178 29628 6184 29640
rect 5482 29600 6184 29628
rect 5482 29597 5494 29600
rect 5436 29591 5494 29597
rect 4430 29520 4436 29572
rect 4488 29560 4494 29572
rect 4614 29560 4620 29572
rect 4488 29532 4620 29560
rect 4488 29520 4494 29532
rect 4614 29520 4620 29532
rect 4672 29560 4678 29572
rect 4982 29560 4988 29572
rect 4672 29532 4988 29560
rect 4672 29520 4678 29532
rect 4982 29520 4988 29532
rect 5040 29560 5046 29572
rect 5184 29560 5212 29591
rect 6178 29588 6184 29600
rect 6236 29588 6242 29640
rect 7009 29631 7067 29637
rect 7009 29597 7021 29631
rect 7055 29597 7067 29631
rect 7009 29591 7067 29597
rect 7276 29631 7334 29637
rect 7276 29597 7288 29631
rect 7322 29628 7334 29631
rect 9122 29628 9128 29640
rect 7322 29600 9128 29628
rect 7322 29597 7334 29600
rect 7276 29591 7334 29597
rect 6914 29560 6920 29572
rect 5040 29532 6920 29560
rect 5040 29520 5046 29532
rect 6914 29520 6920 29532
rect 6972 29560 6978 29572
rect 7024 29560 7052 29591
rect 9122 29588 9128 29600
rect 9180 29588 9186 29640
rect 9582 29588 9588 29640
rect 9640 29628 9646 29640
rect 10045 29631 10103 29637
rect 10045 29628 10057 29631
rect 9640 29600 10057 29628
rect 9640 29588 9646 29600
rect 10045 29597 10057 29600
rect 10091 29597 10103 29631
rect 14642 29628 14648 29640
rect 14603 29600 14648 29628
rect 10045 29591 10103 29597
rect 14642 29588 14648 29600
rect 14700 29628 14706 29640
rect 15930 29628 15936 29640
rect 14700 29600 15936 29628
rect 14700 29588 14706 29600
rect 15930 29588 15936 29600
rect 15988 29588 15994 29640
rect 17034 29628 17040 29640
rect 16995 29600 17040 29628
rect 17034 29588 17040 29600
rect 17092 29588 17098 29640
rect 20892 29631 20950 29637
rect 20892 29597 20904 29631
rect 20938 29628 20950 29631
rect 22002 29628 22008 29640
rect 20938 29600 22008 29628
rect 20938 29597 20950 29600
rect 20892 29591 20950 29597
rect 22002 29588 22008 29600
rect 22060 29588 22066 29640
rect 22465 29631 22523 29637
rect 22465 29597 22477 29631
rect 22511 29597 22523 29631
rect 22465 29591 22523 29597
rect 22732 29631 22790 29637
rect 22732 29597 22744 29631
rect 22778 29628 22790 29631
rect 23842 29628 23848 29640
rect 22778 29600 23848 29628
rect 22778 29597 22790 29600
rect 22732 29591 22790 29597
rect 6972 29532 7052 29560
rect 10312 29563 10370 29569
rect 6972 29520 6978 29532
rect 10312 29529 10324 29563
rect 10358 29560 10370 29563
rect 10962 29560 10968 29572
rect 10358 29532 10968 29560
rect 10358 29529 10370 29532
rect 10312 29523 10370 29529
rect 10962 29520 10968 29532
rect 11020 29520 11026 29572
rect 12152 29563 12210 29569
rect 12152 29529 12164 29563
rect 12198 29560 12210 29563
rect 13538 29560 13544 29572
rect 12198 29532 13544 29560
rect 12198 29529 12210 29532
rect 12152 29523 12210 29529
rect 13538 29520 13544 29532
rect 13596 29520 13602 29572
rect 14912 29563 14970 29569
rect 14912 29529 14924 29563
rect 14958 29560 14970 29563
rect 16114 29560 16120 29572
rect 14958 29532 16120 29560
rect 14958 29529 14970 29532
rect 14912 29523 14970 29529
rect 16114 29520 16120 29532
rect 16172 29520 16178 29572
rect 17310 29569 17316 29572
rect 17304 29523 17316 29569
rect 17368 29560 17374 29572
rect 17368 29532 17404 29560
rect 17310 29520 17316 29523
rect 17368 29520 17374 29532
rect 20622 29520 20628 29572
rect 20680 29560 20686 29572
rect 22480 29560 22508 29591
rect 23842 29588 23848 29600
rect 23900 29588 23906 29640
rect 25038 29588 25044 29640
rect 25096 29628 25102 29640
rect 25777 29631 25835 29637
rect 25777 29628 25789 29631
rect 25096 29600 25789 29628
rect 25096 29588 25102 29600
rect 25777 29597 25789 29600
rect 25823 29628 25835 29631
rect 27522 29628 27528 29640
rect 25823 29600 27528 29628
rect 25823 29597 25835 29600
rect 25777 29591 25835 29597
rect 27522 29588 27528 29600
rect 27580 29628 27586 29640
rect 27617 29631 27675 29637
rect 27617 29628 27629 29631
rect 27580 29600 27629 29628
rect 27580 29588 27586 29600
rect 27617 29597 27629 29600
rect 27663 29597 27675 29631
rect 27617 29591 27675 29597
rect 27884 29631 27942 29637
rect 27884 29597 27896 29631
rect 27930 29628 27942 29631
rect 28994 29628 29000 29640
rect 27930 29600 29000 29628
rect 27930 29597 27942 29600
rect 27884 29591 27942 29597
rect 28994 29588 29000 29600
rect 29052 29588 29058 29640
rect 30276 29631 30334 29637
rect 30276 29597 30288 29631
rect 30322 29628 30334 29631
rect 31754 29628 31760 29640
rect 30322 29600 31760 29628
rect 30322 29597 30334 29600
rect 30276 29591 30334 29597
rect 31754 29588 31760 29600
rect 31812 29588 31818 29640
rect 31849 29631 31907 29637
rect 31849 29597 31861 29631
rect 31895 29628 31907 29631
rect 31938 29628 31944 29640
rect 31895 29600 31944 29628
rect 31895 29597 31907 29600
rect 31849 29591 31907 29597
rect 31938 29588 31944 29600
rect 31996 29588 32002 29640
rect 34698 29628 34704 29640
rect 34659 29600 34704 29628
rect 34698 29588 34704 29600
rect 34756 29588 34762 29640
rect 34968 29631 35026 29637
rect 34968 29597 34980 29631
rect 35014 29628 35026 29631
rect 36078 29628 36084 29640
rect 35014 29600 36084 29628
rect 35014 29597 35026 29600
rect 34968 29591 35026 29597
rect 36078 29588 36084 29600
rect 36136 29588 36142 29640
rect 41500 29631 41558 29637
rect 41500 29597 41512 29631
rect 41546 29628 41558 29631
rect 42610 29628 42616 29640
rect 41546 29600 42616 29628
rect 41546 29597 41558 29600
rect 41500 29591 41558 29597
rect 42610 29588 42616 29600
rect 42668 29588 42674 29640
rect 46008 29631 46066 29637
rect 46008 29597 46020 29631
rect 46054 29628 46066 29631
rect 49602 29628 49608 29640
rect 46054 29600 49608 29628
rect 46054 29597 46066 29600
rect 46008 29591 46066 29597
rect 49602 29588 49608 29600
rect 49660 29588 49666 29640
rect 55398 29588 55404 29640
rect 55456 29628 55462 29640
rect 55565 29631 55623 29637
rect 55565 29628 55577 29631
rect 55456 29600 55577 29628
rect 55456 29588 55462 29600
rect 55565 29597 55577 29600
rect 55611 29597 55623 29631
rect 55565 29591 55623 29597
rect 57054 29588 57060 29640
rect 57112 29628 57118 29640
rect 57149 29631 57207 29637
rect 57149 29628 57161 29631
rect 57112 29600 57161 29628
rect 57112 29588 57118 29600
rect 57149 29597 57161 29600
rect 57195 29597 57207 29631
rect 57149 29591 57207 29597
rect 57238 29588 57244 29640
rect 57296 29628 57302 29640
rect 57405 29631 57463 29637
rect 57405 29628 57417 29631
rect 57296 29600 57417 29628
rect 57296 29588 57302 29600
rect 57405 29597 57417 29600
rect 57451 29597 57463 29631
rect 57405 29591 57463 29597
rect 20680 29532 22508 29560
rect 26044 29563 26102 29569
rect 20680 29520 20686 29532
rect 26044 29529 26056 29563
rect 26090 29560 26102 29563
rect 28350 29560 28356 29572
rect 26090 29532 28356 29560
rect 26090 29529 26102 29532
rect 26044 29523 26102 29529
rect 28350 29520 28356 29532
rect 28408 29520 28414 29572
rect 32116 29563 32174 29569
rect 32116 29529 32128 29563
rect 32162 29560 32174 29563
rect 33778 29560 33784 29572
rect 32162 29532 33784 29560
rect 32162 29529 32174 29532
rect 32116 29523 32174 29529
rect 33778 29520 33784 29532
rect 33836 29520 33842 29572
rect 37728 29563 37786 29569
rect 37728 29529 37740 29563
rect 37774 29560 37786 29563
rect 38746 29560 38752 29572
rect 37774 29532 38752 29560
rect 37774 29529 37786 29532
rect 37728 29523 37786 29529
rect 38746 29520 38752 29532
rect 38804 29520 38810 29572
rect 43340 29563 43398 29569
rect 43340 29529 43352 29563
rect 43386 29560 43398 29563
rect 45094 29560 45100 29572
rect 43386 29532 45100 29560
rect 43386 29529 43398 29532
rect 43340 29523 43398 29529
rect 45094 29520 45100 29532
rect 45152 29520 45158 29572
rect 47581 29563 47639 29569
rect 47581 29529 47593 29563
rect 47627 29560 47639 29563
rect 47946 29560 47952 29572
rect 47627 29532 47952 29560
rect 47627 29529 47639 29532
rect 47581 29523 47639 29529
rect 47946 29520 47952 29532
rect 48004 29560 48010 29572
rect 51810 29560 51816 29572
rect 48004 29532 51816 29560
rect 48004 29520 48010 29532
rect 51810 29520 51816 29532
rect 51868 29520 51874 29572
rect 51988 29563 52046 29569
rect 51988 29529 52000 29563
rect 52034 29560 52046 29563
rect 54570 29560 54576 29572
rect 52034 29532 54576 29560
rect 52034 29529 52046 29532
rect 51988 29523 52046 29529
rect 54570 29520 54576 29532
rect 54628 29520 54634 29572
rect 6546 29492 6552 29504
rect 6507 29464 6552 29492
rect 6546 29452 6552 29464
rect 6604 29452 6610 29504
rect 7098 29452 7104 29504
rect 7156 29492 7162 29504
rect 8389 29495 8447 29501
rect 8389 29492 8401 29495
rect 7156 29464 8401 29492
rect 7156 29452 7162 29464
rect 8389 29461 8401 29464
rect 8435 29461 8447 29495
rect 11422 29492 11428 29504
rect 11383 29464 11428 29492
rect 8389 29455 8447 29461
rect 11422 29452 11428 29464
rect 11480 29452 11486 29504
rect 16022 29492 16028 29504
rect 15983 29464 16028 29492
rect 16022 29452 16028 29464
rect 16080 29452 16086 29504
rect 17954 29452 17960 29504
rect 18012 29492 18018 29504
rect 18417 29495 18475 29501
rect 18417 29492 18429 29495
rect 18012 29464 18429 29492
rect 18012 29452 18018 29464
rect 18417 29461 18429 29464
rect 18463 29461 18475 29495
rect 23842 29492 23848 29504
rect 23803 29464 23848 29492
rect 18417 29455 18475 29461
rect 23842 29452 23848 29464
rect 23900 29452 23906 29504
rect 30466 29452 30472 29504
rect 30524 29492 30530 29504
rect 33229 29495 33287 29501
rect 33229 29492 33241 29495
rect 30524 29464 33241 29492
rect 30524 29452 30530 29464
rect 33229 29461 33241 29464
rect 33275 29461 33287 29495
rect 36078 29492 36084 29504
rect 36039 29464 36084 29492
rect 33229 29455 33287 29461
rect 36078 29452 36084 29464
rect 36136 29452 36142 29504
rect 44450 29492 44456 29504
rect 44411 29464 44456 29492
rect 44450 29452 44456 29464
rect 44508 29452 44514 29504
rect 48314 29452 48320 29504
rect 48372 29492 48378 29504
rect 48869 29495 48927 29501
rect 48869 29492 48881 29495
rect 48372 29464 48881 29492
rect 48372 29452 48378 29464
rect 48869 29461 48881 29464
rect 48915 29461 48927 29495
rect 51828 29492 51856 29520
rect 56502 29492 56508 29504
rect 51828 29464 56508 29492
rect 48869 29455 48927 29461
rect 56502 29452 56508 29464
rect 56560 29452 56566 29504
rect 58529 29495 58587 29501
rect 58529 29461 58541 29495
rect 58575 29492 58587 29495
rect 59541 29495 59599 29501
rect 59541 29492 59553 29495
rect 58575 29464 59553 29492
rect 58575 29461 58587 29464
rect 58529 29455 58587 29461
rect 59541 29461 59553 29464
rect 59587 29461 59599 29495
rect 59541 29455 59599 29461
rect 1104 29402 59340 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 59340 29402
rect 1104 29328 59340 29350
rect 3970 29288 3976 29300
rect 3931 29260 3976 29288
rect 3970 29248 3976 29260
rect 4028 29248 4034 29300
rect 5810 29288 5816 29300
rect 5771 29260 5816 29288
rect 5810 29248 5816 29260
rect 5868 29248 5874 29300
rect 10870 29248 10876 29300
rect 10928 29288 10934 29300
rect 10965 29291 11023 29297
rect 10965 29288 10977 29291
rect 10928 29260 10977 29288
rect 10928 29248 10934 29260
rect 10965 29257 10977 29260
rect 11011 29257 11023 29291
rect 16114 29288 16120 29300
rect 16075 29260 16120 29288
rect 10965 29251 11023 29257
rect 16114 29248 16120 29260
rect 16172 29248 16178 29300
rect 20622 29248 20628 29300
rect 20680 29288 20686 29300
rect 20809 29291 20867 29297
rect 20809 29288 20821 29291
rect 20680 29260 20821 29288
rect 20680 29248 20686 29260
rect 20809 29257 20821 29260
rect 20855 29257 20867 29291
rect 25866 29288 25872 29300
rect 25827 29260 25872 29288
rect 20809 29251 20867 29257
rect 25866 29248 25872 29260
rect 25924 29248 25930 29300
rect 28626 29288 28632 29300
rect 28587 29260 28632 29288
rect 28626 29248 28632 29260
rect 28684 29248 28690 29300
rect 31570 29288 31576 29300
rect 31531 29260 31576 29288
rect 31570 29248 31576 29260
rect 31628 29248 31634 29300
rect 45646 29288 45652 29300
rect 45526 29260 45652 29288
rect 2860 29223 2918 29229
rect 2860 29189 2872 29223
rect 2906 29220 2918 29223
rect 5258 29220 5264 29232
rect 2906 29192 5264 29220
rect 2906 29189 2918 29192
rect 2860 29183 2918 29189
rect 5258 29180 5264 29192
rect 5316 29180 5322 29232
rect 6733 29223 6791 29229
rect 6733 29189 6745 29223
rect 6779 29220 6791 29223
rect 9852 29223 9910 29229
rect 6779 29192 6914 29220
rect 6779 29189 6791 29192
rect 6733 29183 6791 29189
rect 2593 29155 2651 29161
rect 2593 29121 2605 29155
rect 2639 29152 2651 29155
rect 4430 29152 4436 29164
rect 2639 29124 4436 29152
rect 2639 29121 2651 29124
rect 2593 29115 2651 29121
rect 4430 29112 4436 29124
rect 4488 29112 4494 29164
rect 4700 29155 4758 29161
rect 4700 29121 4712 29155
rect 4746 29152 4758 29155
rect 6362 29152 6368 29164
rect 4746 29124 6368 29152
rect 4746 29121 4758 29124
rect 4700 29115 4758 29121
rect 6362 29112 6368 29124
rect 6420 29112 6426 29164
rect 6886 29152 6914 29192
rect 9852 29189 9864 29223
rect 9898 29220 9910 29223
rect 11422 29220 11428 29232
rect 9898 29192 11428 29220
rect 9898 29189 9910 29192
rect 9852 29183 9910 29189
rect 11422 29180 11428 29192
rect 11480 29180 11486 29232
rect 13164 29223 13222 29229
rect 13164 29189 13176 29223
rect 13210 29220 13222 29223
rect 15470 29220 15476 29232
rect 13210 29192 15476 29220
rect 13210 29189 13222 29192
rect 13164 29183 13222 29189
rect 15470 29180 15476 29192
rect 15528 29180 15534 29232
rect 22732 29223 22790 29229
rect 22732 29189 22744 29223
rect 22778 29220 22790 29223
rect 23842 29220 23848 29232
rect 22778 29192 23848 29220
rect 22778 29189 22790 29192
rect 22732 29183 22790 29189
rect 23842 29180 23848 29192
rect 23900 29180 23906 29232
rect 24578 29180 24584 29232
rect 24636 29220 24642 29232
rect 24734 29223 24792 29229
rect 24734 29220 24746 29223
rect 24636 29192 24746 29220
rect 24636 29180 24642 29192
rect 24734 29189 24746 29192
rect 24780 29189 24792 29223
rect 24734 29183 24792 29189
rect 24946 29180 24952 29232
rect 25004 29180 25010 29232
rect 27154 29180 27160 29232
rect 27212 29220 27218 29232
rect 30466 29229 30472 29232
rect 27494 29223 27552 29229
rect 27494 29220 27506 29223
rect 27212 29192 27506 29220
rect 27212 29180 27218 29192
rect 27494 29189 27506 29192
rect 27540 29189 27552 29223
rect 30460 29220 30472 29229
rect 30427 29192 30472 29220
rect 27494 29183 27552 29189
rect 30460 29183 30472 29192
rect 30466 29180 30472 29183
rect 30524 29180 30530 29232
rect 33128 29223 33186 29229
rect 33128 29189 33140 29223
rect 33174 29220 33186 29223
rect 34968 29223 35026 29229
rect 33174 29192 34836 29220
rect 33174 29189 33186 29192
rect 33128 29183 33186 29189
rect 10686 29152 10692 29164
rect 6886 29124 10692 29152
rect 10686 29112 10692 29124
rect 10744 29112 10750 29164
rect 12897 29155 12955 29161
rect 12897 29121 12909 29155
rect 12943 29152 12955 29155
rect 14090 29152 14096 29164
rect 12943 29124 14096 29152
rect 12943 29121 12955 29124
rect 12897 29115 12955 29121
rect 14090 29112 14096 29124
rect 14148 29112 14154 29164
rect 14642 29112 14648 29164
rect 14700 29152 14706 29164
rect 14737 29155 14795 29161
rect 14737 29152 14749 29155
rect 14700 29124 14749 29152
rect 14700 29112 14706 29124
rect 14737 29121 14749 29124
rect 14783 29121 14795 29155
rect 14737 29115 14795 29121
rect 15004 29155 15062 29161
rect 15004 29121 15016 29155
rect 15050 29152 15062 29155
rect 16390 29152 16396 29164
rect 15050 29124 16396 29152
rect 15050 29121 15062 29124
rect 15004 29115 15062 29121
rect 16390 29112 16396 29124
rect 16448 29112 16454 29164
rect 17672 29155 17730 29161
rect 17672 29121 17684 29155
rect 17718 29152 17730 29155
rect 18690 29152 18696 29164
rect 17718 29124 18696 29152
rect 17718 29121 17730 29124
rect 17672 29115 17730 29121
rect 18690 29112 18696 29124
rect 18748 29112 18754 29164
rect 19521 29155 19579 29161
rect 19521 29121 19533 29155
rect 19567 29152 19579 29155
rect 20070 29152 20076 29164
rect 19567 29124 20076 29152
rect 19567 29121 19579 29124
rect 19521 29115 19579 29121
rect 20070 29112 20076 29124
rect 20128 29112 20134 29164
rect 23198 29152 23204 29164
rect 22480 29124 23204 29152
rect 22480 29096 22508 29124
rect 23198 29112 23204 29124
rect 23256 29152 23262 29164
rect 24489 29155 24547 29161
rect 24489 29152 24501 29155
rect 23256 29124 24501 29152
rect 23256 29112 23262 29124
rect 24489 29121 24501 29124
rect 24535 29152 24547 29155
rect 24964 29152 24992 29180
rect 25866 29152 25872 29164
rect 24535 29124 25872 29152
rect 24535 29121 24547 29124
rect 24489 29115 24547 29121
rect 25866 29112 25872 29124
rect 25924 29152 25930 29164
rect 27249 29155 27307 29161
rect 27249 29152 27261 29155
rect 25924 29124 27261 29152
rect 25924 29112 25930 29124
rect 27249 29121 27261 29124
rect 27295 29121 27307 29155
rect 27249 29115 27307 29121
rect 32122 29112 32128 29164
rect 32180 29152 32186 29164
rect 32861 29155 32919 29161
rect 32861 29152 32873 29155
rect 32180 29124 32873 29152
rect 32180 29112 32186 29124
rect 32861 29121 32873 29124
rect 32907 29152 32919 29155
rect 34808 29152 34836 29192
rect 34968 29189 34980 29223
rect 35014 29220 35026 29223
rect 36078 29220 36084 29232
rect 35014 29192 36084 29220
rect 35014 29189 35026 29192
rect 34968 29183 35026 29189
rect 36078 29180 36084 29192
rect 36136 29180 36142 29232
rect 37820 29223 37878 29229
rect 37820 29189 37832 29223
rect 37866 29220 37878 29223
rect 41874 29220 41880 29232
rect 37866 29192 41880 29220
rect 37866 29189 37878 29192
rect 37820 29183 37878 29189
rect 41874 29180 41880 29192
rect 41932 29180 41938 29232
rect 45526 29220 45554 29260
rect 45646 29248 45652 29260
rect 45704 29288 45710 29300
rect 48961 29291 49019 29297
rect 45704 29260 47624 29288
rect 45704 29248 45710 29260
rect 43824 29192 45554 29220
rect 45916 29223 45974 29229
rect 35986 29152 35992 29164
rect 32907 29124 34744 29152
rect 34808 29124 35992 29152
rect 32907 29121 32919 29124
rect 32861 29115 32919 29121
rect 34716 29096 34744 29124
rect 35986 29112 35992 29124
rect 36044 29112 36050 29164
rect 37553 29155 37611 29161
rect 37553 29121 37565 29155
rect 37599 29152 37611 29155
rect 39574 29152 39580 29164
rect 37599 29124 39580 29152
rect 37599 29121 37611 29124
rect 37553 29115 37611 29121
rect 9582 29084 9588 29096
rect 9543 29056 9588 29084
rect 9582 29044 9588 29056
rect 9640 29044 9646 29096
rect 16666 29044 16672 29096
rect 16724 29084 16730 29096
rect 17034 29084 17040 29096
rect 16724 29056 17040 29084
rect 16724 29044 16730 29056
rect 17034 29044 17040 29056
rect 17092 29084 17098 29096
rect 17405 29087 17463 29093
rect 17405 29084 17417 29087
rect 17092 29056 17417 29084
rect 17092 29044 17098 29056
rect 17405 29053 17417 29056
rect 17451 29053 17463 29087
rect 22462 29084 22468 29096
rect 22423 29056 22468 29084
rect 17405 29047 17463 29053
rect 22462 29044 22468 29056
rect 22520 29044 22526 29096
rect 28810 29044 28816 29096
rect 28868 29084 28874 29096
rect 30193 29087 30251 29093
rect 30193 29084 30205 29087
rect 28868 29056 30205 29084
rect 28868 29044 28874 29056
rect 30193 29053 30205 29056
rect 30239 29053 30251 29087
rect 34698 29084 34704 29096
rect 34659 29056 34704 29084
rect 30193 29047 30251 29053
rect 34698 29044 34704 29056
rect 34756 29044 34762 29096
rect 6914 28976 6920 29028
rect 6972 29016 6978 29028
rect 8021 29019 8079 29025
rect 8021 29016 8033 29019
rect 6972 28988 8033 29016
rect 6972 28976 6978 28988
rect 8021 28985 8033 28988
rect 8067 28985 8079 29019
rect 8021 28979 8079 28985
rect 23658 28976 23664 29028
rect 23716 29016 23722 29028
rect 23845 29019 23903 29025
rect 23845 29016 23857 29019
rect 23716 28988 23857 29016
rect 23716 28976 23722 28988
rect 23845 28985 23857 28988
rect 23891 28985 23903 29019
rect 23845 28979 23903 28985
rect 14274 28948 14280 28960
rect 14235 28920 14280 28948
rect 14274 28908 14280 28920
rect 14332 28908 14338 28960
rect 18782 28948 18788 28960
rect 18743 28920 18788 28948
rect 18782 28908 18788 28920
rect 18840 28908 18846 28960
rect 34238 28948 34244 28960
rect 34199 28920 34244 28948
rect 34238 28908 34244 28920
rect 34296 28908 34302 28960
rect 36078 28948 36084 28960
rect 36039 28920 36084 28948
rect 36078 28908 36084 28920
rect 36136 28908 36142 28960
rect 37366 28908 37372 28960
rect 37424 28948 37430 28960
rect 37568 28948 37596 29115
rect 39574 29112 39580 29124
rect 39632 29152 39638 29164
rect 39669 29155 39727 29161
rect 39669 29152 39681 29155
rect 39632 29124 39681 29152
rect 39632 29112 39638 29124
rect 39669 29121 39681 29124
rect 39715 29121 39727 29155
rect 39669 29115 39727 29121
rect 39936 29155 39994 29161
rect 39936 29121 39948 29155
rect 39982 29152 39994 29155
rect 41506 29152 41512 29164
rect 39982 29124 41512 29152
rect 39982 29121 39994 29124
rect 39936 29115 39994 29121
rect 41506 29112 41512 29124
rect 41564 29112 41570 29164
rect 42978 29112 42984 29164
rect 43036 29152 43042 29164
rect 43824 29161 43852 29192
rect 45916 29189 45928 29223
rect 45962 29220 45974 29223
rect 47026 29220 47032 29232
rect 45962 29192 47032 29220
rect 45962 29189 45974 29192
rect 45916 29183 45974 29189
rect 47026 29180 47032 29192
rect 47084 29180 47090 29232
rect 47596 29220 47624 29260
rect 48961 29257 48973 29291
rect 49007 29288 49019 29291
rect 49786 29288 49792 29300
rect 49007 29260 49792 29288
rect 49007 29257 49019 29260
rect 48961 29251 49019 29257
rect 49786 29248 49792 29260
rect 49844 29248 49850 29300
rect 56594 29248 56600 29300
rect 56652 29288 56658 29300
rect 56689 29291 56747 29297
rect 56689 29288 56701 29291
rect 56652 29260 56701 29288
rect 56652 29248 56658 29260
rect 56689 29257 56701 29260
rect 56735 29257 56747 29291
rect 56689 29251 56747 29257
rect 48314 29220 48320 29232
rect 47596 29192 48320 29220
rect 43809 29155 43867 29161
rect 43809 29152 43821 29155
rect 43036 29124 43821 29152
rect 43036 29112 43042 29124
rect 43809 29121 43821 29124
rect 43855 29121 43867 29155
rect 43809 29115 43867 29121
rect 44076 29155 44134 29161
rect 44076 29121 44088 29155
rect 44122 29152 44134 29155
rect 47118 29152 47124 29164
rect 44122 29124 47124 29152
rect 44122 29121 44134 29124
rect 44076 29115 44134 29121
rect 47118 29112 47124 29124
rect 47176 29112 47182 29164
rect 47596 29161 47624 29192
rect 48314 29180 48320 29192
rect 48372 29180 48378 29232
rect 51810 29180 51816 29232
rect 51868 29220 51874 29232
rect 53101 29223 53159 29229
rect 53101 29220 53113 29223
rect 51868 29192 53113 29220
rect 51868 29180 51874 29192
rect 53101 29189 53113 29192
rect 53147 29189 53159 29223
rect 53101 29183 53159 29189
rect 54110 29180 54116 29232
rect 54168 29220 54174 29232
rect 55554 29223 55612 29229
rect 55554 29220 55566 29223
rect 54168 29192 55566 29220
rect 54168 29180 54174 29192
rect 55554 29189 55566 29192
rect 55600 29189 55612 29223
rect 55554 29183 55612 29189
rect 47581 29155 47639 29161
rect 47581 29121 47593 29155
rect 47627 29121 47639 29155
rect 47581 29115 47639 29121
rect 47848 29155 47906 29161
rect 47848 29121 47860 29155
rect 47894 29152 47906 29155
rect 48958 29152 48964 29164
rect 47894 29124 48964 29152
rect 47894 29121 47906 29124
rect 47848 29115 47906 29121
rect 48958 29112 48964 29124
rect 49016 29112 49022 29164
rect 49688 29155 49746 29161
rect 49688 29121 49700 29155
rect 49734 29152 49746 29155
rect 50890 29152 50896 29164
rect 49734 29124 50896 29152
rect 49734 29121 49746 29124
rect 49688 29115 49746 29121
rect 50890 29112 50896 29124
rect 50948 29112 50954 29164
rect 55309 29155 55367 29161
rect 55309 29121 55321 29155
rect 55355 29152 55367 29155
rect 57054 29152 57060 29164
rect 55355 29124 57060 29152
rect 55355 29121 55367 29124
rect 55309 29115 55367 29121
rect 57054 29112 57060 29124
rect 57112 29112 57118 29164
rect 45646 29084 45652 29096
rect 45607 29056 45652 29084
rect 45646 29044 45652 29056
rect 45704 29044 45710 29096
rect 49418 29084 49424 29096
rect 49379 29056 49424 29084
rect 49418 29044 49424 29056
rect 49476 29044 49482 29096
rect 41046 29016 41052 29028
rect 41007 28988 41052 29016
rect 41046 28976 41052 28988
rect 41104 28976 41110 29028
rect 46934 28976 46940 29028
rect 46992 29016 46998 29028
rect 47029 29019 47087 29025
rect 47029 29016 47041 29019
rect 46992 28988 47041 29016
rect 46992 28976 46998 28988
rect 47029 28985 47041 28988
rect 47075 28985 47087 29019
rect 47029 28979 47087 28985
rect 50706 28976 50712 29028
rect 50764 29016 50770 29028
rect 50801 29019 50859 29025
rect 50801 29016 50813 29019
rect 50764 28988 50813 29016
rect 50764 28976 50770 28988
rect 50801 28985 50813 28988
rect 50847 28985 50859 29019
rect 50801 28979 50859 28985
rect 53190 28976 53196 29028
rect 53248 29016 53254 29028
rect 54389 29019 54447 29025
rect 54389 29016 54401 29019
rect 53248 28988 54401 29016
rect 53248 28976 53254 28988
rect 54389 28985 54401 28988
rect 54435 28985 54447 29019
rect 54389 28979 54447 28985
rect 38930 28948 38936 28960
rect 37424 28920 37596 28948
rect 38891 28920 38936 28948
rect 37424 28908 37430 28920
rect 38930 28908 38936 28920
rect 38988 28908 38994 28960
rect 45186 28948 45192 28960
rect 45147 28920 45192 28948
rect 45186 28908 45192 28920
rect 45244 28908 45250 28960
rect 1104 28858 59340 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 59340 28858
rect 1104 28784 59340 28806
rect 6362 28744 6368 28756
rect 6323 28716 6368 28744
rect 6362 28704 6368 28716
rect 6420 28704 6426 28756
rect 8386 28744 8392 28756
rect 8347 28716 8392 28744
rect 8386 28704 8392 28716
rect 8444 28704 8450 28756
rect 11514 28704 11520 28756
rect 11572 28744 11578 28756
rect 11977 28747 12035 28753
rect 11977 28744 11989 28747
rect 11572 28716 11989 28744
rect 11572 28704 11578 28716
rect 11977 28713 11989 28716
rect 12023 28713 12035 28747
rect 18690 28744 18696 28756
rect 18651 28716 18696 28744
rect 11977 28707 12035 28713
rect 18690 28704 18696 28716
rect 18748 28704 18754 28756
rect 19978 28704 19984 28756
rect 20036 28744 20042 28756
rect 20625 28747 20683 28753
rect 20625 28744 20637 28747
rect 20036 28716 20637 28744
rect 20036 28704 20042 28716
rect 20625 28713 20637 28716
rect 20671 28713 20683 28747
rect 33778 28744 33784 28756
rect 33739 28716 33784 28744
rect 20625 28707 20683 28713
rect 33778 28704 33784 28716
rect 33836 28704 33842 28756
rect 38746 28744 38752 28756
rect 38707 28716 38752 28744
rect 38746 28704 38752 28716
rect 38804 28704 38810 28756
rect 41506 28744 41512 28756
rect 41467 28716 41512 28744
rect 41506 28704 41512 28716
rect 41564 28704 41570 28756
rect 44358 28704 44364 28756
rect 44416 28744 44422 28756
rect 44453 28747 44511 28753
rect 44453 28744 44465 28747
rect 44416 28716 44465 28744
rect 44416 28704 44422 28716
rect 44453 28713 44465 28716
rect 44499 28713 44511 28747
rect 48958 28744 48964 28756
rect 48919 28716 48964 28744
rect 44453 28707 44511 28713
rect 48958 28704 48964 28716
rect 49016 28704 49022 28756
rect 54570 28744 54576 28756
rect 54531 28716 54576 28744
rect 54570 28704 54576 28716
rect 54628 28704 54634 28756
rect 4982 28608 4988 28620
rect 4943 28580 4988 28608
rect 4982 28568 4988 28580
rect 5040 28568 5046 28620
rect 37366 28608 37372 28620
rect 37327 28580 37372 28608
rect 37366 28568 37372 28580
rect 37424 28568 37430 28620
rect 39574 28568 39580 28620
rect 39632 28608 39638 28620
rect 39942 28608 39948 28620
rect 39632 28580 39948 28608
rect 39632 28568 39638 28580
rect 39942 28568 39948 28580
rect 40000 28608 40006 28620
rect 40129 28611 40187 28617
rect 40129 28608 40141 28611
rect 40000 28580 40141 28608
rect 40000 28568 40006 28580
rect 40129 28577 40141 28580
rect 40175 28577 40187 28611
rect 40129 28571 40187 28577
rect 42978 28568 42984 28620
rect 43036 28608 43042 28620
rect 43073 28611 43131 28617
rect 43073 28608 43085 28611
rect 43036 28580 43085 28608
rect 43036 28568 43042 28580
rect 43073 28577 43085 28580
rect 43119 28577 43131 28611
rect 43073 28571 43131 28577
rect 52730 28568 52736 28620
rect 52788 28608 52794 28620
rect 53190 28608 53196 28620
rect 52788 28580 53196 28608
rect 52788 28568 52794 28580
rect 53190 28568 53196 28580
rect 53248 28568 53254 28620
rect 5252 28543 5310 28549
rect 5252 28509 5264 28543
rect 5298 28540 5310 28543
rect 6546 28540 6552 28552
rect 5298 28512 6552 28540
rect 5298 28509 5310 28512
rect 5252 28503 5310 28509
rect 6546 28500 6552 28512
rect 6604 28500 6610 28552
rect 7009 28543 7067 28549
rect 7009 28509 7021 28543
rect 7055 28540 7067 28543
rect 8294 28540 8300 28552
rect 7055 28512 8300 28540
rect 7055 28509 7067 28512
rect 7009 28503 7067 28509
rect 8294 28500 8300 28512
rect 8352 28500 8358 28552
rect 10686 28540 10692 28552
rect 10647 28512 10692 28540
rect 10686 28500 10692 28512
rect 10744 28540 10750 28552
rect 12526 28540 12532 28552
rect 10744 28512 12532 28540
rect 10744 28500 10750 28512
rect 12526 28500 12532 28512
rect 12584 28500 12590 28552
rect 15473 28543 15531 28549
rect 15473 28509 15485 28543
rect 15519 28540 15531 28543
rect 16666 28540 16672 28552
rect 15519 28512 16672 28540
rect 15519 28509 15531 28512
rect 15473 28503 15531 28509
rect 16666 28500 16672 28512
rect 16724 28500 16730 28552
rect 17313 28543 17371 28549
rect 17313 28509 17325 28543
rect 17359 28540 17371 28543
rect 18046 28540 18052 28552
rect 17359 28512 18052 28540
rect 17359 28509 17371 28512
rect 17313 28503 17371 28509
rect 18046 28500 18052 28512
rect 18104 28540 18110 28552
rect 19242 28540 19248 28552
rect 18104 28512 19248 28540
rect 18104 28500 18110 28512
rect 19242 28500 19248 28512
rect 19300 28500 19306 28552
rect 19512 28543 19570 28549
rect 19512 28509 19524 28543
rect 19558 28540 19570 28543
rect 20990 28540 20996 28552
rect 19558 28512 20996 28540
rect 19558 28509 19570 28512
rect 19512 28503 19570 28509
rect 20990 28500 20996 28512
rect 21048 28500 21054 28552
rect 21821 28543 21879 28549
rect 21821 28509 21833 28543
rect 21867 28540 21879 28543
rect 22462 28540 22468 28552
rect 21867 28512 22468 28540
rect 21867 28509 21879 28512
rect 21821 28503 21879 28509
rect 22462 28500 22468 28512
rect 22520 28500 22526 28552
rect 25130 28540 25136 28552
rect 25091 28512 25136 28540
rect 25130 28500 25136 28512
rect 25188 28500 25194 28552
rect 26973 28543 27031 28549
rect 26973 28509 26985 28543
rect 27019 28540 27031 28543
rect 27614 28540 27620 28552
rect 27019 28512 27620 28540
rect 27019 28509 27031 28512
rect 26973 28503 27031 28509
rect 27614 28500 27620 28512
rect 27672 28500 27678 28552
rect 29546 28540 29552 28552
rect 29507 28512 29552 28540
rect 29546 28500 29552 28512
rect 29604 28500 29610 28552
rect 32401 28543 32459 28549
rect 32401 28509 32413 28543
rect 32447 28509 32459 28543
rect 32401 28503 32459 28509
rect 32668 28543 32726 28549
rect 32668 28509 32680 28543
rect 32714 28540 32726 28543
rect 34238 28540 34244 28552
rect 32714 28512 34244 28540
rect 32714 28509 32726 28512
rect 32668 28503 32726 28509
rect 7276 28475 7334 28481
rect 7276 28441 7288 28475
rect 7322 28472 7334 28475
rect 9122 28472 9128 28484
rect 7322 28444 9128 28472
rect 7322 28441 7334 28444
rect 7276 28435 7334 28441
rect 9122 28432 9128 28444
rect 9180 28432 9186 28484
rect 15740 28475 15798 28481
rect 15740 28441 15752 28475
rect 15786 28472 15798 28475
rect 17580 28475 17638 28481
rect 15786 28444 17540 28472
rect 15786 28441 15798 28444
rect 15740 28435 15798 28441
rect 16850 28404 16856 28416
rect 16811 28376 16856 28404
rect 16850 28364 16856 28376
rect 16908 28364 16914 28416
rect 17512 28404 17540 28444
rect 17580 28441 17592 28475
rect 17626 28472 17638 28475
rect 22088 28475 22146 28481
rect 17626 28444 19472 28472
rect 17626 28441 17638 28444
rect 17580 28435 17638 28441
rect 18046 28404 18052 28416
rect 17512 28376 18052 28404
rect 18046 28364 18052 28376
rect 18104 28364 18110 28416
rect 19444 28404 19472 28444
rect 22088 28441 22100 28475
rect 22134 28472 22146 28475
rect 23474 28472 23480 28484
rect 22134 28444 23480 28472
rect 22134 28441 22146 28444
rect 22088 28435 22146 28441
rect 23474 28432 23480 28444
rect 23532 28432 23538 28484
rect 25400 28475 25458 28481
rect 25400 28441 25412 28475
rect 25446 28472 25458 28475
rect 27062 28472 27068 28484
rect 25446 28444 27068 28472
rect 25446 28441 25458 28444
rect 25400 28435 25458 28441
rect 27062 28432 27068 28444
rect 27120 28432 27126 28484
rect 27240 28475 27298 28481
rect 27240 28441 27252 28475
rect 27286 28472 27298 28475
rect 28074 28472 28080 28484
rect 27286 28444 28080 28472
rect 27286 28441 27298 28444
rect 27240 28435 27298 28441
rect 28074 28432 28080 28444
rect 28132 28432 28138 28484
rect 29794 28475 29852 28481
rect 29794 28472 29806 28475
rect 28184 28444 29806 28472
rect 20530 28404 20536 28416
rect 19444 28376 20536 28404
rect 20530 28364 20536 28376
rect 20588 28364 20594 28416
rect 23198 28404 23204 28416
rect 23159 28376 23204 28404
rect 23198 28364 23204 28376
rect 23256 28364 23262 28416
rect 26513 28407 26571 28413
rect 26513 28373 26525 28407
rect 26559 28404 26571 28407
rect 28184 28404 28212 28444
rect 29794 28441 29806 28444
rect 29840 28441 29852 28475
rect 32416 28472 32444 28503
rect 34238 28500 34244 28512
rect 34296 28500 34302 28552
rect 34698 28500 34704 28552
rect 34756 28540 34762 28552
rect 34793 28543 34851 28549
rect 34793 28540 34805 28543
rect 34756 28512 34805 28540
rect 34756 28500 34762 28512
rect 34793 28509 34805 28512
rect 34839 28509 34851 28543
rect 34793 28503 34851 28509
rect 35060 28543 35118 28549
rect 35060 28509 35072 28543
rect 35106 28540 35118 28543
rect 36078 28540 36084 28552
rect 35106 28512 36084 28540
rect 35106 28509 35118 28512
rect 35060 28503 35118 28509
rect 36078 28500 36084 28512
rect 36136 28500 36142 28552
rect 37636 28543 37694 28549
rect 37636 28509 37648 28543
rect 37682 28540 37694 28543
rect 38930 28540 38936 28552
rect 37682 28512 38936 28540
rect 37682 28509 37694 28512
rect 37636 28503 37694 28509
rect 38930 28500 38936 28512
rect 38988 28500 38994 28552
rect 43340 28543 43398 28549
rect 43340 28509 43352 28543
rect 43386 28540 43398 28543
rect 44450 28540 44456 28552
rect 43386 28512 44456 28540
rect 43386 28509 43398 28512
rect 43340 28503 43398 28509
rect 44450 28500 44456 28512
rect 44508 28500 44514 28552
rect 45741 28543 45799 28549
rect 45741 28509 45753 28543
rect 45787 28509 45799 28543
rect 45741 28503 45799 28509
rect 33134 28472 33140 28484
rect 32416 28444 33140 28472
rect 29794 28435 29852 28441
rect 33134 28432 33140 28444
rect 33192 28432 33198 28484
rect 40396 28475 40454 28481
rect 40396 28441 40408 28475
rect 40442 28472 40454 28475
rect 40678 28472 40684 28484
rect 40442 28444 40684 28472
rect 40442 28441 40454 28444
rect 40396 28435 40454 28441
rect 40678 28432 40684 28444
rect 40736 28432 40742 28484
rect 45646 28432 45652 28484
rect 45704 28472 45710 28484
rect 45756 28472 45784 28503
rect 45830 28500 45836 28552
rect 45888 28540 45894 28552
rect 45997 28543 46055 28549
rect 45997 28540 46009 28543
rect 45888 28512 46009 28540
rect 45888 28500 45894 28512
rect 45997 28509 46009 28512
rect 46043 28509 46055 28543
rect 45997 28503 46055 28509
rect 47581 28543 47639 28549
rect 47581 28509 47593 28543
rect 47627 28540 47639 28543
rect 48314 28540 48320 28552
rect 47627 28512 48320 28540
rect 47627 28509 47639 28512
rect 47581 28503 47639 28509
rect 47596 28472 47624 28503
rect 48314 28500 48320 28512
rect 48372 28500 48378 28552
rect 50154 28540 50160 28552
rect 50067 28512 50160 28540
rect 50154 28500 50160 28512
rect 50212 28540 50218 28552
rect 50798 28540 50804 28552
rect 50212 28512 50804 28540
rect 50212 28500 50218 28512
rect 50798 28500 50804 28512
rect 50856 28500 50862 28552
rect 57054 28540 57060 28552
rect 57015 28512 57060 28540
rect 57054 28500 57060 28512
rect 57112 28500 57118 28552
rect 45704 28444 47624 28472
rect 47848 28475 47906 28481
rect 45704 28432 45710 28444
rect 47848 28441 47860 28475
rect 47894 28472 47906 28475
rect 49050 28472 49056 28484
rect 47894 28444 49056 28472
rect 47894 28441 47906 28444
rect 47848 28435 47906 28441
rect 49050 28432 49056 28444
rect 49108 28432 49114 28484
rect 50424 28475 50482 28481
rect 50424 28441 50436 28475
rect 50470 28472 50482 28475
rect 51442 28472 51448 28484
rect 50470 28444 51448 28472
rect 50470 28441 50482 28444
rect 50424 28435 50482 28441
rect 51442 28432 51448 28444
rect 51500 28432 51506 28484
rect 53460 28475 53518 28481
rect 53460 28441 53472 28475
rect 53506 28472 53518 28475
rect 54754 28472 54760 28484
rect 53506 28444 54760 28472
rect 53506 28441 53518 28444
rect 53460 28435 53518 28441
rect 54754 28432 54760 28444
rect 54812 28432 54818 28484
rect 56686 28432 56692 28484
rect 56744 28472 56750 28484
rect 57302 28475 57360 28481
rect 57302 28472 57314 28475
rect 56744 28444 57314 28472
rect 56744 28432 56750 28444
rect 57302 28441 57314 28444
rect 57348 28441 57360 28475
rect 57302 28435 57360 28441
rect 28350 28404 28356 28416
rect 26559 28376 28212 28404
rect 28311 28376 28356 28404
rect 26559 28373 26571 28376
rect 26513 28367 26571 28373
rect 28350 28364 28356 28376
rect 28408 28364 28414 28416
rect 30929 28407 30987 28413
rect 30929 28373 30941 28407
rect 30975 28404 30987 28407
rect 31478 28404 31484 28416
rect 30975 28376 31484 28404
rect 30975 28373 30987 28376
rect 30929 28367 30987 28373
rect 31478 28364 31484 28376
rect 31536 28364 31542 28416
rect 36170 28404 36176 28416
rect 36131 28376 36176 28404
rect 36170 28364 36176 28376
rect 36228 28364 36234 28416
rect 47118 28404 47124 28416
rect 47079 28376 47124 28404
rect 47118 28364 47124 28376
rect 47176 28364 47182 28416
rect 50614 28364 50620 28416
rect 50672 28404 50678 28416
rect 51537 28407 51595 28413
rect 51537 28404 51549 28407
rect 50672 28376 51549 28404
rect 50672 28364 50678 28376
rect 51537 28373 51549 28376
rect 51583 28373 51595 28407
rect 51537 28367 51595 28373
rect 58437 28407 58495 28413
rect 58437 28373 58449 28407
rect 58483 28404 58495 28407
rect 59449 28407 59507 28413
rect 59449 28404 59461 28407
rect 58483 28376 59461 28404
rect 58483 28373 58495 28376
rect 58437 28367 58495 28373
rect 59449 28373 59461 28376
rect 59495 28373 59507 28407
rect 59449 28367 59507 28373
rect 1104 28314 59340 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 59340 28314
rect 1104 28240 59340 28262
rect 9122 28200 9128 28212
rect 9083 28172 9128 28200
rect 9122 28160 9128 28172
rect 9180 28160 9186 28212
rect 10962 28200 10968 28212
rect 10923 28172 10968 28200
rect 10962 28160 10968 28172
rect 11020 28160 11026 28212
rect 25866 28200 25872 28212
rect 25827 28172 25872 28200
rect 25866 28160 25872 28172
rect 25924 28160 25930 28212
rect 27062 28160 27068 28212
rect 27120 28200 27126 28212
rect 30193 28203 30251 28209
rect 30193 28200 30205 28203
rect 27120 28172 30205 28200
rect 27120 28160 27126 28172
rect 30193 28169 30205 28172
rect 30239 28169 30251 28203
rect 39942 28200 39948 28212
rect 39903 28172 39948 28200
rect 30193 28163 30251 28169
rect 39942 28160 39948 28172
rect 40000 28160 40006 28212
rect 42978 28160 42984 28212
rect 43036 28200 43042 28212
rect 45646 28200 45652 28212
rect 43036 28172 45652 28200
rect 43036 28160 43042 28172
rect 45646 28160 45652 28172
rect 45704 28160 45710 28212
rect 47026 28200 47032 28212
rect 46987 28172 47032 28200
rect 47026 28160 47032 28172
rect 47084 28160 47090 28212
rect 49050 28200 49056 28212
rect 49011 28172 49056 28200
rect 49050 28160 49056 28172
rect 49108 28160 49114 28212
rect 50890 28200 50896 28212
rect 50851 28172 50896 28200
rect 50890 28160 50896 28172
rect 50948 28160 50954 28212
rect 54754 28200 54760 28212
rect 54715 28172 54760 28200
rect 54754 28160 54760 28172
rect 54812 28160 54818 28212
rect 8012 28135 8070 28141
rect 8012 28101 8024 28135
rect 8058 28132 8070 28135
rect 9674 28132 9680 28144
rect 8058 28104 9680 28132
rect 8058 28101 8070 28104
rect 8012 28095 8070 28101
rect 9674 28092 9680 28104
rect 9732 28092 9738 28144
rect 9852 28135 9910 28141
rect 9852 28101 9864 28135
rect 9898 28132 9910 28135
rect 12434 28132 12440 28144
rect 9898 28104 12440 28132
rect 9898 28101 9910 28104
rect 9852 28095 9910 28101
rect 12434 28092 12440 28104
rect 12492 28092 12498 28144
rect 12980 28135 13038 28141
rect 12980 28101 12992 28135
rect 13026 28132 13038 28135
rect 14274 28132 14280 28144
rect 13026 28104 14280 28132
rect 13026 28101 13038 28104
rect 12980 28095 13038 28101
rect 14274 28092 14280 28104
rect 14332 28092 14338 28144
rect 15004 28135 15062 28141
rect 15004 28101 15016 28135
rect 15050 28132 15062 28135
rect 16850 28132 16856 28144
rect 15050 28104 16856 28132
rect 15050 28101 15062 28104
rect 15004 28095 15062 28101
rect 16850 28092 16856 28104
rect 16908 28092 16914 28144
rect 17304 28135 17362 28141
rect 17304 28101 17316 28135
rect 17350 28132 17362 28135
rect 18782 28132 18788 28144
rect 17350 28104 18788 28132
rect 17350 28101 17362 28104
rect 17304 28095 17362 28101
rect 18782 28092 18788 28104
rect 18840 28092 18846 28144
rect 19426 28092 19432 28144
rect 19484 28141 19490 28144
rect 19484 28135 19548 28141
rect 19484 28101 19502 28135
rect 19536 28101 19548 28135
rect 27614 28132 27620 28144
rect 19484 28095 19548 28101
rect 26988 28104 27620 28132
rect 19484 28092 19490 28095
rect 7745 28067 7803 28073
rect 7745 28033 7757 28067
rect 7791 28064 7803 28067
rect 8294 28064 8300 28076
rect 7791 28036 8300 28064
rect 7791 28033 7803 28036
rect 7745 28027 7803 28033
rect 8294 28024 8300 28036
rect 8352 28064 8358 28076
rect 8352 28036 9628 28064
rect 8352 28024 8358 28036
rect 9600 28008 9628 28036
rect 12250 28024 12256 28076
rect 12308 28064 12314 28076
rect 12713 28067 12771 28073
rect 12713 28064 12725 28067
rect 12308 28036 12725 28064
rect 12308 28024 12314 28036
rect 12713 28033 12725 28036
rect 12759 28064 12771 28067
rect 14090 28064 14096 28076
rect 12759 28036 14096 28064
rect 12759 28033 12771 28036
rect 12713 28027 12771 28033
rect 14090 28024 14096 28036
rect 14148 28064 14154 28076
rect 14737 28067 14795 28073
rect 14737 28064 14749 28067
rect 14148 28036 14749 28064
rect 14148 28024 14154 28036
rect 14737 28033 14749 28036
rect 14783 28033 14795 28067
rect 19242 28064 19248 28076
rect 19203 28036 19248 28064
rect 14737 28027 14795 28033
rect 19242 28024 19248 28036
rect 19300 28024 19306 28076
rect 23008 28067 23066 28073
rect 23008 28033 23020 28067
rect 23054 28064 23066 28067
rect 24486 28064 24492 28076
rect 23054 28036 24492 28064
rect 23054 28033 23066 28036
rect 23008 28027 23066 28033
rect 24486 28024 24492 28036
rect 24544 28024 24550 28076
rect 24581 28067 24639 28073
rect 24581 28033 24593 28067
rect 24627 28064 24639 28067
rect 24762 28064 24768 28076
rect 24627 28036 24768 28064
rect 24627 28033 24639 28036
rect 24581 28027 24639 28033
rect 24762 28024 24768 28036
rect 24820 28024 24826 28076
rect 26988 28073 27016 28104
rect 27614 28092 27620 28104
rect 27672 28132 27678 28144
rect 27672 28104 28304 28132
rect 27672 28092 27678 28104
rect 26973 28067 27031 28073
rect 26973 28033 26985 28067
rect 27019 28033 27031 28067
rect 26973 28027 27031 28033
rect 27240 28067 27298 28073
rect 27240 28033 27252 28067
rect 27286 28064 27298 28067
rect 28166 28064 28172 28076
rect 27286 28036 28172 28064
rect 27286 28033 27298 28036
rect 27240 28027 27298 28033
rect 28166 28024 28172 28036
rect 28224 28024 28230 28076
rect 28276 28064 28304 28104
rect 28350 28092 28356 28144
rect 28408 28132 28414 28144
rect 29058 28135 29116 28141
rect 29058 28132 29070 28135
rect 28408 28104 29070 28132
rect 28408 28092 28414 28104
rect 29058 28101 29070 28104
rect 29104 28101 29116 28135
rect 29058 28095 29116 28101
rect 35060 28135 35118 28141
rect 35060 28101 35072 28135
rect 35106 28132 35118 28135
rect 36170 28132 36176 28144
rect 35106 28104 36176 28132
rect 35106 28101 35118 28104
rect 35060 28095 35118 28101
rect 36170 28092 36176 28104
rect 36228 28092 36234 28144
rect 38654 28132 38660 28144
rect 38615 28104 38660 28132
rect 38654 28092 38660 28104
rect 38712 28132 38718 28144
rect 42058 28132 42064 28144
rect 38712 28104 42064 28132
rect 38712 28092 38718 28104
rect 42058 28092 42064 28104
rect 42116 28092 42122 28144
rect 44076 28135 44134 28141
rect 44076 28101 44088 28135
rect 44122 28132 44134 28135
rect 45186 28132 45192 28144
rect 44122 28104 45192 28132
rect 44122 28101 44134 28104
rect 44076 28095 44134 28101
rect 45186 28092 45192 28104
rect 45244 28092 45250 28144
rect 45916 28135 45974 28141
rect 45916 28101 45928 28135
rect 45962 28132 45974 28135
rect 47118 28132 47124 28144
rect 45962 28104 47124 28132
rect 45962 28101 45974 28104
rect 45916 28095 45974 28101
rect 47118 28092 47124 28104
rect 47176 28092 47182 28144
rect 48314 28132 48320 28144
rect 47688 28104 48320 28132
rect 28810 28064 28816 28076
rect 28276 28036 28816 28064
rect 28810 28024 28816 28036
rect 28868 28064 28874 28076
rect 32125 28067 32183 28073
rect 32125 28064 32137 28067
rect 28868 28036 32137 28064
rect 28868 28024 28874 28036
rect 32125 28033 32137 28036
rect 32171 28033 32183 28067
rect 32125 28027 32183 28033
rect 32392 28067 32450 28073
rect 32392 28033 32404 28067
rect 32438 28064 32450 28067
rect 32674 28064 32680 28076
rect 32438 28036 32680 28064
rect 32438 28033 32450 28036
rect 32392 28027 32450 28033
rect 32674 28024 32680 28036
rect 32732 28024 32738 28076
rect 43809 28067 43867 28073
rect 43809 28033 43821 28067
rect 43855 28064 43867 28067
rect 44358 28064 44364 28076
rect 43855 28036 44364 28064
rect 43855 28033 43867 28036
rect 43809 28027 43867 28033
rect 44358 28024 44364 28036
rect 44416 28024 44422 28076
rect 45646 28064 45652 28076
rect 45607 28036 45652 28064
rect 45646 28024 45652 28036
rect 45704 28024 45710 28076
rect 47688 28073 47716 28104
rect 48314 28092 48320 28104
rect 48372 28132 48378 28144
rect 49418 28132 49424 28144
rect 48372 28104 49424 28132
rect 48372 28092 48378 28104
rect 49418 28092 49424 28104
rect 49476 28092 49482 28144
rect 49786 28141 49792 28144
rect 49780 28132 49792 28141
rect 49747 28104 49792 28132
rect 49780 28095 49792 28104
rect 49786 28092 49792 28095
rect 49844 28092 49850 28144
rect 57054 28132 57060 28144
rect 55968 28104 57060 28132
rect 47673 28067 47731 28073
rect 47673 28033 47685 28067
rect 47719 28033 47731 28067
rect 47673 28027 47731 28033
rect 47940 28067 47998 28073
rect 47940 28033 47952 28067
rect 47986 28064 47998 28067
rect 48958 28064 48964 28076
rect 47986 28036 48964 28064
rect 47986 28033 47998 28036
rect 47940 28027 47998 28033
rect 48958 28024 48964 28036
rect 49016 28024 49022 28076
rect 53190 28024 53196 28076
rect 53248 28064 53254 28076
rect 53377 28067 53435 28073
rect 53377 28064 53389 28067
rect 53248 28036 53389 28064
rect 53248 28024 53254 28036
rect 53377 28033 53389 28036
rect 53423 28033 53435 28067
rect 53377 28027 53435 28033
rect 53644 28067 53702 28073
rect 53644 28033 53656 28067
rect 53690 28064 53702 28067
rect 54754 28064 54760 28076
rect 53690 28036 54760 28064
rect 53690 28033 53702 28036
rect 53644 28027 53702 28033
rect 54754 28024 54760 28036
rect 54812 28024 54818 28076
rect 55968 28073 55996 28104
rect 57054 28092 57060 28104
rect 57112 28092 57118 28144
rect 55953 28067 56011 28073
rect 55953 28033 55965 28067
rect 55999 28033 56011 28067
rect 55953 28027 56011 28033
rect 56220 28067 56278 28073
rect 56220 28033 56232 28067
rect 56266 28064 56278 28067
rect 57238 28064 57244 28076
rect 56266 28036 57244 28064
rect 56266 28033 56278 28036
rect 56220 28027 56278 28033
rect 57238 28024 57244 28036
rect 57296 28024 57302 28076
rect 9582 27996 9588 28008
rect 9543 27968 9588 27996
rect 9582 27956 9588 27968
rect 9640 27956 9646 28008
rect 16666 27956 16672 28008
rect 16724 27996 16730 28008
rect 17037 27999 17095 28005
rect 17037 27996 17049 27999
rect 16724 27968 17049 27996
rect 16724 27956 16730 27968
rect 17037 27965 17049 27968
rect 17083 27965 17095 27999
rect 17037 27959 17095 27965
rect 22462 27956 22468 28008
rect 22520 27996 22526 28008
rect 22741 27999 22799 28005
rect 22741 27996 22753 27999
rect 22520 27968 22753 27996
rect 22520 27956 22526 27968
rect 22741 27965 22753 27968
rect 22787 27965 22799 27999
rect 22741 27959 22799 27965
rect 34698 27956 34704 28008
rect 34756 27996 34762 28008
rect 34793 27999 34851 28005
rect 34793 27996 34805 27999
rect 34756 27968 34805 27996
rect 34756 27956 34762 27968
rect 34793 27965 34805 27968
rect 34839 27965 34851 27999
rect 34793 27959 34851 27965
rect 49418 27956 49424 28008
rect 49476 27996 49482 28008
rect 49513 27999 49571 28005
rect 49513 27996 49525 27999
rect 49476 27968 49525 27996
rect 49476 27956 49482 27968
rect 49513 27965 49525 27968
rect 49559 27965 49571 27999
rect 49513 27959 49571 27965
rect 28074 27888 28080 27940
rect 28132 27928 28138 27940
rect 28353 27931 28411 27937
rect 28353 27928 28365 27931
rect 28132 27900 28365 27928
rect 28132 27888 28138 27900
rect 28353 27897 28365 27900
rect 28399 27897 28411 27931
rect 28353 27891 28411 27897
rect 45094 27888 45100 27940
rect 45152 27928 45158 27940
rect 45189 27931 45247 27937
rect 45189 27928 45201 27931
rect 45152 27900 45201 27928
rect 45152 27888 45158 27900
rect 45189 27897 45201 27900
rect 45235 27897 45247 27931
rect 45189 27891 45247 27897
rect 14090 27860 14096 27872
rect 14051 27832 14096 27860
rect 14090 27820 14096 27832
rect 14148 27820 14154 27872
rect 16114 27860 16120 27872
rect 16075 27832 16120 27860
rect 16114 27820 16120 27832
rect 16172 27820 16178 27872
rect 18414 27860 18420 27872
rect 18375 27832 18420 27860
rect 18414 27820 18420 27832
rect 18472 27820 18478 27872
rect 20622 27860 20628 27872
rect 20583 27832 20628 27860
rect 20622 27820 20628 27832
rect 20680 27820 20686 27872
rect 24118 27860 24124 27872
rect 24079 27832 24124 27860
rect 24118 27820 24124 27832
rect 24176 27820 24182 27872
rect 25866 27820 25872 27872
rect 25924 27860 25930 27872
rect 29546 27860 29552 27872
rect 25924 27832 29552 27860
rect 25924 27820 25930 27832
rect 29546 27820 29552 27832
rect 29604 27820 29610 27872
rect 33502 27860 33508 27872
rect 33463 27832 33508 27860
rect 33502 27820 33508 27832
rect 33560 27820 33566 27872
rect 36170 27860 36176 27872
rect 36131 27832 36176 27860
rect 36170 27820 36176 27832
rect 36228 27820 36234 27872
rect 56594 27820 56600 27872
rect 56652 27860 56658 27872
rect 57333 27863 57391 27869
rect 57333 27860 57345 27863
rect 56652 27832 57345 27860
rect 56652 27820 56658 27832
rect 57333 27829 57345 27832
rect 57379 27829 57391 27863
rect 57333 27823 57391 27829
rect 1104 27770 59340 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 59340 27770
rect 1104 27696 59340 27718
rect 8202 27588 8208 27600
rect 8163 27560 8208 27588
rect 8202 27548 8208 27560
rect 8260 27548 8266 27600
rect 13538 27588 13544 27600
rect 13499 27560 13544 27588
rect 13538 27548 13544 27560
rect 13596 27548 13602 27600
rect 16390 27588 16396 27600
rect 16351 27560 16396 27588
rect 16390 27548 16396 27560
rect 16448 27548 16454 27600
rect 20530 27548 20536 27600
rect 20588 27588 20594 27600
rect 20625 27591 20683 27597
rect 20625 27588 20637 27591
rect 20588 27560 20637 27588
rect 20588 27548 20594 27560
rect 20625 27557 20637 27560
rect 20671 27557 20683 27591
rect 20625 27551 20683 27557
rect 28166 27548 28172 27600
rect 28224 27588 28230 27600
rect 28353 27591 28411 27597
rect 28353 27588 28365 27591
rect 28224 27560 28365 27588
rect 28224 27548 28230 27560
rect 28353 27557 28365 27560
rect 28399 27557 28411 27591
rect 41874 27588 41880 27600
rect 41835 27560 41880 27588
rect 28353 27551 28411 27557
rect 41874 27548 41880 27560
rect 41932 27548 41938 27600
rect 44266 27548 44272 27600
rect 44324 27588 44330 27600
rect 44453 27591 44511 27597
rect 44453 27588 44465 27591
rect 44324 27560 44465 27588
rect 44324 27548 44330 27560
rect 44453 27557 44465 27560
rect 44499 27557 44511 27591
rect 54754 27588 54760 27600
rect 54715 27560 54760 27588
rect 44453 27551 44511 27557
rect 54754 27548 54760 27560
rect 54812 27548 54818 27600
rect 19242 27520 19248 27532
rect 19203 27492 19248 27520
rect 19242 27480 19248 27492
rect 19300 27480 19306 27532
rect 39942 27480 39948 27532
rect 40000 27520 40006 27532
rect 40497 27523 40555 27529
rect 40497 27520 40509 27523
rect 40000 27492 40509 27520
rect 40000 27480 40006 27492
rect 40497 27489 40509 27492
rect 40543 27489 40555 27523
rect 40497 27483 40555 27489
rect 42978 27480 42984 27532
rect 43036 27520 43042 27532
rect 43073 27523 43131 27529
rect 43073 27520 43085 27523
rect 43036 27492 43085 27520
rect 43036 27480 43042 27492
rect 43073 27489 43085 27492
rect 43119 27489 43131 27523
rect 50154 27520 50160 27532
rect 50115 27492 50160 27520
rect 43073 27483 43131 27489
rect 50154 27480 50160 27492
rect 50212 27480 50218 27532
rect 6825 27455 6883 27461
rect 6825 27421 6837 27455
rect 6871 27452 6883 27455
rect 6914 27452 6920 27464
rect 6871 27424 6920 27452
rect 6871 27421 6883 27424
rect 6825 27415 6883 27421
rect 6914 27412 6920 27424
rect 6972 27412 6978 27464
rect 7098 27461 7104 27464
rect 7092 27452 7104 27461
rect 7059 27424 7104 27452
rect 7092 27415 7104 27424
rect 7098 27412 7104 27415
rect 7156 27412 7162 27464
rect 12161 27455 12219 27461
rect 12161 27421 12173 27455
rect 12207 27452 12219 27455
rect 12250 27452 12256 27464
rect 12207 27424 12256 27452
rect 12207 27421 12219 27424
rect 12161 27415 12219 27421
rect 12250 27412 12256 27424
rect 12308 27412 12314 27464
rect 12428 27455 12486 27461
rect 12428 27421 12440 27455
rect 12474 27452 12486 27455
rect 14090 27452 14096 27464
rect 12474 27424 14096 27452
rect 12474 27421 12486 27424
rect 12428 27415 12486 27421
rect 14090 27412 14096 27424
rect 14148 27412 14154 27464
rect 14734 27412 14740 27464
rect 14792 27452 14798 27464
rect 15013 27455 15071 27461
rect 15013 27452 15025 27455
rect 14792 27424 15025 27452
rect 14792 27412 14798 27424
rect 15013 27421 15025 27424
rect 15059 27421 15071 27455
rect 15013 27415 15071 27421
rect 15280 27455 15338 27461
rect 15280 27421 15292 27455
rect 15326 27452 15338 27455
rect 16114 27452 16120 27464
rect 15326 27424 16120 27452
rect 15326 27421 15338 27424
rect 15280 27415 15338 27421
rect 16114 27412 16120 27424
rect 16172 27412 16178 27464
rect 16666 27412 16672 27464
rect 16724 27452 16730 27464
rect 16853 27455 16911 27461
rect 16853 27452 16865 27455
rect 16724 27424 16865 27452
rect 16724 27412 16730 27424
rect 16853 27421 16865 27424
rect 16899 27421 16911 27455
rect 16853 27415 16911 27421
rect 17120 27455 17178 27461
rect 17120 27421 17132 27455
rect 17166 27452 17178 27455
rect 18414 27452 18420 27464
rect 17166 27424 18420 27452
rect 17166 27421 17178 27424
rect 17120 27415 17178 27421
rect 18414 27412 18420 27424
rect 18472 27412 18478 27464
rect 19512 27455 19570 27461
rect 19512 27421 19524 27455
rect 19558 27452 19570 27455
rect 20622 27452 20628 27464
rect 19558 27424 20628 27452
rect 19558 27421 19570 27424
rect 19512 27415 19570 27421
rect 20622 27412 20628 27424
rect 20680 27412 20686 27464
rect 22462 27452 22468 27464
rect 22423 27424 22468 27452
rect 22462 27412 22468 27424
rect 22520 27412 22526 27464
rect 22732 27455 22790 27461
rect 22732 27421 22744 27455
rect 22778 27452 22790 27455
rect 24118 27452 24124 27464
rect 22778 27424 24124 27452
rect 22778 27421 22790 27424
rect 22732 27415 22790 27421
rect 24118 27412 24124 27424
rect 24176 27412 24182 27464
rect 24397 27455 24455 27461
rect 24397 27421 24409 27455
rect 24443 27421 24455 27455
rect 24397 27415 24455 27421
rect 23382 27344 23388 27396
rect 23440 27384 23446 27396
rect 24412 27384 24440 27415
rect 25130 27412 25136 27464
rect 25188 27452 25194 27464
rect 26973 27455 27031 27461
rect 26973 27452 26985 27455
rect 25188 27424 26985 27452
rect 25188 27412 25194 27424
rect 26973 27421 26985 27424
rect 27019 27452 27031 27455
rect 27614 27452 27620 27464
rect 27019 27424 27620 27452
rect 27019 27421 27031 27424
rect 26973 27415 27031 27421
rect 27614 27412 27620 27424
rect 27672 27412 27678 27464
rect 29549 27455 29607 27461
rect 29549 27421 29561 27455
rect 29595 27452 29607 27455
rect 30098 27452 30104 27464
rect 29595 27424 30104 27452
rect 29595 27421 29607 27424
rect 29549 27415 29607 27421
rect 30098 27412 30104 27424
rect 30156 27452 30162 27464
rect 31389 27455 31447 27461
rect 31389 27452 31401 27455
rect 30156 27424 31401 27452
rect 30156 27412 30162 27424
rect 31389 27421 31401 27424
rect 31435 27421 31447 27455
rect 31389 27415 31447 27421
rect 31478 27412 31484 27464
rect 31536 27452 31542 27464
rect 31645 27455 31703 27461
rect 31645 27452 31657 27455
rect 31536 27424 31657 27452
rect 31536 27412 31542 27424
rect 31645 27421 31657 27424
rect 31691 27421 31703 27455
rect 34698 27452 34704 27464
rect 34659 27424 34704 27452
rect 31645 27415 31703 27421
rect 34698 27412 34704 27424
rect 34756 27412 34762 27464
rect 34968 27455 35026 27461
rect 34968 27421 34980 27455
rect 35014 27452 35026 27455
rect 36170 27452 36176 27464
rect 35014 27424 36176 27452
rect 35014 27421 35026 27424
rect 34968 27415 35026 27421
rect 36170 27412 36176 27424
rect 36228 27412 36234 27464
rect 37274 27452 37280 27464
rect 37235 27424 37280 27452
rect 37274 27412 37280 27424
rect 37332 27412 37338 27464
rect 40764 27455 40822 27461
rect 40764 27421 40776 27455
rect 40810 27452 40822 27455
rect 41046 27452 41052 27464
rect 40810 27424 41052 27452
rect 40810 27421 40822 27424
rect 40764 27415 40822 27421
rect 41046 27412 41052 27424
rect 41104 27412 41110 27464
rect 43340 27455 43398 27461
rect 43340 27421 43352 27455
rect 43386 27452 43398 27455
rect 44174 27452 44180 27464
rect 43386 27424 44180 27452
rect 43386 27421 43398 27424
rect 43340 27415 43398 27421
rect 44174 27412 44180 27424
rect 44232 27412 44238 27464
rect 44358 27412 44364 27464
rect 44416 27452 44422 27464
rect 45005 27455 45063 27461
rect 45005 27452 45017 27455
rect 44416 27424 45017 27452
rect 44416 27412 44422 27424
rect 45005 27421 45017 27424
rect 45051 27452 45063 27455
rect 46845 27455 46903 27461
rect 46845 27452 46857 27455
rect 45051 27424 46857 27452
rect 45051 27421 45063 27424
rect 45005 27415 45063 27421
rect 46845 27421 46857 27424
rect 46891 27421 46903 27455
rect 46845 27415 46903 27421
rect 53377 27455 53435 27461
rect 53377 27421 53389 27455
rect 53423 27452 53435 27455
rect 54110 27452 54116 27464
rect 53423 27424 54116 27452
rect 53423 27421 53435 27424
rect 53377 27415 53435 27421
rect 54110 27412 54116 27424
rect 54168 27412 54174 27464
rect 56505 27455 56563 27461
rect 56505 27421 56517 27455
rect 56551 27452 56563 27455
rect 57054 27452 57060 27464
rect 56551 27424 57060 27452
rect 56551 27421 56563 27424
rect 56505 27415 56563 27421
rect 57054 27412 57060 27424
rect 57112 27412 57118 27464
rect 23440 27356 24440 27384
rect 24664 27387 24722 27393
rect 23440 27344 23446 27356
rect 24664 27353 24676 27387
rect 24710 27384 24722 27387
rect 25314 27384 25320 27396
rect 24710 27356 25320 27384
rect 24710 27353 24722 27356
rect 24664 27347 24722 27353
rect 25314 27344 25320 27356
rect 25372 27344 25378 27396
rect 27240 27387 27298 27393
rect 27240 27353 27252 27387
rect 27286 27384 27298 27387
rect 28994 27384 29000 27396
rect 27286 27356 29000 27384
rect 27286 27353 27298 27356
rect 27240 27347 27298 27353
rect 28994 27344 29000 27356
rect 29052 27344 29058 27396
rect 29816 27387 29874 27393
rect 29816 27353 29828 27387
rect 29862 27384 29874 27387
rect 32582 27384 32588 27396
rect 29862 27356 32588 27384
rect 29862 27353 29874 27356
rect 29816 27347 29874 27353
rect 32582 27344 32588 27356
rect 32640 27344 32646 27396
rect 37544 27387 37602 27393
rect 37544 27353 37556 27387
rect 37590 27384 37602 27387
rect 40402 27384 40408 27396
rect 37590 27356 40408 27384
rect 37590 27353 37602 27356
rect 37544 27347 37602 27353
rect 40402 27344 40408 27356
rect 40460 27344 40466 27396
rect 45272 27387 45330 27393
rect 45272 27353 45284 27387
rect 45318 27384 45330 27387
rect 45646 27384 45652 27396
rect 45318 27356 45652 27384
rect 45318 27353 45330 27356
rect 45272 27347 45330 27353
rect 45646 27344 45652 27356
rect 45704 27344 45710 27396
rect 47112 27387 47170 27393
rect 47112 27353 47124 27387
rect 47158 27384 47170 27387
rect 48130 27384 48136 27396
rect 47158 27356 48136 27384
rect 47158 27353 47170 27356
rect 47112 27347 47170 27353
rect 48130 27344 48136 27356
rect 48188 27344 48194 27396
rect 50424 27387 50482 27393
rect 50424 27353 50436 27387
rect 50470 27384 50482 27387
rect 50798 27384 50804 27396
rect 50470 27356 50804 27384
rect 50470 27353 50482 27356
rect 50424 27347 50482 27353
rect 50798 27344 50804 27356
rect 50856 27344 50862 27396
rect 53644 27387 53702 27393
rect 53644 27353 53656 27387
rect 53690 27384 53702 27387
rect 54662 27384 54668 27396
rect 53690 27356 54668 27384
rect 53690 27353 53702 27356
rect 53644 27347 53702 27353
rect 54662 27344 54668 27356
rect 54720 27344 54726 27396
rect 56772 27387 56830 27393
rect 56772 27353 56784 27387
rect 56818 27384 56830 27387
rect 57330 27384 57336 27396
rect 56818 27356 57336 27384
rect 56818 27353 56830 27356
rect 56772 27347 56830 27353
rect 57330 27344 57336 27356
rect 57388 27344 57394 27396
rect 18230 27316 18236 27328
rect 18191 27288 18236 27316
rect 18230 27276 18236 27288
rect 18288 27276 18294 27328
rect 23842 27316 23848 27328
rect 23803 27288 23848 27316
rect 23842 27276 23848 27288
rect 23900 27276 23906 27328
rect 24486 27276 24492 27328
rect 24544 27316 24550 27328
rect 25777 27319 25835 27325
rect 25777 27316 25789 27319
rect 24544 27288 25789 27316
rect 24544 27276 24550 27288
rect 25777 27285 25789 27288
rect 25823 27285 25835 27319
rect 25777 27279 25835 27285
rect 27890 27276 27896 27328
rect 27948 27316 27954 27328
rect 30929 27319 30987 27325
rect 30929 27316 30941 27319
rect 27948 27288 30941 27316
rect 27948 27276 27954 27288
rect 30929 27285 30941 27288
rect 30975 27285 30987 27319
rect 32766 27316 32772 27328
rect 32727 27288 32772 27316
rect 30929 27279 30987 27285
rect 32766 27276 32772 27288
rect 32824 27276 32830 27328
rect 36078 27316 36084 27328
rect 36039 27288 36084 27316
rect 36078 27276 36084 27288
rect 36136 27276 36142 27328
rect 38657 27319 38715 27325
rect 38657 27285 38669 27319
rect 38703 27316 38715 27319
rect 39298 27316 39304 27328
rect 38703 27288 39304 27316
rect 38703 27285 38715 27288
rect 38657 27279 38715 27285
rect 39298 27276 39304 27288
rect 39356 27276 39362 27328
rect 46385 27319 46443 27325
rect 46385 27285 46397 27319
rect 46431 27316 46443 27319
rect 46934 27316 46940 27328
rect 46431 27288 46940 27316
rect 46431 27285 46443 27288
rect 46385 27279 46443 27285
rect 46934 27276 46940 27288
rect 46992 27276 46998 27328
rect 48222 27316 48228 27328
rect 48183 27288 48228 27316
rect 48222 27276 48228 27288
rect 48280 27276 48286 27328
rect 51534 27316 51540 27328
rect 51495 27288 51540 27316
rect 51534 27276 51540 27288
rect 51592 27276 51598 27328
rect 57882 27316 57888 27328
rect 57843 27288 57888 27316
rect 57882 27276 57888 27288
rect 57940 27276 57946 27328
rect 1104 27226 59340 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 59340 27226
rect 1104 27152 59340 27174
rect 18046 27112 18052 27124
rect 18007 27084 18052 27112
rect 18046 27072 18052 27084
rect 18104 27072 18110 27124
rect 23474 27112 23480 27124
rect 23435 27084 23480 27112
rect 23474 27072 23480 27084
rect 23532 27072 23538 27124
rect 25314 27112 25320 27124
rect 25275 27084 25320 27112
rect 25314 27072 25320 27084
rect 25372 27072 25378 27124
rect 45646 27112 45652 27124
rect 45607 27084 45652 27112
rect 45646 27072 45652 27084
rect 45704 27072 45710 27124
rect 48958 27112 48964 27124
rect 48919 27084 48964 27112
rect 48958 27072 48964 27084
rect 49016 27072 49022 27124
rect 50798 27112 50804 27124
rect 50759 27084 50804 27112
rect 50798 27072 50804 27084
rect 50856 27072 50862 27124
rect 54662 27072 54668 27124
rect 54720 27112 54726 27124
rect 54757 27115 54815 27121
rect 54757 27112 54769 27115
rect 54720 27084 54769 27112
rect 54720 27072 54726 27084
rect 54757 27081 54769 27084
rect 54803 27081 54815 27115
rect 54757 27075 54815 27081
rect 57238 27072 57244 27124
rect 57296 27112 57302 27124
rect 57333 27115 57391 27121
rect 57333 27112 57345 27115
rect 57296 27084 57345 27112
rect 57296 27072 57302 27084
rect 57333 27081 57345 27084
rect 57379 27081 57391 27115
rect 57333 27075 57391 27081
rect 12250 27044 12256 27056
rect 11532 27016 12256 27044
rect 6914 26936 6920 26988
rect 6972 26976 6978 26988
rect 7653 26979 7711 26985
rect 7653 26976 7665 26979
rect 6972 26948 7665 26976
rect 6972 26936 6978 26948
rect 7653 26945 7665 26948
rect 7699 26945 7711 26979
rect 7653 26939 7711 26945
rect 7920 26979 7978 26985
rect 7920 26945 7932 26979
rect 7966 26976 7978 26979
rect 8478 26976 8484 26988
rect 7966 26948 8484 26976
rect 7966 26945 7978 26948
rect 7920 26939 7978 26945
rect 8478 26936 8484 26948
rect 8536 26936 8542 26988
rect 11532 26985 11560 27016
rect 12250 27004 12256 27016
rect 12308 27004 12314 27056
rect 12526 27004 12532 27056
rect 12584 27044 12590 27056
rect 13541 27047 13599 27053
rect 13541 27044 13553 27047
rect 12584 27016 13553 27044
rect 12584 27004 12590 27016
rect 13541 27013 13553 27016
rect 13587 27013 13599 27047
rect 13541 27007 13599 27013
rect 16936 27047 16994 27053
rect 16936 27013 16948 27047
rect 16982 27044 16994 27047
rect 18230 27044 18236 27056
rect 16982 27016 18236 27044
rect 16982 27013 16994 27016
rect 16936 27007 16994 27013
rect 18230 27004 18236 27016
rect 18288 27004 18294 27056
rect 22364 27047 22422 27053
rect 22364 27013 22376 27047
rect 22410 27044 22422 27047
rect 23842 27044 23848 27056
rect 22410 27016 23848 27044
rect 22410 27013 22422 27016
rect 22364 27007 22422 27013
rect 23842 27004 23848 27016
rect 23900 27004 23906 27056
rect 24762 27004 24768 27056
rect 24820 27044 24826 27056
rect 32760 27047 32818 27053
rect 24820 27016 27844 27044
rect 24820 27004 24826 27016
rect 27816 26988 27844 27016
rect 32760 27013 32772 27047
rect 32806 27044 32818 27047
rect 33502 27044 33508 27056
rect 32806 27016 33508 27044
rect 32806 27013 32818 27016
rect 32760 27007 32818 27013
rect 33502 27004 33508 27016
rect 33560 27004 33566 27056
rect 34968 27047 35026 27053
rect 34968 27013 34980 27047
rect 35014 27044 35026 27047
rect 36078 27044 36084 27056
rect 35014 27016 36084 27044
rect 35014 27013 35026 27016
rect 34968 27007 35026 27013
rect 36078 27004 36084 27016
rect 36136 27004 36142 27056
rect 37274 27004 37280 27056
rect 37332 27044 37338 27056
rect 39942 27044 39948 27056
rect 37332 27016 39948 27044
rect 37332 27004 37338 27016
rect 11790 26985 11796 26988
rect 11517 26979 11575 26985
rect 11517 26945 11529 26979
rect 11563 26945 11575 26979
rect 11517 26939 11575 26945
rect 11784 26939 11796 26985
rect 11848 26976 11854 26988
rect 11848 26948 11884 26976
rect 11790 26936 11796 26939
rect 11848 26936 11854 26948
rect 13630 26936 13636 26988
rect 13688 26976 13694 26988
rect 17954 26976 17960 26988
rect 13688 26948 17960 26976
rect 13688 26936 13694 26948
rect 17954 26936 17960 26948
rect 18012 26936 18018 26988
rect 19242 26936 19248 26988
rect 19300 26976 19306 26988
rect 19889 26979 19947 26985
rect 19889 26976 19901 26979
rect 19300 26948 19901 26976
rect 19300 26936 19306 26948
rect 19889 26945 19901 26948
rect 19935 26945 19947 26979
rect 19889 26939 19947 26945
rect 20156 26979 20214 26985
rect 20156 26945 20168 26979
rect 20202 26976 20214 26979
rect 23106 26976 23112 26988
rect 20202 26948 23112 26976
rect 20202 26945 20214 26948
rect 20156 26939 20214 26945
rect 16666 26908 16672 26920
rect 16627 26880 16672 26908
rect 16666 26868 16672 26880
rect 16724 26868 16730 26920
rect 9030 26772 9036 26784
rect 8991 26744 9036 26772
rect 9030 26732 9036 26744
rect 9088 26732 9094 26784
rect 9122 26732 9128 26784
rect 9180 26772 9186 26784
rect 12897 26775 12955 26781
rect 12897 26772 12909 26775
rect 9180 26744 12909 26772
rect 9180 26732 9186 26744
rect 12897 26741 12909 26744
rect 12943 26741 12955 26775
rect 12897 26735 12955 26741
rect 15013 26775 15071 26781
rect 15013 26741 15025 26775
rect 15059 26772 15071 26775
rect 15102 26772 15108 26784
rect 15059 26744 15108 26772
rect 15059 26741 15071 26744
rect 15013 26735 15071 26741
rect 15102 26732 15108 26744
rect 15160 26732 15166 26784
rect 19904 26772 19932 26939
rect 23106 26936 23112 26948
rect 23164 26936 23170 26988
rect 24204 26979 24262 26985
rect 24204 26945 24216 26979
rect 24250 26976 24262 26979
rect 25774 26976 25780 26988
rect 24250 26948 25780 26976
rect 24250 26945 24262 26948
rect 24204 26939 24262 26945
rect 25774 26936 25780 26948
rect 25832 26936 25838 26988
rect 27798 26936 27804 26988
rect 27856 26976 27862 26988
rect 28721 26979 28779 26985
rect 28721 26976 28733 26979
rect 27856 26948 28733 26976
rect 27856 26936 27862 26948
rect 28721 26945 28733 26948
rect 28767 26945 28779 26979
rect 28721 26939 28779 26945
rect 30098 26936 30104 26988
rect 30156 26976 30162 26988
rect 32493 26979 32551 26985
rect 32493 26976 32505 26979
rect 30156 26948 32505 26976
rect 30156 26936 30162 26948
rect 32493 26945 32505 26948
rect 32539 26976 32551 26979
rect 33134 26976 33140 26988
rect 32539 26948 33140 26976
rect 32539 26945 32551 26948
rect 32493 26939 32551 26945
rect 33134 26936 33140 26948
rect 33192 26936 33198 26988
rect 34698 26976 34704 26988
rect 34611 26948 34704 26976
rect 34698 26936 34704 26948
rect 34756 26976 34762 26988
rect 35710 26976 35716 26988
rect 34756 26948 35716 26976
rect 34756 26936 34762 26948
rect 35710 26936 35716 26948
rect 35768 26936 35774 26988
rect 37660 26985 37688 27016
rect 37645 26979 37703 26985
rect 37645 26945 37657 26979
rect 37691 26945 37703 26979
rect 37645 26939 37703 26945
rect 37912 26979 37970 26985
rect 37912 26945 37924 26979
rect 37958 26976 37970 26979
rect 38654 26976 38660 26988
rect 37958 26948 38660 26976
rect 37958 26945 37970 26948
rect 37912 26939 37970 26945
rect 38654 26936 38660 26948
rect 38712 26936 38718 26988
rect 39500 26985 39528 27016
rect 39942 27004 39948 27016
rect 40000 27004 40006 27056
rect 42696 27047 42754 27053
rect 42696 27013 42708 27047
rect 42742 27044 42754 27047
rect 46290 27044 46296 27056
rect 42742 27016 46296 27044
rect 42742 27013 42754 27016
rect 42696 27007 42754 27013
rect 46290 27004 46296 27016
rect 46348 27004 46354 27056
rect 47848 27047 47906 27053
rect 47848 27013 47860 27047
rect 47894 27044 47906 27047
rect 48222 27044 48228 27056
rect 47894 27016 48228 27044
rect 47894 27013 47906 27016
rect 47848 27007 47906 27013
rect 48222 27004 48228 27016
rect 48280 27004 48286 27056
rect 49688 27047 49746 27053
rect 49688 27013 49700 27047
rect 49734 27044 49746 27047
rect 50706 27044 50712 27056
rect 49734 27016 50712 27044
rect 49734 27013 49746 27016
rect 49688 27007 49746 27013
rect 50706 27004 50712 27016
rect 50764 27004 50770 27056
rect 56220 27047 56278 27053
rect 56220 27013 56232 27047
rect 56266 27044 56278 27047
rect 57882 27044 57888 27056
rect 56266 27016 57888 27044
rect 56266 27013 56278 27016
rect 56220 27007 56278 27013
rect 57882 27004 57888 27016
rect 57940 27004 57946 27056
rect 39485 26979 39543 26985
rect 39485 26945 39497 26979
rect 39531 26945 39543 26979
rect 39485 26939 39543 26945
rect 39752 26979 39810 26985
rect 39752 26945 39764 26979
rect 39798 26976 39810 26979
rect 41230 26976 41236 26988
rect 39798 26948 41236 26976
rect 39798 26945 39810 26948
rect 39752 26939 39810 26945
rect 41230 26936 41236 26948
rect 41288 26936 41294 26988
rect 42429 26979 42487 26985
rect 42429 26945 42441 26979
rect 42475 26976 42487 26979
rect 42518 26976 42524 26988
rect 42475 26948 42524 26976
rect 42475 26945 42487 26948
rect 42429 26939 42487 26945
rect 42518 26936 42524 26948
rect 42576 26936 42582 26988
rect 44269 26979 44327 26985
rect 44269 26945 44281 26979
rect 44315 26976 44327 26979
rect 44358 26976 44364 26988
rect 44315 26948 44364 26976
rect 44315 26945 44327 26948
rect 44269 26939 44327 26945
rect 44358 26936 44364 26948
rect 44416 26936 44422 26988
rect 44536 26979 44594 26985
rect 44536 26945 44548 26979
rect 44582 26976 44594 26979
rect 46382 26976 46388 26988
rect 44582 26948 46388 26976
rect 44582 26945 44594 26948
rect 44536 26939 44594 26945
rect 46382 26936 46388 26948
rect 46440 26936 46446 26988
rect 49418 26976 49424 26988
rect 49379 26948 49424 26976
rect 49418 26936 49424 26948
rect 49476 26936 49482 26988
rect 53190 26936 53196 26988
rect 53248 26976 53254 26988
rect 53377 26979 53435 26985
rect 53377 26976 53389 26979
rect 53248 26948 53389 26976
rect 53248 26936 53254 26948
rect 53377 26945 53389 26948
rect 53423 26945 53435 26979
rect 53377 26939 53435 26945
rect 53644 26979 53702 26985
rect 53644 26945 53656 26979
rect 53690 26976 53702 26979
rect 54754 26976 54760 26988
rect 53690 26948 54760 26976
rect 53690 26945 53702 26948
rect 53644 26939 53702 26945
rect 54754 26936 54760 26948
rect 54812 26936 54818 26988
rect 55953 26979 56011 26985
rect 55953 26945 55965 26979
rect 55999 26976 56011 26979
rect 57054 26976 57060 26988
rect 55999 26948 57060 26976
rect 55999 26945 56011 26948
rect 55953 26939 56011 26945
rect 57054 26936 57060 26948
rect 57112 26936 57118 26988
rect 22097 26911 22155 26917
rect 22097 26908 22109 26911
rect 20916 26880 22109 26908
rect 20916 26772 20944 26880
rect 22097 26877 22109 26880
rect 22143 26877 22155 26911
rect 22097 26871 22155 26877
rect 23382 26868 23388 26920
rect 23440 26908 23446 26920
rect 23937 26911 23995 26917
rect 23937 26908 23949 26911
rect 23440 26880 23949 26908
rect 23440 26868 23446 26880
rect 23937 26877 23949 26880
rect 23983 26877 23995 26911
rect 23937 26871 23995 26877
rect 46842 26868 46848 26920
rect 46900 26908 46906 26920
rect 47581 26911 47639 26917
rect 47581 26908 47593 26911
rect 46900 26880 47593 26908
rect 46900 26868 46906 26880
rect 47581 26877 47593 26880
rect 47627 26877 47639 26911
rect 47581 26871 47639 26877
rect 35986 26800 35992 26852
rect 36044 26840 36050 26852
rect 36081 26843 36139 26849
rect 36081 26840 36093 26843
rect 36044 26812 36093 26840
rect 36044 26800 36050 26812
rect 36081 26809 36093 26812
rect 36127 26809 36139 26843
rect 36081 26803 36139 26809
rect 21266 26772 21272 26784
rect 19904 26744 20944 26772
rect 21227 26744 21272 26772
rect 21266 26732 21272 26744
rect 21324 26732 21330 26784
rect 30190 26772 30196 26784
rect 30151 26744 30196 26772
rect 30190 26732 30196 26744
rect 30248 26732 30254 26784
rect 32398 26732 32404 26784
rect 32456 26772 32462 26784
rect 33873 26775 33931 26781
rect 33873 26772 33885 26775
rect 32456 26744 33885 26772
rect 32456 26732 32462 26744
rect 33873 26741 33885 26744
rect 33919 26741 33931 26775
rect 39022 26772 39028 26784
rect 38983 26744 39028 26772
rect 33873 26735 33931 26741
rect 39022 26732 39028 26744
rect 39080 26732 39086 26784
rect 40865 26775 40923 26781
rect 40865 26741 40877 26775
rect 40911 26772 40923 26775
rect 41782 26772 41788 26784
rect 40911 26744 41788 26772
rect 40911 26741 40923 26744
rect 40865 26735 40923 26741
rect 41782 26732 41788 26744
rect 41840 26732 41846 26784
rect 43809 26775 43867 26781
rect 43809 26741 43821 26775
rect 43855 26772 43867 26775
rect 44450 26772 44456 26784
rect 43855 26744 44456 26772
rect 43855 26741 43867 26744
rect 43809 26735 43867 26741
rect 44450 26732 44456 26744
rect 44508 26732 44514 26784
rect 1104 26682 59340 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 59340 26682
rect 1104 26608 59340 26630
rect 6914 26568 6920 26580
rect 6656 26540 6920 26568
rect 6656 26441 6684 26540
rect 6914 26528 6920 26540
rect 6972 26528 6978 26580
rect 11701 26571 11759 26577
rect 11701 26537 11713 26571
rect 11747 26568 11759 26571
rect 11790 26568 11796 26580
rect 11747 26540 11796 26568
rect 11747 26537 11759 26540
rect 11701 26531 11759 26537
rect 11790 26528 11796 26540
rect 11848 26528 11854 26580
rect 13541 26571 13599 26577
rect 13541 26537 13553 26571
rect 13587 26568 13599 26571
rect 16850 26568 16856 26580
rect 13587 26540 16856 26568
rect 13587 26537 13599 26540
rect 13541 26531 13599 26537
rect 16850 26528 16856 26540
rect 16908 26528 16914 26580
rect 17310 26568 17316 26580
rect 17271 26540 17316 26568
rect 17310 26528 17316 26540
rect 17368 26528 17374 26580
rect 23106 26568 23112 26580
rect 23067 26540 23112 26568
rect 23106 26528 23112 26540
rect 23164 26528 23170 26580
rect 25774 26568 25780 26580
rect 25735 26540 25780 26568
rect 25774 26528 25780 26540
rect 25832 26528 25838 26580
rect 28994 26568 29000 26580
rect 28955 26540 29000 26568
rect 28994 26528 29000 26540
rect 29052 26528 29058 26580
rect 41230 26568 41236 26580
rect 41191 26540 41236 26568
rect 41230 26528 41236 26540
rect 41288 26528 41294 26580
rect 42518 26528 42524 26580
rect 42576 26568 42582 26580
rect 43349 26571 43407 26577
rect 43349 26568 43361 26571
rect 42576 26540 43361 26568
rect 42576 26528 42582 26540
rect 43349 26537 43361 26540
rect 43395 26537 43407 26571
rect 46382 26568 46388 26580
rect 46343 26540 46388 26568
rect 43349 26531 43407 26537
rect 46382 26528 46388 26540
rect 46440 26528 46446 26580
rect 48130 26528 48136 26580
rect 48188 26568 48194 26580
rect 48225 26571 48283 26577
rect 48225 26568 48237 26571
rect 48188 26540 48237 26568
rect 48188 26528 48194 26540
rect 48225 26537 48237 26540
rect 48271 26537 48283 26571
rect 48225 26531 48283 26537
rect 51442 26528 51448 26580
rect 51500 26568 51506 26580
rect 51537 26571 51595 26577
rect 51537 26568 51549 26571
rect 51500 26540 51549 26568
rect 51500 26528 51506 26540
rect 51537 26537 51549 26540
rect 51583 26537 51595 26571
rect 54754 26568 54760 26580
rect 54715 26540 54760 26568
rect 51537 26531 51595 26537
rect 54754 26528 54760 26540
rect 54812 26528 54818 26580
rect 15470 26500 15476 26512
rect 15431 26472 15476 26500
rect 15470 26460 15476 26472
rect 15528 26460 15534 26512
rect 30929 26503 30987 26509
rect 30929 26469 30941 26503
rect 30975 26500 30987 26503
rect 31202 26500 31208 26512
rect 30975 26472 31208 26500
rect 30975 26469 30987 26472
rect 30929 26463 30987 26469
rect 31202 26460 31208 26472
rect 31260 26460 31266 26512
rect 57054 26460 57060 26512
rect 57112 26500 57118 26512
rect 57793 26503 57851 26509
rect 57793 26500 57805 26503
rect 57112 26472 57805 26500
rect 57112 26460 57118 26472
rect 57793 26469 57805 26472
rect 57839 26469 57851 26503
rect 57793 26463 57851 26469
rect 6641 26435 6699 26441
rect 6641 26401 6653 26435
rect 6687 26401 6699 26435
rect 6641 26395 6699 26401
rect 19242 26392 19248 26444
rect 19300 26432 19306 26444
rect 19889 26435 19947 26441
rect 19889 26432 19901 26435
rect 19300 26404 19901 26432
rect 19300 26392 19306 26404
rect 19889 26401 19901 26404
rect 19935 26401 19947 26435
rect 46842 26432 46848 26444
rect 46803 26404 46848 26432
rect 19889 26395 19947 26401
rect 46842 26392 46848 26404
rect 46900 26392 46906 26444
rect 50154 26432 50160 26444
rect 50115 26404 50160 26432
rect 50154 26392 50160 26404
rect 50212 26392 50218 26444
rect 6908 26367 6966 26373
rect 6908 26333 6920 26367
rect 6954 26364 6966 26367
rect 9122 26364 9128 26376
rect 6954 26336 9128 26364
rect 6954 26333 6966 26336
rect 6908 26327 6966 26333
rect 9122 26324 9128 26336
rect 9180 26324 9186 26376
rect 10318 26364 10324 26376
rect 10279 26336 10324 26364
rect 10318 26324 10324 26336
rect 10376 26324 10382 26376
rect 12066 26324 12072 26376
rect 12124 26364 12130 26376
rect 12161 26367 12219 26373
rect 12161 26364 12173 26367
rect 12124 26336 12173 26364
rect 12124 26324 12130 26336
rect 12161 26333 12173 26336
rect 12207 26364 12219 26367
rect 12250 26364 12256 26376
rect 12207 26336 12256 26364
rect 12207 26333 12219 26336
rect 12161 26327 12219 26333
rect 12250 26324 12256 26336
rect 12308 26324 12314 26376
rect 13630 26364 13636 26376
rect 12360 26336 13636 26364
rect 10588 26299 10646 26305
rect 10588 26265 10600 26299
rect 10634 26296 10646 26299
rect 12360 26296 12388 26336
rect 13630 26324 13636 26336
rect 13688 26324 13694 26376
rect 14090 26364 14096 26376
rect 14003 26336 14096 26364
rect 14090 26324 14096 26336
rect 14148 26364 14154 26376
rect 15102 26364 15108 26376
rect 14148 26336 15108 26364
rect 14148 26324 14154 26336
rect 15102 26324 15108 26336
rect 15160 26364 15166 26376
rect 15930 26364 15936 26376
rect 15160 26336 15936 26364
rect 15160 26324 15166 26336
rect 15930 26324 15936 26336
rect 15988 26324 15994 26376
rect 20156 26367 20214 26373
rect 20156 26333 20168 26367
rect 20202 26364 20214 26367
rect 21266 26364 21272 26376
rect 20202 26336 21272 26364
rect 20202 26333 20214 26336
rect 20156 26327 20214 26333
rect 21266 26324 21272 26336
rect 21324 26324 21330 26376
rect 21729 26367 21787 26373
rect 21729 26333 21741 26367
rect 21775 26333 21787 26367
rect 21729 26327 21787 26333
rect 21996 26367 22054 26373
rect 21996 26333 22008 26367
rect 22042 26364 22054 26367
rect 23198 26364 23204 26376
rect 22042 26336 23204 26364
rect 22042 26333 22054 26336
rect 21996 26327 22054 26333
rect 10634 26268 12388 26296
rect 12428 26299 12486 26305
rect 10634 26265 10646 26268
rect 10588 26259 10646 26265
rect 12428 26265 12440 26299
rect 12474 26296 12486 26299
rect 14182 26296 14188 26308
rect 12474 26268 14188 26296
rect 12474 26265 12486 26268
rect 12428 26259 12486 26265
rect 14182 26256 14188 26268
rect 14240 26256 14246 26308
rect 14360 26299 14418 26305
rect 14360 26265 14372 26299
rect 14406 26296 14418 26299
rect 16022 26296 16028 26308
rect 14406 26268 16028 26296
rect 14406 26265 14418 26268
rect 14360 26259 14418 26265
rect 16022 26256 16028 26268
rect 16080 26256 16086 26308
rect 16200 26299 16258 26305
rect 16200 26265 16212 26299
rect 16246 26296 16258 26299
rect 17862 26296 17868 26308
rect 16246 26268 17868 26296
rect 16246 26265 16258 26268
rect 16200 26259 16258 26265
rect 17862 26256 17868 26268
rect 17920 26256 17926 26308
rect 19978 26256 19984 26308
rect 20036 26296 20042 26308
rect 21744 26296 21772 26327
rect 23198 26324 23204 26336
rect 23256 26324 23262 26376
rect 24397 26367 24455 26373
rect 24397 26333 24409 26367
rect 24443 26364 24455 26367
rect 25130 26364 25136 26376
rect 24443 26336 25136 26364
rect 24443 26333 24455 26336
rect 24397 26327 24455 26333
rect 25130 26324 25136 26336
rect 25188 26324 25194 26376
rect 27614 26364 27620 26376
rect 27527 26336 27620 26364
rect 27614 26324 27620 26336
rect 27672 26324 27678 26376
rect 27890 26373 27896 26376
rect 27884 26364 27896 26373
rect 27851 26336 27896 26364
rect 27884 26327 27896 26336
rect 27890 26324 27896 26327
rect 27948 26324 27954 26376
rect 28902 26324 28908 26376
rect 28960 26364 28966 26376
rect 29546 26364 29552 26376
rect 28960 26336 29552 26364
rect 28960 26324 28966 26336
rect 29546 26324 29552 26336
rect 29604 26364 29610 26376
rect 30190 26364 30196 26376
rect 29604 26336 30196 26364
rect 29604 26324 29610 26336
rect 30190 26324 30196 26336
rect 30248 26364 30254 26376
rect 31389 26367 31447 26373
rect 31389 26364 31401 26367
rect 30248 26336 31401 26364
rect 30248 26324 30254 26336
rect 31389 26333 31401 26336
rect 31435 26333 31447 26367
rect 31389 26327 31447 26333
rect 31656 26367 31714 26373
rect 31656 26333 31668 26367
rect 31702 26364 31714 26367
rect 32766 26364 32772 26376
rect 31702 26336 32772 26364
rect 31702 26333 31714 26336
rect 31656 26327 31714 26333
rect 32766 26324 32772 26336
rect 32824 26324 32830 26376
rect 33962 26324 33968 26376
rect 34020 26364 34026 26376
rect 34701 26367 34759 26373
rect 34701 26364 34713 26367
rect 34020 26336 34713 26364
rect 34020 26324 34026 26336
rect 34701 26333 34713 26336
rect 34747 26333 34759 26367
rect 34701 26327 34759 26333
rect 36541 26367 36599 26373
rect 36541 26333 36553 26367
rect 36587 26364 36599 26367
rect 37274 26364 37280 26376
rect 36587 26336 37280 26364
rect 36587 26333 36599 26336
rect 36541 26327 36599 26333
rect 37274 26324 37280 26336
rect 37332 26324 37338 26376
rect 39850 26364 39856 26376
rect 39811 26336 39856 26364
rect 39850 26324 39856 26336
rect 39908 26324 39914 26376
rect 42058 26364 42064 26376
rect 42019 26336 42064 26364
rect 42058 26324 42064 26336
rect 42116 26324 42122 26376
rect 45002 26364 45008 26376
rect 44963 26336 45008 26364
rect 45002 26324 45008 26336
rect 45060 26324 45066 26376
rect 50424 26367 50482 26373
rect 50424 26333 50436 26367
rect 50470 26364 50482 26367
rect 51534 26364 51540 26376
rect 50470 26336 51540 26364
rect 50470 26333 50482 26336
rect 50424 26327 50482 26333
rect 51534 26324 51540 26336
rect 51592 26324 51598 26376
rect 53377 26367 53435 26373
rect 53377 26333 53389 26367
rect 53423 26364 53435 26367
rect 54110 26364 54116 26376
rect 53423 26336 54116 26364
rect 53423 26333 53435 26336
rect 53377 26327 53435 26333
rect 54110 26324 54116 26336
rect 54168 26324 54174 26376
rect 56502 26364 56508 26376
rect 56463 26336 56508 26364
rect 56502 26324 56508 26336
rect 56560 26324 56566 26376
rect 22462 26296 22468 26308
rect 20036 26268 22468 26296
rect 20036 26256 20042 26268
rect 22462 26256 22468 26268
rect 22520 26296 22526 26308
rect 23382 26296 23388 26308
rect 22520 26268 23388 26296
rect 22520 26256 22526 26268
rect 23382 26256 23388 26268
rect 23440 26256 23446 26308
rect 24664 26299 24722 26305
rect 24664 26265 24676 26299
rect 24710 26296 24722 26299
rect 25498 26296 25504 26308
rect 24710 26268 25504 26296
rect 24710 26265 24722 26268
rect 24664 26259 24722 26265
rect 25498 26256 25504 26268
rect 25556 26256 25562 26308
rect 26970 26256 26976 26308
rect 27028 26296 27034 26308
rect 27632 26296 27660 26324
rect 28920 26296 28948 26324
rect 27028 26268 28948 26296
rect 29816 26299 29874 26305
rect 27028 26256 27034 26268
rect 29816 26265 29828 26299
rect 29862 26296 29874 26299
rect 31294 26296 31300 26308
rect 29862 26268 31300 26296
rect 29862 26265 29874 26268
rect 29816 26259 29874 26265
rect 31294 26256 31300 26268
rect 31352 26256 31358 26308
rect 34514 26256 34520 26308
rect 34572 26296 34578 26308
rect 34946 26299 35004 26305
rect 34946 26296 34958 26299
rect 34572 26268 34958 26296
rect 34572 26256 34578 26268
rect 34946 26265 34958 26268
rect 34992 26265 35004 26299
rect 34946 26259 35004 26265
rect 36170 26256 36176 26308
rect 36228 26296 36234 26308
rect 36786 26299 36844 26305
rect 36786 26296 36798 26299
rect 36228 26268 36798 26296
rect 36228 26256 36234 26268
rect 36786 26265 36798 26268
rect 36832 26265 36844 26299
rect 36786 26259 36844 26265
rect 40120 26299 40178 26305
rect 40120 26265 40132 26299
rect 40166 26296 40178 26299
rect 41138 26296 41144 26308
rect 40166 26268 41144 26296
rect 40166 26265 40178 26268
rect 40120 26259 40178 26265
rect 41138 26256 41144 26268
rect 41196 26256 41202 26308
rect 45272 26299 45330 26305
rect 45272 26265 45284 26299
rect 45318 26296 45330 26299
rect 45922 26296 45928 26308
rect 45318 26268 45928 26296
rect 45318 26265 45330 26268
rect 45272 26259 45330 26265
rect 45922 26256 45928 26268
rect 45980 26256 45986 26308
rect 47112 26299 47170 26305
rect 47112 26265 47124 26299
rect 47158 26296 47170 26299
rect 48130 26296 48136 26308
rect 47158 26268 48136 26296
rect 47158 26265 47170 26268
rect 47112 26259 47170 26265
rect 48130 26256 48136 26268
rect 48188 26256 48194 26308
rect 53644 26299 53702 26305
rect 53644 26265 53656 26299
rect 53690 26296 53702 26299
rect 54754 26296 54760 26308
rect 53690 26268 54760 26296
rect 53690 26265 53702 26268
rect 53644 26259 53702 26265
rect 54754 26256 54760 26268
rect 54812 26256 54818 26308
rect 8018 26228 8024 26240
rect 7979 26200 8024 26228
rect 8018 26188 8024 26200
rect 8076 26188 8082 26240
rect 21266 26228 21272 26240
rect 21227 26200 21272 26228
rect 21266 26188 21272 26200
rect 21324 26188 21330 26240
rect 32766 26228 32772 26240
rect 32727 26200 32772 26228
rect 32766 26188 32772 26200
rect 32824 26188 32830 26240
rect 36078 26228 36084 26240
rect 36039 26200 36084 26228
rect 36078 26188 36084 26200
rect 36136 26188 36142 26240
rect 37918 26228 37924 26240
rect 37879 26200 37924 26228
rect 37918 26188 37924 26200
rect 37976 26188 37982 26240
rect 1104 26138 59340 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 59340 26138
rect 1104 26064 59340 26086
rect 8478 26024 8484 26036
rect 8439 25996 8484 26024
rect 8478 25984 8484 25996
rect 8536 25984 8542 26036
rect 13541 26027 13599 26033
rect 13541 25993 13553 26027
rect 13587 25993 13599 26027
rect 13541 25987 13599 25993
rect 7368 25959 7426 25965
rect 7368 25925 7380 25959
rect 7414 25956 7426 25959
rect 8018 25956 8024 25968
rect 7414 25928 8024 25956
rect 7414 25925 7426 25928
rect 7368 25919 7426 25925
rect 8018 25916 8024 25928
rect 8076 25916 8082 25968
rect 9030 25916 9036 25968
rect 9088 25956 9094 25968
rect 9186 25959 9244 25965
rect 9186 25956 9198 25959
rect 9088 25928 9198 25956
rect 9088 25916 9094 25928
rect 9186 25925 9198 25928
rect 9232 25925 9244 25959
rect 13556 25956 13584 25987
rect 16850 25984 16856 26036
rect 16908 26024 16914 26036
rect 16908 25996 16988 26024
rect 16908 25984 16914 25996
rect 16960 25965 16988 25996
rect 17862 25984 17868 26036
rect 17920 26024 17926 26036
rect 18049 26027 18107 26033
rect 18049 26024 18061 26027
rect 17920 25996 18061 26024
rect 17920 25984 17926 25996
rect 18049 25993 18061 25996
rect 18095 25993 18107 26027
rect 25498 26024 25504 26036
rect 25459 25996 25504 26024
rect 18049 25987 18107 25993
rect 25498 25984 25504 25996
rect 25556 25984 25562 26036
rect 31294 25984 31300 26036
rect 31352 26024 31358 26036
rect 31389 26027 31447 26033
rect 31389 26024 31401 26027
rect 31352 25996 31401 26024
rect 31352 25984 31358 25996
rect 31389 25993 31401 25996
rect 31435 25993 31447 26027
rect 38654 26024 38660 26036
rect 38615 25996 38660 26024
rect 31389 25987 31447 25993
rect 38654 25984 38660 25996
rect 38712 25984 38718 26036
rect 39298 25984 39304 26036
rect 39356 26024 39362 26036
rect 39356 25996 39436 26024
rect 39356 25984 39362 25996
rect 14246 25959 14304 25965
rect 14246 25956 14258 25959
rect 13556 25928 14258 25956
rect 9186 25919 9244 25925
rect 14246 25925 14258 25928
rect 14292 25925 14304 25959
rect 14246 25919 14304 25925
rect 16936 25959 16994 25965
rect 16936 25925 16948 25959
rect 16982 25925 16994 25959
rect 16936 25919 16994 25925
rect 23474 25916 23480 25968
rect 23532 25956 23538 25968
rect 24946 25956 24952 25968
rect 23532 25928 24952 25956
rect 23532 25916 23538 25928
rect 4700 25891 4758 25897
rect 4700 25857 4712 25891
rect 4746 25888 4758 25891
rect 5166 25888 5172 25900
rect 4746 25860 5172 25888
rect 4746 25857 4758 25860
rect 4700 25851 4758 25857
rect 5166 25848 5172 25860
rect 5224 25848 5230 25900
rect 6914 25848 6920 25900
rect 6972 25888 6978 25900
rect 7101 25891 7159 25897
rect 7101 25888 7113 25891
rect 6972 25860 7113 25888
rect 6972 25848 6978 25860
rect 7101 25857 7113 25860
rect 7147 25857 7159 25891
rect 9582 25888 9588 25900
rect 7101 25851 7159 25857
rect 8956 25860 9588 25888
rect 8956 25832 8984 25860
rect 9582 25848 9588 25860
rect 9640 25888 9646 25900
rect 10318 25888 10324 25900
rect 9640 25860 10324 25888
rect 9640 25848 9646 25860
rect 10318 25848 10324 25860
rect 10376 25848 10382 25900
rect 12428 25891 12486 25897
rect 12428 25857 12440 25891
rect 12474 25888 12486 25891
rect 13538 25888 13544 25900
rect 12474 25860 13544 25888
rect 12474 25857 12486 25860
rect 12428 25851 12486 25857
rect 13538 25848 13544 25860
rect 13596 25848 13602 25900
rect 14090 25848 14096 25900
rect 14148 25848 14154 25900
rect 15470 25848 15476 25900
rect 15528 25888 15534 25900
rect 15930 25888 15936 25900
rect 15528 25860 15936 25888
rect 15528 25848 15534 25860
rect 15930 25848 15936 25860
rect 15988 25888 15994 25900
rect 16669 25891 16727 25897
rect 16669 25888 16681 25891
rect 15988 25860 16681 25888
rect 15988 25848 15994 25860
rect 16669 25857 16681 25860
rect 16715 25857 16727 25891
rect 16669 25851 16727 25857
rect 18601 25891 18659 25897
rect 18601 25857 18613 25891
rect 18647 25888 18659 25891
rect 20070 25888 20076 25900
rect 18647 25860 20076 25888
rect 18647 25857 18659 25860
rect 18601 25851 18659 25857
rect 20070 25848 20076 25860
rect 20128 25888 20134 25900
rect 20898 25888 20904 25900
rect 20128 25860 20904 25888
rect 20128 25848 20134 25860
rect 20898 25848 20904 25860
rect 20956 25848 20962 25900
rect 22088 25891 22146 25897
rect 22088 25857 22100 25891
rect 22134 25888 22146 25891
rect 23106 25888 23112 25900
rect 22134 25860 23112 25888
rect 22134 25857 22146 25860
rect 22088 25851 22146 25857
rect 23106 25848 23112 25860
rect 23164 25848 23170 25900
rect 24136 25897 24164 25928
rect 24946 25916 24952 25928
rect 25004 25916 25010 25968
rect 35428 25959 35486 25965
rect 35428 25925 35440 25959
rect 35474 25956 35486 25959
rect 36078 25956 36084 25968
rect 35474 25928 36084 25956
rect 35474 25925 35486 25928
rect 35428 25919 35486 25925
rect 36078 25916 36084 25928
rect 36136 25916 36142 25968
rect 39408 25965 39436 25996
rect 44450 25984 44456 26036
rect 44508 26024 44514 26036
rect 57330 26024 57336 26036
rect 44508 25996 44588 26024
rect 57291 25996 57336 26024
rect 44508 25984 44514 25996
rect 44560 25965 44588 25996
rect 57330 25984 57336 25996
rect 57388 25984 57394 26036
rect 39384 25959 39442 25965
rect 39384 25925 39396 25959
rect 39430 25925 39442 25959
rect 39384 25919 39442 25925
rect 44536 25959 44594 25965
rect 44536 25925 44548 25959
rect 44582 25925 44594 25959
rect 44536 25919 44594 25925
rect 50424 25959 50482 25965
rect 50424 25925 50436 25959
rect 50470 25956 50482 25959
rect 50614 25956 50620 25968
rect 50470 25928 50620 25956
rect 50470 25925 50482 25928
rect 50424 25919 50482 25925
rect 50614 25916 50620 25928
rect 50672 25916 50678 25968
rect 54380 25959 54438 25965
rect 54380 25925 54392 25959
rect 54426 25956 54438 25959
rect 56594 25956 56600 25968
rect 54426 25928 56600 25956
rect 54426 25925 54438 25928
rect 54380 25919 54438 25925
rect 56594 25916 56600 25928
rect 56652 25916 56658 25968
rect 24121 25891 24179 25897
rect 24121 25857 24133 25891
rect 24167 25857 24179 25891
rect 24121 25851 24179 25857
rect 24388 25891 24446 25897
rect 24388 25857 24400 25891
rect 24434 25888 24446 25891
rect 25498 25888 25504 25900
rect 24434 25860 25504 25888
rect 24434 25857 24446 25860
rect 24388 25851 24446 25857
rect 25498 25848 25504 25860
rect 25556 25848 25562 25900
rect 26970 25888 26976 25900
rect 26931 25860 26976 25888
rect 26970 25848 26976 25860
rect 27028 25848 27034 25900
rect 27240 25891 27298 25897
rect 27240 25857 27252 25891
rect 27286 25888 27298 25891
rect 27706 25888 27712 25900
rect 27286 25860 27712 25888
rect 27286 25857 27298 25860
rect 27240 25851 27298 25857
rect 27706 25848 27712 25860
rect 27764 25848 27770 25900
rect 30009 25891 30067 25897
rect 30009 25857 30021 25891
rect 30055 25888 30067 25891
rect 30098 25888 30104 25900
rect 30055 25860 30104 25888
rect 30055 25857 30067 25860
rect 30009 25851 30067 25857
rect 30098 25848 30104 25860
rect 30156 25848 30162 25900
rect 30276 25891 30334 25897
rect 30276 25857 30288 25891
rect 30322 25888 30334 25891
rect 30834 25888 30840 25900
rect 30322 25860 30840 25888
rect 30322 25857 30334 25860
rect 30276 25851 30334 25857
rect 30834 25848 30840 25860
rect 30892 25848 30898 25900
rect 32950 25888 32956 25900
rect 32911 25860 32956 25888
rect 32950 25848 32956 25860
rect 33008 25848 33014 25900
rect 37544 25891 37602 25897
rect 37544 25857 37556 25891
rect 37590 25888 37602 25891
rect 38654 25888 38660 25900
rect 37590 25860 38660 25888
rect 37590 25857 37602 25860
rect 37544 25851 37602 25857
rect 38654 25848 38660 25860
rect 38712 25848 38718 25900
rect 39117 25891 39175 25897
rect 39117 25857 39129 25891
rect 39163 25888 39175 25891
rect 39850 25888 39856 25900
rect 39163 25860 39856 25888
rect 39163 25857 39175 25860
rect 39117 25851 39175 25857
rect 39850 25848 39856 25860
rect 39908 25848 39914 25900
rect 42696 25891 42754 25897
rect 42696 25857 42708 25891
rect 42742 25888 42754 25891
rect 43070 25888 43076 25900
rect 42742 25860 43076 25888
rect 42742 25857 42754 25860
rect 42696 25851 42754 25857
rect 43070 25848 43076 25860
rect 43128 25848 43134 25900
rect 44269 25891 44327 25897
rect 44269 25857 44281 25891
rect 44315 25888 44327 25891
rect 44358 25888 44364 25900
rect 44315 25860 44364 25888
rect 44315 25857 44327 25860
rect 44269 25851 44327 25857
rect 44358 25848 44364 25860
rect 44416 25848 44422 25900
rect 47946 25888 47952 25900
rect 47859 25860 47952 25888
rect 47946 25848 47952 25860
rect 48004 25888 48010 25900
rect 49418 25888 49424 25900
rect 48004 25860 49424 25888
rect 48004 25848 48010 25860
rect 49418 25848 49424 25860
rect 49476 25848 49482 25900
rect 50154 25888 50160 25900
rect 50115 25860 50160 25888
rect 50154 25848 50160 25860
rect 50212 25848 50218 25900
rect 56220 25891 56278 25897
rect 56220 25857 56232 25891
rect 56266 25888 56278 25891
rect 58158 25888 58164 25900
rect 56266 25860 58164 25888
rect 56266 25857 56278 25860
rect 56220 25851 56278 25857
rect 58158 25848 58164 25860
rect 58216 25848 58222 25900
rect 4433 25823 4491 25829
rect 4433 25789 4445 25823
rect 4479 25789 4491 25823
rect 8938 25820 8944 25832
rect 8899 25792 8944 25820
rect 4433 25783 4491 25789
rect 4448 25684 4476 25783
rect 8938 25780 8944 25792
rect 8996 25780 9002 25832
rect 12066 25780 12072 25832
rect 12124 25820 12130 25832
rect 12161 25823 12219 25829
rect 12161 25820 12173 25823
rect 12124 25792 12173 25820
rect 12124 25780 12130 25792
rect 12161 25789 12173 25792
rect 12207 25789 12219 25823
rect 12161 25783 12219 25789
rect 14001 25823 14059 25829
rect 14001 25789 14013 25823
rect 14047 25820 14059 25823
rect 14108 25820 14136 25848
rect 14047 25792 14136 25820
rect 14047 25789 14059 25792
rect 14001 25783 14059 25789
rect 4614 25684 4620 25696
rect 4448 25656 4620 25684
rect 4614 25644 4620 25656
rect 4672 25644 4678 25696
rect 5810 25684 5816 25696
rect 5771 25656 5816 25684
rect 5810 25644 5816 25656
rect 5868 25644 5874 25696
rect 10318 25684 10324 25696
rect 10279 25656 10324 25684
rect 10318 25644 10324 25656
rect 10376 25644 10382 25696
rect 12176 25684 12204 25783
rect 14016 25684 14044 25783
rect 19886 25780 19892 25832
rect 19944 25820 19950 25832
rect 20349 25823 20407 25829
rect 20349 25820 20361 25823
rect 19944 25792 20361 25820
rect 19944 25780 19950 25792
rect 20349 25789 20361 25792
rect 20395 25820 20407 25823
rect 21818 25820 21824 25832
rect 20395 25792 21824 25820
rect 20395 25789 20407 25792
rect 20349 25783 20407 25789
rect 21818 25780 21824 25792
rect 21876 25780 21882 25832
rect 35161 25823 35219 25829
rect 35161 25820 35173 25823
rect 34256 25792 35173 25820
rect 15378 25684 15384 25696
rect 12176 25656 14044 25684
rect 15339 25656 15384 25684
rect 15378 25644 15384 25656
rect 15436 25644 15442 25696
rect 23201 25687 23259 25693
rect 23201 25653 23213 25687
rect 23247 25684 23259 25687
rect 24486 25684 24492 25696
rect 23247 25656 24492 25684
rect 23247 25653 23259 25656
rect 23201 25647 23259 25653
rect 24486 25644 24492 25656
rect 24544 25644 24550 25696
rect 28353 25687 28411 25693
rect 28353 25653 28365 25687
rect 28399 25684 28411 25687
rect 29086 25684 29092 25696
rect 28399 25656 29092 25684
rect 28399 25653 28411 25656
rect 28353 25647 28411 25653
rect 29086 25644 29092 25656
rect 29144 25644 29150 25696
rect 33962 25644 33968 25696
rect 34020 25684 34026 25696
rect 34256 25693 34284 25792
rect 35161 25789 35173 25792
rect 35207 25789 35219 25823
rect 37274 25820 37280 25832
rect 37235 25792 37280 25820
rect 35161 25783 35219 25789
rect 37274 25780 37280 25792
rect 37332 25780 37338 25832
rect 42426 25820 42432 25832
rect 42387 25792 42432 25820
rect 42426 25780 42432 25792
rect 42484 25780 42490 25832
rect 54110 25820 54116 25832
rect 54071 25792 54116 25820
rect 54110 25780 54116 25792
rect 54168 25780 54174 25832
rect 55953 25823 56011 25829
rect 55953 25789 55965 25823
rect 55999 25789 56011 25823
rect 55953 25783 56011 25789
rect 34241 25687 34299 25693
rect 34241 25684 34253 25687
rect 34020 25656 34253 25684
rect 34020 25644 34026 25656
rect 34241 25653 34253 25656
rect 34287 25653 34299 25687
rect 34241 25647 34299 25653
rect 35434 25644 35440 25696
rect 35492 25684 35498 25696
rect 36541 25687 36599 25693
rect 36541 25684 36553 25687
rect 35492 25656 36553 25684
rect 35492 25644 35498 25656
rect 36541 25653 36553 25656
rect 36587 25653 36599 25687
rect 40494 25684 40500 25696
rect 40455 25656 40500 25684
rect 36541 25647 36599 25653
rect 40494 25644 40500 25656
rect 40552 25644 40558 25696
rect 43806 25684 43812 25696
rect 43767 25656 43812 25684
rect 43806 25644 43812 25656
rect 43864 25644 43870 25696
rect 45646 25684 45652 25696
rect 45607 25656 45652 25684
rect 45646 25644 45652 25656
rect 45704 25644 45710 25696
rect 49421 25687 49479 25693
rect 49421 25653 49433 25687
rect 49467 25684 49479 25687
rect 49510 25684 49516 25696
rect 49467 25656 49516 25684
rect 49467 25653 49479 25656
rect 49421 25647 49479 25653
rect 49510 25644 49516 25656
rect 49568 25644 49574 25696
rect 51534 25684 51540 25696
rect 51495 25656 51540 25684
rect 51534 25644 51540 25656
rect 51592 25644 51598 25696
rect 55490 25684 55496 25696
rect 55451 25656 55496 25684
rect 55490 25644 55496 25656
rect 55548 25644 55554 25696
rect 55968 25684 55996 25783
rect 56870 25684 56876 25696
rect 55968 25656 56876 25684
rect 56870 25644 56876 25656
rect 56928 25644 56934 25696
rect 1104 25594 59340 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 59340 25594
rect 1104 25520 59340 25542
rect 13538 25480 13544 25492
rect 13499 25452 13544 25480
rect 13538 25440 13544 25452
rect 13596 25440 13602 25492
rect 14182 25440 14188 25492
rect 14240 25480 14246 25492
rect 16485 25483 16543 25489
rect 16485 25480 16497 25483
rect 14240 25452 16497 25480
rect 14240 25440 14246 25452
rect 16485 25449 16497 25452
rect 16531 25449 16543 25483
rect 23106 25480 23112 25492
rect 23067 25452 23112 25480
rect 16485 25443 16543 25449
rect 23106 25440 23112 25452
rect 23164 25440 23170 25492
rect 30834 25440 30840 25492
rect 30892 25480 30898 25492
rect 30929 25483 30987 25489
rect 30929 25480 30941 25483
rect 30892 25452 30941 25480
rect 30892 25440 30898 25452
rect 30929 25449 30941 25452
rect 30975 25449 30987 25483
rect 30929 25443 30987 25449
rect 32674 25440 32680 25492
rect 32732 25480 32738 25492
rect 32769 25483 32827 25489
rect 32769 25480 32781 25483
rect 32732 25452 32781 25480
rect 32732 25440 32738 25452
rect 32769 25449 32781 25452
rect 32815 25449 32827 25483
rect 43070 25480 43076 25492
rect 43031 25452 43076 25480
rect 32769 25443 32827 25449
rect 43070 25440 43076 25452
rect 43128 25440 43134 25492
rect 45922 25440 45928 25492
rect 45980 25480 45986 25492
rect 46385 25483 46443 25489
rect 46385 25480 46397 25483
rect 45980 25452 46397 25480
rect 45980 25440 45986 25452
rect 46385 25449 46397 25452
rect 46431 25449 46443 25483
rect 46385 25443 46443 25449
rect 48130 25440 48136 25492
rect 48188 25480 48194 25492
rect 48225 25483 48283 25489
rect 48225 25480 48237 25483
rect 48188 25452 48237 25480
rect 48188 25440 48194 25452
rect 48225 25449 48237 25452
rect 48271 25449 48283 25483
rect 54754 25480 54760 25492
rect 54715 25452 54760 25480
rect 48225 25443 48283 25449
rect 54754 25440 54760 25452
rect 54812 25440 54818 25492
rect 57054 25480 57060 25492
rect 56796 25452 57060 25480
rect 12161 25347 12219 25353
rect 12161 25344 12173 25347
rect 12084 25316 12173 25344
rect 4522 25276 4528 25288
rect 4483 25248 4528 25276
rect 4522 25236 4528 25248
rect 4580 25236 4586 25288
rect 6362 25276 6368 25288
rect 6323 25248 6368 25276
rect 6362 25236 6368 25248
rect 6420 25236 6426 25288
rect 8941 25279 8999 25285
rect 8941 25245 8953 25279
rect 8987 25245 8999 25279
rect 8941 25239 8999 25245
rect 9208 25279 9266 25285
rect 9208 25245 9220 25279
rect 9254 25276 9266 25279
rect 10318 25276 10324 25288
rect 9254 25248 10324 25276
rect 9254 25245 9266 25248
rect 9208 25239 9266 25245
rect 4792 25211 4850 25217
rect 4792 25177 4804 25211
rect 4838 25208 4850 25211
rect 4838 25180 6040 25208
rect 4838 25177 4850 25180
rect 4792 25171 4850 25177
rect 4338 25100 4344 25152
rect 4396 25140 4402 25152
rect 5905 25143 5963 25149
rect 5905 25140 5917 25143
rect 4396 25112 5917 25140
rect 4396 25100 4402 25112
rect 5905 25109 5917 25112
rect 5951 25109 5963 25143
rect 6012 25140 6040 25180
rect 6086 25168 6092 25220
rect 6144 25208 6150 25220
rect 6610 25211 6668 25217
rect 6610 25208 6622 25211
rect 6144 25180 6622 25208
rect 6144 25168 6150 25180
rect 6610 25177 6622 25180
rect 6656 25177 6668 25211
rect 8956 25208 8984 25239
rect 10318 25236 10324 25248
rect 10376 25236 10382 25288
rect 12084 25220 12112 25316
rect 12161 25313 12173 25316
rect 12207 25313 12219 25347
rect 12161 25307 12219 25313
rect 14734 25304 14740 25356
rect 14792 25344 14798 25356
rect 15105 25347 15163 25353
rect 15105 25344 15117 25347
rect 14792 25316 15117 25344
rect 14792 25304 14798 25316
rect 15105 25313 15117 25316
rect 15151 25313 15163 25347
rect 19886 25344 19892 25356
rect 19847 25316 19892 25344
rect 15105 25307 15163 25313
rect 12066 25208 12072 25220
rect 8956 25180 12072 25208
rect 6610 25171 6668 25177
rect 12066 25168 12072 25180
rect 12124 25168 12130 25220
rect 12428 25211 12486 25217
rect 12428 25177 12440 25211
rect 12474 25208 12486 25211
rect 13446 25208 13452 25220
rect 12474 25180 13452 25208
rect 12474 25177 12486 25180
rect 12428 25171 12486 25177
rect 13446 25168 13452 25180
rect 13504 25168 13510 25220
rect 15120 25208 15148 25307
rect 19886 25304 19892 25316
rect 19944 25304 19950 25356
rect 29546 25344 29552 25356
rect 29507 25316 29552 25344
rect 29546 25304 29552 25316
rect 29604 25304 29610 25356
rect 35710 25304 35716 25356
rect 35768 25344 35774 25356
rect 36541 25347 36599 25353
rect 36541 25344 36553 25347
rect 35768 25316 36553 25344
rect 35768 25304 35774 25316
rect 36541 25313 36553 25316
rect 36587 25313 36599 25347
rect 45002 25344 45008 25356
rect 44963 25316 45008 25344
rect 36541 25307 36599 25313
rect 45002 25304 45008 25316
rect 45060 25304 45066 25356
rect 56594 25304 56600 25356
rect 56652 25344 56658 25356
rect 56796 25353 56824 25452
rect 57054 25440 57060 25452
rect 57112 25440 57118 25492
rect 58158 25480 58164 25492
rect 58119 25452 58164 25480
rect 58158 25440 58164 25452
rect 58216 25440 58222 25492
rect 56781 25347 56839 25353
rect 56781 25344 56793 25347
rect 56652 25316 56793 25344
rect 56652 25304 56658 25316
rect 56781 25313 56793 25316
rect 56827 25313 56839 25347
rect 56781 25307 56839 25313
rect 15378 25285 15384 25288
rect 15372 25276 15384 25285
rect 15339 25248 15384 25276
rect 15372 25239 15384 25248
rect 15378 25236 15384 25239
rect 15436 25236 15442 25288
rect 16666 25276 16672 25288
rect 16546 25248 16672 25276
rect 16546 25208 16574 25248
rect 16666 25236 16672 25248
rect 16724 25276 16730 25288
rect 17310 25276 17316 25288
rect 16724 25248 17316 25276
rect 16724 25236 16730 25248
rect 17310 25236 17316 25248
rect 17368 25236 17374 25288
rect 20156 25279 20214 25285
rect 20156 25245 20168 25279
rect 20202 25276 20214 25279
rect 21266 25276 21272 25288
rect 20202 25248 21272 25276
rect 20202 25245 20214 25248
rect 20156 25239 20214 25245
rect 21266 25236 21272 25248
rect 21324 25236 21330 25288
rect 21726 25276 21732 25288
rect 21687 25248 21732 25276
rect 21726 25236 21732 25248
rect 21784 25236 21790 25288
rect 24397 25279 24455 25285
rect 24397 25245 24409 25279
rect 24443 25276 24455 25279
rect 24946 25276 24952 25288
rect 24443 25248 24952 25276
rect 24443 25245 24455 25248
rect 24397 25239 24455 25245
rect 24946 25236 24952 25248
rect 25004 25276 25010 25288
rect 26237 25279 26295 25285
rect 26237 25276 26249 25279
rect 25004 25248 26249 25276
rect 25004 25236 25010 25248
rect 26237 25245 26249 25248
rect 26283 25245 26295 25279
rect 26237 25239 26295 25245
rect 30098 25236 30104 25288
rect 30156 25276 30162 25288
rect 31386 25276 31392 25288
rect 30156 25248 31392 25276
rect 30156 25236 30162 25248
rect 31386 25236 31392 25248
rect 31444 25236 31450 25288
rect 31656 25279 31714 25285
rect 31656 25245 31668 25279
rect 31702 25276 31714 25279
rect 32766 25276 32772 25288
rect 31702 25248 32772 25276
rect 31702 25245 31714 25248
rect 31656 25239 31714 25245
rect 32766 25236 32772 25248
rect 32824 25236 32830 25288
rect 34701 25279 34759 25285
rect 34701 25245 34713 25279
rect 34747 25276 34759 25279
rect 36808 25279 36866 25285
rect 34747 25248 35894 25276
rect 34747 25245 34759 25248
rect 34701 25239 34759 25245
rect 15120 25180 16574 25208
rect 17580 25211 17638 25217
rect 17580 25177 17592 25211
rect 17626 25208 17638 25211
rect 19242 25208 19248 25220
rect 17626 25180 19248 25208
rect 17626 25177 17638 25180
rect 17580 25171 17638 25177
rect 19242 25168 19248 25180
rect 19300 25168 19306 25220
rect 21996 25211 22054 25217
rect 21996 25177 22008 25211
rect 22042 25208 22054 25211
rect 23198 25208 23204 25220
rect 22042 25180 23204 25208
rect 22042 25177 22054 25180
rect 21996 25171 22054 25177
rect 23198 25168 23204 25180
rect 23256 25168 23262 25220
rect 24664 25211 24722 25217
rect 24664 25177 24676 25211
rect 24710 25208 24722 25211
rect 25314 25208 25320 25220
rect 24710 25180 25320 25208
rect 24710 25177 24722 25180
rect 24664 25171 24722 25177
rect 25314 25168 25320 25180
rect 25372 25168 25378 25220
rect 26482 25211 26540 25217
rect 26482 25208 26494 25211
rect 26206 25180 26494 25208
rect 7745 25143 7803 25149
rect 7745 25140 7757 25143
rect 6012 25112 7757 25140
rect 5905 25103 5963 25109
rect 7745 25109 7757 25112
rect 7791 25109 7803 25143
rect 10318 25140 10324 25152
rect 10279 25112 10324 25140
rect 7745 25103 7803 25109
rect 10318 25100 10324 25112
rect 10376 25100 10382 25152
rect 18690 25140 18696 25152
rect 18651 25112 18696 25140
rect 18690 25100 18696 25112
rect 18748 25100 18754 25152
rect 21266 25140 21272 25152
rect 21227 25112 21272 25140
rect 21266 25100 21272 25112
rect 21324 25100 21330 25152
rect 25777 25143 25835 25149
rect 25777 25109 25789 25143
rect 25823 25140 25835 25143
rect 26206 25140 26234 25180
rect 26482 25177 26494 25180
rect 26528 25177 26540 25211
rect 26482 25171 26540 25177
rect 29816 25211 29874 25217
rect 29816 25177 29828 25211
rect 29862 25208 29874 25211
rect 30190 25208 30196 25220
rect 29862 25180 30196 25208
rect 29862 25177 29874 25180
rect 29816 25171 29874 25177
rect 30190 25168 30196 25180
rect 30248 25168 30254 25220
rect 34968 25211 35026 25217
rect 34968 25177 34980 25211
rect 35014 25208 35026 25211
rect 35434 25208 35440 25220
rect 35014 25180 35440 25208
rect 35014 25177 35026 25180
rect 34968 25171 35026 25177
rect 35434 25168 35440 25180
rect 35492 25168 35498 25220
rect 35866 25208 35894 25248
rect 36808 25245 36820 25279
rect 36854 25276 36866 25279
rect 37918 25276 37924 25288
rect 36854 25248 37924 25276
rect 36854 25245 36866 25248
rect 36808 25239 36866 25245
rect 37918 25236 37924 25248
rect 37976 25236 37982 25288
rect 39850 25276 39856 25288
rect 39811 25248 39856 25276
rect 39850 25236 39856 25248
rect 39908 25236 39914 25288
rect 40120 25279 40178 25285
rect 40120 25245 40132 25279
rect 40166 25276 40178 25279
rect 40494 25276 40500 25288
rect 40166 25248 40500 25276
rect 40166 25245 40178 25248
rect 40120 25239 40178 25245
rect 40494 25236 40500 25248
rect 40552 25236 40558 25288
rect 41693 25279 41751 25285
rect 41693 25245 41705 25279
rect 41739 25245 41751 25279
rect 41693 25239 41751 25245
rect 37274 25208 37280 25220
rect 35866 25180 37280 25208
rect 37274 25168 37280 25180
rect 37332 25168 37338 25220
rect 41708 25208 41736 25239
rect 41782 25236 41788 25288
rect 41840 25276 41846 25288
rect 41949 25279 42007 25285
rect 41949 25276 41961 25279
rect 41840 25248 41961 25276
rect 41840 25236 41846 25248
rect 41949 25245 41961 25248
rect 41995 25245 42007 25279
rect 41949 25239 42007 25245
rect 45272 25279 45330 25285
rect 45272 25245 45284 25279
rect 45318 25276 45330 25279
rect 45646 25276 45652 25288
rect 45318 25248 45652 25276
rect 45318 25245 45330 25248
rect 45272 25239 45330 25245
rect 45646 25236 45652 25248
rect 45704 25236 45710 25288
rect 46842 25276 46848 25288
rect 46803 25248 46848 25276
rect 46842 25236 46848 25248
rect 46900 25236 46906 25288
rect 46934 25236 46940 25288
rect 46992 25276 46998 25288
rect 47101 25279 47159 25285
rect 47101 25276 47113 25279
rect 46992 25248 47113 25276
rect 46992 25236 46998 25248
rect 47101 25245 47113 25248
rect 47147 25245 47159 25279
rect 47101 25239 47159 25245
rect 49510 25236 49516 25288
rect 49568 25276 49574 25288
rect 50157 25279 50215 25285
rect 50157 25276 50169 25279
rect 49568 25248 50169 25276
rect 49568 25236 49574 25248
rect 50157 25245 50169 25248
rect 50203 25245 50215 25279
rect 50157 25239 50215 25245
rect 50424 25279 50482 25285
rect 50424 25245 50436 25279
rect 50470 25276 50482 25279
rect 51534 25276 51540 25288
rect 50470 25248 51540 25276
rect 50470 25245 50482 25248
rect 50424 25239 50482 25245
rect 51534 25236 51540 25248
rect 51592 25236 51598 25288
rect 53377 25279 53435 25285
rect 53377 25245 53389 25279
rect 53423 25276 53435 25279
rect 54110 25276 54116 25288
rect 53423 25248 54116 25276
rect 53423 25245 53435 25248
rect 53377 25239 53435 25245
rect 54110 25236 54116 25248
rect 54168 25236 54174 25288
rect 42426 25208 42432 25220
rect 41708 25180 42432 25208
rect 42426 25168 42432 25180
rect 42484 25168 42490 25220
rect 44358 25168 44364 25220
rect 44416 25208 44422 25220
rect 44910 25208 44916 25220
rect 44416 25180 44916 25208
rect 44416 25168 44422 25180
rect 44910 25168 44916 25180
rect 44968 25208 44974 25220
rect 46860 25208 46888 25236
rect 44968 25180 46888 25208
rect 53644 25211 53702 25217
rect 44968 25168 44974 25180
rect 53644 25177 53656 25211
rect 53690 25208 53702 25211
rect 54754 25208 54760 25220
rect 53690 25180 54760 25208
rect 53690 25177 53702 25180
rect 53644 25171 53702 25177
rect 54754 25168 54760 25180
rect 54812 25168 54818 25220
rect 57048 25211 57106 25217
rect 57048 25177 57060 25211
rect 57094 25208 57106 25211
rect 57330 25208 57336 25220
rect 57094 25180 57336 25208
rect 57094 25177 57106 25180
rect 57048 25171 57106 25177
rect 57330 25168 57336 25180
rect 57388 25168 57394 25220
rect 27614 25140 27620 25152
rect 25823 25112 26234 25140
rect 27575 25112 27620 25140
rect 25823 25109 25835 25112
rect 25777 25103 25835 25109
rect 27614 25100 27620 25112
rect 27672 25100 27678 25152
rect 36078 25140 36084 25152
rect 36039 25112 36084 25140
rect 36078 25100 36084 25112
rect 36136 25100 36142 25152
rect 37918 25140 37924 25152
rect 37879 25112 37924 25140
rect 37918 25100 37924 25112
rect 37976 25100 37982 25152
rect 41230 25140 41236 25152
rect 41191 25112 41236 25140
rect 41230 25100 41236 25112
rect 41288 25100 41294 25152
rect 51534 25140 51540 25152
rect 51495 25112 51540 25140
rect 51534 25100 51540 25112
rect 51592 25100 51598 25152
rect 1104 25050 59340 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 59340 25050
rect 1104 24976 59340 24998
rect 5166 24936 5172 24948
rect 5127 24908 5172 24936
rect 5166 24896 5172 24908
rect 5224 24896 5230 24948
rect 13446 24896 13452 24948
rect 13504 24936 13510 24948
rect 13541 24939 13599 24945
rect 13541 24936 13553 24939
rect 13504 24908 13553 24936
rect 13504 24896 13510 24908
rect 13541 24905 13553 24908
rect 13587 24905 13599 24939
rect 23198 24936 23204 24948
rect 23159 24908 23204 24936
rect 13541 24899 13599 24905
rect 23198 24896 23204 24908
rect 23256 24896 23262 24948
rect 25498 24936 25504 24948
rect 25459 24908 25504 24936
rect 25498 24896 25504 24908
rect 25556 24896 25562 24948
rect 30190 24936 30196 24948
rect 30151 24908 30196 24936
rect 30190 24896 30196 24908
rect 30248 24896 30254 24948
rect 38654 24936 38660 24948
rect 38615 24908 38660 24936
rect 38654 24896 38660 24908
rect 38712 24896 38718 24948
rect 57330 24936 57336 24948
rect 57291 24908 57336 24936
rect 57330 24896 57336 24908
rect 57388 24896 57394 24948
rect 4522 24868 4528 24880
rect 2148 24840 3648 24868
rect 2148 24800 2176 24840
rect 1964 24772 2176 24800
rect 2216 24803 2274 24809
rect 1854 24692 1860 24744
rect 1912 24732 1918 24744
rect 1964 24741 1992 24772
rect 2216 24769 2228 24803
rect 2262 24800 2274 24803
rect 3620 24800 3648 24840
rect 3988 24840 4528 24868
rect 3789 24803 3847 24809
rect 3789 24800 3801 24803
rect 2262 24772 3556 24800
rect 3620 24772 3801 24800
rect 2262 24769 2274 24772
rect 2216 24763 2274 24769
rect 1949 24735 2007 24741
rect 1949 24732 1961 24735
rect 1912 24704 1961 24732
rect 1912 24692 1918 24704
rect 1949 24701 1961 24704
rect 1995 24701 2007 24735
rect 1949 24695 2007 24701
rect 3326 24596 3332 24608
rect 3287 24568 3332 24596
rect 3326 24556 3332 24568
rect 3384 24556 3390 24608
rect 3528 24596 3556 24772
rect 3789 24769 3801 24772
rect 3835 24800 3847 24803
rect 3988 24800 4016 24840
rect 4522 24828 4528 24840
rect 4580 24828 4586 24880
rect 8938 24828 8944 24880
rect 8996 24868 9002 24880
rect 8996 24840 9076 24868
rect 8996 24828 9002 24840
rect 3835 24772 4016 24800
rect 4056 24803 4114 24809
rect 3835 24769 3847 24772
rect 3789 24763 3847 24769
rect 4056 24769 4068 24803
rect 4102 24800 4114 24803
rect 4338 24800 4344 24812
rect 4102 24772 4344 24800
rect 4102 24769 4114 24772
rect 4056 24763 4114 24769
rect 4338 24760 4344 24772
rect 4396 24760 4402 24812
rect 4540 24800 4568 24828
rect 6362 24800 6368 24812
rect 4540 24772 6368 24800
rect 6362 24760 6368 24772
rect 6420 24760 6426 24812
rect 6632 24803 6690 24809
rect 6632 24769 6644 24803
rect 6678 24800 6690 24803
rect 8018 24800 8024 24812
rect 6678 24772 8024 24800
rect 6678 24769 6690 24772
rect 6632 24763 6690 24769
rect 8018 24760 8024 24772
rect 8076 24760 8082 24812
rect 9048 24809 9076 24840
rect 19978 24828 19984 24880
rect 20036 24828 20042 24880
rect 37544 24871 37602 24877
rect 37544 24837 37556 24871
rect 37590 24868 37602 24871
rect 37918 24868 37924 24880
rect 37590 24840 37924 24868
rect 37590 24837 37602 24840
rect 37544 24831 37602 24837
rect 37918 24828 37924 24840
rect 37976 24828 37982 24880
rect 56870 24868 56876 24880
rect 47780 24840 49464 24868
rect 9033 24803 9091 24809
rect 9033 24769 9045 24803
rect 9079 24769 9091 24803
rect 9033 24763 9091 24769
rect 9300 24803 9358 24809
rect 9300 24769 9312 24803
rect 9346 24800 9358 24803
rect 10318 24800 10324 24812
rect 9346 24772 10324 24800
rect 9346 24769 9358 24772
rect 9300 24763 9358 24769
rect 10318 24760 10324 24772
rect 10376 24760 10382 24812
rect 12066 24760 12072 24812
rect 12124 24800 12130 24812
rect 12161 24803 12219 24809
rect 12161 24800 12173 24803
rect 12124 24772 12173 24800
rect 12124 24760 12130 24772
rect 12161 24769 12173 24772
rect 12207 24769 12219 24803
rect 12161 24763 12219 24769
rect 12428 24803 12486 24809
rect 12428 24769 12440 24803
rect 12474 24800 12486 24803
rect 13446 24800 13452 24812
rect 12474 24772 13452 24800
rect 12474 24769 12486 24772
rect 12428 24763 12486 24769
rect 13446 24760 13452 24772
rect 13504 24760 13510 24812
rect 14734 24800 14740 24812
rect 14695 24772 14740 24800
rect 14734 24760 14740 24772
rect 14792 24760 14798 24812
rect 15004 24803 15062 24809
rect 15004 24769 15016 24803
rect 15050 24800 15062 24803
rect 17580 24803 17638 24809
rect 15050 24772 16574 24800
rect 15050 24769 15062 24772
rect 15004 24763 15062 24769
rect 5810 24596 5816 24608
rect 3528 24568 5816 24596
rect 5810 24556 5816 24568
rect 5868 24556 5874 24608
rect 6178 24556 6184 24608
rect 6236 24596 6242 24608
rect 7745 24599 7803 24605
rect 7745 24596 7757 24599
rect 6236 24568 7757 24596
rect 6236 24556 6242 24568
rect 7745 24565 7757 24568
rect 7791 24565 7803 24599
rect 10410 24596 10416 24608
rect 10371 24568 10416 24596
rect 7745 24559 7803 24565
rect 10410 24556 10416 24568
rect 10468 24556 10474 24608
rect 16114 24596 16120 24608
rect 16075 24568 16120 24596
rect 16114 24556 16120 24568
rect 16172 24556 16178 24608
rect 16546 24596 16574 24772
rect 17580 24769 17592 24803
rect 17626 24800 17638 24803
rect 18690 24800 18696 24812
rect 17626 24772 18696 24800
rect 17626 24769 17638 24772
rect 17580 24763 17638 24769
rect 18690 24760 18696 24772
rect 18748 24760 18754 24812
rect 19797 24803 19855 24809
rect 19797 24769 19809 24803
rect 19843 24800 19855 24803
rect 19996 24800 20024 24828
rect 19843 24772 20024 24800
rect 20064 24803 20122 24809
rect 19843 24769 19855 24772
rect 19797 24763 19855 24769
rect 20064 24769 20076 24803
rect 20110 24800 20122 24803
rect 21266 24800 21272 24812
rect 20110 24772 21272 24800
rect 20110 24769 20122 24772
rect 20064 24763 20122 24769
rect 21266 24760 21272 24772
rect 21324 24760 21330 24812
rect 21726 24760 21732 24812
rect 21784 24800 21790 24812
rect 21821 24803 21879 24809
rect 21821 24800 21833 24803
rect 21784 24772 21833 24800
rect 21784 24760 21790 24772
rect 21821 24769 21833 24772
rect 21867 24769 21879 24803
rect 21821 24763 21879 24769
rect 22088 24803 22146 24809
rect 22088 24769 22100 24803
rect 22134 24800 22146 24803
rect 23198 24800 23204 24812
rect 22134 24772 23204 24800
rect 22134 24769 22146 24772
rect 22088 24763 22146 24769
rect 23198 24760 23204 24772
rect 23256 24760 23262 24812
rect 24388 24803 24446 24809
rect 24388 24769 24400 24803
rect 24434 24800 24446 24803
rect 25498 24800 25504 24812
rect 24434 24772 25504 24800
rect 24434 24769 24446 24772
rect 24388 24763 24446 24769
rect 25498 24760 25504 24772
rect 25556 24760 25562 24812
rect 27240 24803 27298 24809
rect 27240 24769 27252 24803
rect 27286 24800 27298 24803
rect 28350 24800 28356 24812
rect 27286 24772 28356 24800
rect 27286 24769 27298 24772
rect 27240 24763 27298 24769
rect 28350 24760 28356 24772
rect 28408 24760 28414 24812
rect 28813 24803 28871 24809
rect 28813 24769 28825 24803
rect 28859 24800 28871 24803
rect 28902 24800 28908 24812
rect 28859 24772 28908 24800
rect 28859 24769 28871 24772
rect 28813 24763 28871 24769
rect 28902 24760 28908 24772
rect 28960 24760 28966 24812
rect 29080 24803 29138 24809
rect 29080 24769 29092 24803
rect 29126 24800 29138 24803
rect 30926 24800 30932 24812
rect 29126 24772 30932 24800
rect 29126 24769 29138 24772
rect 29080 24763 29138 24769
rect 30926 24760 30932 24772
rect 30984 24760 30990 24812
rect 31386 24760 31392 24812
rect 31444 24800 31450 24812
rect 32398 24809 32404 24812
rect 32125 24803 32183 24809
rect 32125 24800 32137 24803
rect 31444 24772 32137 24800
rect 31444 24760 31450 24772
rect 32125 24769 32137 24772
rect 32171 24769 32183 24803
rect 32392 24800 32404 24809
rect 32359 24772 32404 24800
rect 32125 24763 32183 24769
rect 32392 24763 32404 24772
rect 32398 24760 32404 24763
rect 32456 24760 32462 24812
rect 34221 24803 34279 24809
rect 34221 24800 34233 24803
rect 33520 24772 34233 24800
rect 17310 24732 17316 24744
rect 17271 24704 17316 24732
rect 17310 24692 17316 24704
rect 17368 24692 17374 24744
rect 24118 24732 24124 24744
rect 24079 24704 24124 24732
rect 24118 24692 24124 24704
rect 24176 24692 24182 24744
rect 26234 24692 26240 24744
rect 26292 24732 26298 24744
rect 26973 24735 27031 24741
rect 26973 24732 26985 24735
rect 26292 24704 26985 24732
rect 26292 24692 26298 24704
rect 26973 24701 26985 24704
rect 27019 24701 27031 24735
rect 26973 24695 27031 24701
rect 33520 24673 33548 24772
rect 34221 24769 34233 24772
rect 34267 24769 34279 24803
rect 37274 24800 37280 24812
rect 37187 24772 37280 24800
rect 34221 24763 34279 24769
rect 37274 24760 37280 24772
rect 37332 24800 37338 24812
rect 37826 24800 37832 24812
rect 37332 24772 37832 24800
rect 37332 24760 37338 24772
rect 37826 24760 37832 24772
rect 37884 24760 37890 24812
rect 38010 24760 38016 24812
rect 38068 24800 38074 24812
rect 39373 24803 39431 24809
rect 39373 24800 39385 24803
rect 38068 24772 39385 24800
rect 38068 24760 38074 24772
rect 39373 24769 39385 24772
rect 39419 24769 39431 24803
rect 39373 24763 39431 24769
rect 43070 24760 43076 24812
rect 43128 24800 43134 24812
rect 43421 24803 43479 24809
rect 43421 24800 43433 24803
rect 43128 24772 43433 24800
rect 43128 24760 43134 24772
rect 43421 24769 43433 24772
rect 43467 24769 43479 24803
rect 45261 24803 45319 24809
rect 45261 24800 45273 24803
rect 43421 24763 43479 24769
rect 44560 24772 45273 24800
rect 33962 24732 33968 24744
rect 33923 24704 33968 24732
rect 33962 24692 33968 24704
rect 34020 24692 34026 24744
rect 39117 24735 39175 24741
rect 39117 24701 39129 24735
rect 39163 24701 39175 24735
rect 39117 24695 39175 24701
rect 33505 24667 33563 24673
rect 33505 24633 33517 24667
rect 33551 24633 33563 24667
rect 33505 24627 33563 24633
rect 18506 24596 18512 24608
rect 16546 24568 18512 24596
rect 18506 24556 18512 24568
rect 18564 24556 18570 24608
rect 18690 24596 18696 24608
rect 18651 24568 18696 24596
rect 18690 24556 18696 24568
rect 18748 24556 18754 24608
rect 21174 24596 21180 24608
rect 21135 24568 21180 24596
rect 21174 24556 21180 24568
rect 21232 24556 21238 24608
rect 27890 24556 27896 24608
rect 27948 24596 27954 24608
rect 28353 24599 28411 24605
rect 28353 24596 28365 24599
rect 27948 24568 28365 24596
rect 27948 24556 27954 24568
rect 28353 24565 28365 24568
rect 28399 24565 28411 24599
rect 28353 24559 28411 24565
rect 32398 24556 32404 24608
rect 32456 24596 32462 24608
rect 35345 24599 35403 24605
rect 35345 24596 35357 24599
rect 32456 24568 35357 24596
rect 32456 24556 32462 24568
rect 35345 24565 35357 24568
rect 35391 24565 35403 24599
rect 39132 24596 39160 24695
rect 42426 24692 42432 24744
rect 42484 24732 42490 24744
rect 43165 24735 43223 24741
rect 43165 24732 43177 24735
rect 42484 24704 43177 24732
rect 42484 24692 42490 24704
rect 43165 24701 43177 24704
rect 43211 24701 43223 24735
rect 43165 24695 43223 24701
rect 40402 24624 40408 24676
rect 40460 24664 40466 24676
rect 40497 24667 40555 24673
rect 40497 24664 40509 24667
rect 40460 24636 40509 24664
rect 40460 24624 40466 24636
rect 40497 24633 40509 24636
rect 40543 24633 40555 24667
rect 40497 24627 40555 24633
rect 39850 24596 39856 24608
rect 39132 24568 39856 24596
rect 35345 24559 35403 24565
rect 39850 24556 39856 24568
rect 39908 24556 39914 24608
rect 43180 24596 43208 24695
rect 44560 24673 44588 24772
rect 45261 24769 45273 24772
rect 45307 24769 45319 24803
rect 45261 24763 45319 24769
rect 46842 24760 46848 24812
rect 46900 24800 46906 24812
rect 47581 24803 47639 24809
rect 47581 24800 47593 24803
rect 46900 24772 47593 24800
rect 46900 24760 46906 24772
rect 47581 24769 47593 24772
rect 47627 24800 47639 24803
rect 47780 24800 47808 24840
rect 47627 24772 47808 24800
rect 47848 24803 47906 24809
rect 47627 24769 47639 24772
rect 47581 24763 47639 24769
rect 47848 24769 47860 24803
rect 47894 24800 47906 24803
rect 48958 24800 48964 24812
rect 47894 24772 48964 24800
rect 47894 24769 47906 24772
rect 47848 24763 47906 24769
rect 48958 24760 48964 24772
rect 49016 24760 49022 24812
rect 49436 24809 49464 24840
rect 55968 24840 56876 24868
rect 49421 24803 49479 24809
rect 49421 24769 49433 24803
rect 49467 24800 49479 24803
rect 49510 24800 49516 24812
rect 49467 24772 49516 24800
rect 49467 24769 49479 24772
rect 49421 24763 49479 24769
rect 49510 24760 49516 24772
rect 49568 24760 49574 24812
rect 49688 24803 49746 24809
rect 49688 24769 49700 24803
rect 49734 24800 49746 24803
rect 51534 24800 51540 24812
rect 49734 24772 51540 24800
rect 49734 24769 49746 24772
rect 49688 24763 49746 24769
rect 51534 24760 51540 24772
rect 51592 24760 51598 24812
rect 54380 24803 54438 24809
rect 54380 24769 54392 24803
rect 54426 24800 54438 24803
rect 55490 24800 55496 24812
rect 54426 24772 55496 24800
rect 54426 24769 54438 24772
rect 54380 24763 54438 24769
rect 55490 24760 55496 24772
rect 55548 24760 55554 24812
rect 55968 24809 55996 24840
rect 56870 24828 56876 24840
rect 56928 24828 56934 24880
rect 55953 24803 56011 24809
rect 55953 24769 55965 24803
rect 55999 24769 56011 24803
rect 55953 24763 56011 24769
rect 56220 24803 56278 24809
rect 56220 24769 56232 24803
rect 56266 24800 56278 24803
rect 57330 24800 57336 24812
rect 56266 24772 57336 24800
rect 56266 24769 56278 24772
rect 56220 24763 56278 24769
rect 57330 24760 57336 24772
rect 57388 24760 57394 24812
rect 45002 24732 45008 24744
rect 44963 24704 45008 24732
rect 45002 24692 45008 24704
rect 45060 24692 45066 24744
rect 54110 24732 54116 24744
rect 54071 24704 54116 24732
rect 54110 24692 54116 24704
rect 54168 24692 54174 24744
rect 44545 24667 44603 24673
rect 44545 24633 44557 24667
rect 44591 24633 44603 24667
rect 44545 24627 44603 24633
rect 45020 24596 45048 24692
rect 46290 24624 46296 24676
rect 46348 24664 46354 24676
rect 46385 24667 46443 24673
rect 46385 24664 46397 24667
rect 46348 24636 46397 24664
rect 46348 24624 46354 24636
rect 46385 24633 46397 24636
rect 46431 24633 46443 24667
rect 46385 24627 46443 24633
rect 43180 24568 45048 24596
rect 45922 24556 45928 24608
rect 45980 24596 45986 24608
rect 48961 24599 49019 24605
rect 48961 24596 48973 24599
rect 45980 24568 48973 24596
rect 45980 24556 45986 24568
rect 48961 24565 48973 24568
rect 49007 24565 49019 24599
rect 48961 24559 49019 24565
rect 49694 24556 49700 24608
rect 49752 24596 49758 24608
rect 50801 24599 50859 24605
rect 50801 24596 50813 24599
rect 49752 24568 50813 24596
rect 49752 24556 49758 24568
rect 50801 24565 50813 24568
rect 50847 24565 50859 24599
rect 50801 24559 50859 24565
rect 55493 24599 55551 24605
rect 55493 24565 55505 24599
rect 55539 24596 55551 24599
rect 56686 24596 56692 24608
rect 55539 24568 56692 24596
rect 55539 24565 55551 24568
rect 55493 24559 55551 24565
rect 56686 24556 56692 24568
rect 56744 24556 56750 24608
rect 1104 24506 59340 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 59340 24506
rect 1104 24432 59340 24454
rect 6362 24352 6368 24404
rect 6420 24392 6426 24404
rect 6549 24395 6607 24401
rect 6549 24392 6561 24395
rect 6420 24364 6561 24392
rect 6420 24352 6426 24364
rect 6549 24361 6561 24364
rect 6595 24361 6607 24395
rect 6549 24355 6607 24361
rect 11514 24352 11520 24404
rect 11572 24392 11578 24404
rect 12434 24392 12440 24404
rect 11572 24364 12440 24392
rect 11572 24352 11578 24364
rect 12434 24352 12440 24364
rect 12492 24352 12498 24404
rect 13446 24392 13452 24404
rect 13407 24364 13452 24392
rect 13446 24352 13452 24364
rect 13504 24352 13510 24404
rect 25314 24352 25320 24404
rect 25372 24392 25378 24404
rect 25777 24395 25835 24401
rect 25777 24392 25789 24395
rect 25372 24364 25789 24392
rect 25372 24352 25378 24364
rect 25777 24361 25789 24364
rect 25823 24361 25835 24395
rect 30926 24392 30932 24404
rect 30887 24364 30932 24392
rect 25777 24355 25835 24361
rect 30926 24352 30932 24364
rect 30984 24352 30990 24404
rect 32582 24352 32588 24404
rect 32640 24392 32646 24404
rect 32769 24395 32827 24401
rect 32769 24392 32781 24395
rect 32640 24364 32781 24392
rect 32640 24352 32646 24364
rect 32769 24361 32781 24364
rect 32815 24361 32827 24395
rect 32769 24355 32827 24361
rect 37921 24395 37979 24401
rect 37921 24361 37933 24395
rect 37967 24392 37979 24395
rect 38010 24392 38016 24404
rect 37967 24364 38016 24392
rect 37967 24361 37979 24364
rect 37921 24355 37979 24361
rect 38010 24352 38016 24364
rect 38068 24352 38074 24404
rect 41138 24352 41144 24404
rect 41196 24392 41202 24404
rect 41233 24395 41291 24401
rect 41233 24392 41245 24395
rect 41196 24364 41245 24392
rect 41196 24352 41202 24364
rect 41233 24361 41245 24364
rect 41279 24361 41291 24395
rect 42426 24392 42432 24404
rect 41233 24355 41291 24361
rect 41708 24364 42432 24392
rect 1854 24256 1860 24268
rect 1815 24228 1860 24256
rect 1854 24216 1860 24228
rect 1912 24216 1918 24268
rect 15470 24256 15476 24268
rect 15431 24228 15476 24256
rect 15470 24216 15476 24228
rect 15528 24216 15534 24268
rect 31386 24256 31392 24268
rect 31347 24228 31392 24256
rect 31386 24216 31392 24228
rect 31444 24216 31450 24268
rect 33962 24216 33968 24268
rect 34020 24256 34026 24268
rect 34701 24259 34759 24265
rect 34701 24256 34713 24259
rect 34020 24228 34713 24256
rect 34020 24216 34026 24228
rect 34701 24225 34713 24228
rect 34747 24225 34759 24259
rect 34701 24219 34759 24225
rect 2124 24191 2182 24197
rect 2124 24157 2136 24191
rect 2170 24188 2182 24191
rect 3326 24188 3332 24200
rect 2170 24160 3332 24188
rect 2170 24157 2182 24160
rect 2124 24151 2182 24157
rect 3326 24148 3332 24160
rect 3384 24148 3390 24200
rect 9214 24148 9220 24200
rect 9272 24188 9278 24200
rect 9309 24191 9367 24197
rect 9309 24188 9321 24191
rect 9272 24160 9321 24188
rect 9272 24148 9278 24160
rect 9309 24157 9321 24160
rect 9355 24157 9367 24191
rect 9309 24151 9367 24157
rect 9576 24191 9634 24197
rect 9576 24157 9588 24191
rect 9622 24188 9634 24191
rect 10410 24188 10416 24200
rect 9622 24160 10416 24188
rect 9622 24157 9634 24160
rect 9576 24151 9634 24157
rect 10410 24148 10416 24160
rect 10468 24148 10474 24200
rect 11609 24191 11667 24197
rect 11609 24157 11621 24191
rect 11655 24157 11667 24191
rect 12066 24188 12072 24200
rect 12027 24160 12072 24188
rect 11609 24151 11667 24157
rect 5258 24120 5264 24132
rect 5219 24092 5264 24120
rect 5258 24080 5264 24092
rect 5316 24120 5322 24132
rect 5316 24092 11468 24120
rect 5316 24080 5322 24092
rect 3234 24052 3240 24064
rect 3195 24024 3240 24052
rect 3234 24012 3240 24024
rect 3292 24012 3298 24064
rect 10686 24052 10692 24064
rect 10647 24024 10692 24052
rect 10686 24012 10692 24024
rect 10744 24012 10750 24064
rect 11440 24061 11468 24092
rect 11425 24055 11483 24061
rect 11425 24021 11437 24055
rect 11471 24052 11483 24055
rect 11514 24052 11520 24064
rect 11471 24024 11520 24052
rect 11471 24021 11483 24024
rect 11425 24015 11483 24021
rect 11514 24012 11520 24024
rect 11572 24012 11578 24064
rect 11624 24052 11652 24151
rect 12066 24148 12072 24160
rect 12124 24148 12130 24200
rect 15740 24191 15798 24197
rect 15740 24157 15752 24191
rect 15786 24188 15798 24191
rect 16114 24188 16120 24200
rect 15786 24160 16120 24188
rect 15786 24157 15798 24160
rect 15740 24151 15798 24157
rect 16114 24148 16120 24160
rect 16172 24148 16178 24200
rect 17310 24188 17316 24200
rect 17223 24160 17316 24188
rect 17310 24148 17316 24160
rect 17368 24148 17374 24200
rect 17580 24191 17638 24197
rect 17580 24157 17592 24191
rect 17626 24188 17638 24191
rect 18690 24188 18696 24200
rect 17626 24160 18696 24188
rect 17626 24157 17638 24160
rect 17580 24151 17638 24157
rect 18690 24148 18696 24160
rect 18748 24148 18754 24200
rect 19429 24191 19487 24197
rect 19429 24157 19441 24191
rect 19475 24157 19487 24191
rect 19429 24151 19487 24157
rect 19696 24191 19754 24197
rect 19696 24157 19708 24191
rect 19742 24188 19754 24191
rect 21174 24188 21180 24200
rect 19742 24160 21180 24188
rect 19742 24157 19754 24160
rect 19696 24151 19754 24157
rect 12336 24123 12394 24129
rect 12336 24089 12348 24123
rect 12382 24120 12394 24123
rect 13262 24120 13268 24132
rect 12382 24092 13268 24120
rect 12382 24089 12394 24092
rect 12336 24083 12394 24089
rect 13262 24080 13268 24092
rect 13320 24080 13326 24132
rect 17328 24120 17356 24148
rect 19334 24120 19340 24132
rect 17328 24092 19340 24120
rect 19334 24080 19340 24092
rect 19392 24120 19398 24132
rect 19444 24120 19472 24151
rect 21174 24148 21180 24160
rect 21232 24148 21238 24200
rect 21269 24191 21327 24197
rect 21269 24157 21281 24191
rect 21315 24188 21327 24191
rect 21818 24188 21824 24200
rect 21315 24160 21824 24188
rect 21315 24157 21327 24160
rect 21269 24151 21327 24157
rect 21284 24120 21312 24151
rect 21818 24148 21824 24160
rect 21876 24188 21882 24200
rect 24397 24191 24455 24197
rect 24397 24188 24409 24191
rect 21876 24160 24409 24188
rect 21876 24148 21882 24160
rect 24397 24157 24409 24160
rect 24443 24157 24455 24191
rect 24397 24151 24455 24157
rect 24486 24148 24492 24200
rect 24544 24188 24550 24200
rect 24653 24191 24711 24197
rect 24653 24188 24665 24191
rect 24544 24160 24665 24188
rect 24544 24148 24550 24160
rect 24653 24157 24665 24160
rect 24699 24157 24711 24191
rect 24653 24151 24711 24157
rect 26234 24148 26240 24200
rect 26292 24188 26298 24200
rect 26504 24191 26562 24197
rect 26292 24160 26337 24188
rect 26292 24148 26298 24160
rect 26504 24157 26516 24191
rect 26550 24188 26562 24191
rect 27614 24188 27620 24200
rect 26550 24160 27620 24188
rect 26550 24157 26562 24160
rect 26504 24151 26562 24157
rect 27614 24148 27620 24160
rect 27672 24148 27678 24200
rect 29549 24191 29607 24197
rect 29549 24157 29561 24191
rect 29595 24188 29607 24191
rect 30282 24188 30288 24200
rect 29595 24160 30288 24188
rect 29595 24157 29607 24160
rect 29549 24151 29607 24157
rect 30282 24148 30288 24160
rect 30340 24148 30346 24200
rect 19392 24092 21312 24120
rect 21536 24123 21594 24129
rect 19392 24080 19398 24092
rect 21536 24089 21548 24123
rect 21582 24120 21594 24123
rect 23106 24120 23112 24132
rect 21582 24092 23112 24120
rect 21582 24089 21594 24092
rect 21536 24083 21594 24089
rect 23106 24080 23112 24092
rect 23164 24080 23170 24132
rect 29816 24123 29874 24129
rect 29816 24089 29828 24123
rect 29862 24120 29874 24123
rect 30926 24120 30932 24132
rect 29862 24092 30932 24120
rect 29862 24089 29874 24092
rect 29816 24083 29874 24089
rect 30926 24080 30932 24092
rect 30984 24080 30990 24132
rect 31202 24080 31208 24132
rect 31260 24120 31266 24132
rect 31634 24123 31692 24129
rect 31634 24120 31646 24123
rect 31260 24092 31646 24120
rect 31260 24080 31266 24092
rect 31634 24089 31646 24092
rect 31680 24089 31692 24123
rect 34716 24120 34744 24219
rect 41414 24216 41420 24268
rect 41472 24256 41478 24268
rect 41708 24265 41736 24364
rect 42426 24352 42432 24364
rect 42484 24352 42490 24404
rect 43070 24392 43076 24404
rect 43031 24364 43076 24392
rect 43070 24352 43076 24364
rect 43128 24352 43134 24404
rect 48958 24392 48964 24404
rect 48919 24364 48964 24392
rect 48958 24352 48964 24364
rect 49016 24352 49022 24404
rect 54110 24392 54116 24404
rect 53116 24364 54116 24392
rect 41693 24259 41751 24265
rect 41693 24256 41705 24259
rect 41472 24228 41705 24256
rect 41472 24216 41478 24228
rect 41693 24225 41705 24228
rect 41739 24225 41751 24259
rect 41693 24219 41751 24225
rect 44910 24216 44916 24268
rect 44968 24256 44974 24268
rect 53116 24265 53144 24364
rect 54110 24352 54116 24364
rect 54168 24392 54174 24404
rect 56502 24392 56508 24404
rect 54168 24364 56508 24392
rect 54168 24352 54174 24364
rect 55324 24265 55352 24364
rect 56502 24352 56508 24364
rect 56560 24352 56566 24404
rect 56689 24395 56747 24401
rect 56689 24361 56701 24395
rect 56735 24392 56747 24395
rect 56778 24392 56784 24404
rect 56735 24364 56784 24392
rect 56735 24361 56747 24364
rect 56689 24355 56747 24361
rect 56778 24352 56784 24364
rect 56836 24352 56842 24404
rect 59541 24395 59599 24401
rect 59541 24392 59553 24395
rect 57072 24364 59553 24392
rect 45005 24259 45063 24265
rect 45005 24256 45017 24259
rect 44968 24228 45017 24256
rect 44968 24216 44974 24228
rect 45005 24225 45017 24228
rect 45051 24225 45063 24259
rect 45005 24219 45063 24225
rect 53101 24259 53159 24265
rect 53101 24225 53113 24259
rect 53147 24225 53159 24259
rect 53101 24219 53159 24225
rect 55309 24259 55367 24265
rect 55309 24225 55321 24259
rect 55355 24225 55367 24259
rect 55309 24219 55367 24225
rect 34968 24191 35026 24197
rect 34968 24157 34980 24191
rect 35014 24188 35026 24191
rect 36078 24188 36084 24200
rect 35014 24160 36084 24188
rect 35014 24157 35026 24160
rect 34968 24151 35026 24157
rect 36078 24148 36084 24160
rect 36136 24148 36142 24200
rect 36541 24191 36599 24197
rect 36541 24157 36553 24191
rect 36587 24157 36599 24191
rect 36541 24151 36599 24157
rect 36808 24191 36866 24197
rect 36808 24157 36820 24191
rect 36854 24188 36866 24191
rect 39022 24188 39028 24200
rect 36854 24160 39028 24188
rect 36854 24157 36866 24160
rect 36808 24151 36866 24157
rect 35342 24120 35348 24132
rect 34716 24092 35348 24120
rect 31634 24083 31692 24089
rect 35342 24080 35348 24092
rect 35400 24120 35406 24132
rect 36556 24120 36584 24151
rect 39022 24148 39028 24160
rect 39080 24148 39086 24200
rect 39850 24188 39856 24200
rect 39763 24160 39856 24188
rect 39850 24148 39856 24160
rect 39908 24148 39914 24200
rect 40120 24191 40178 24197
rect 40120 24157 40132 24191
rect 40166 24188 40178 24191
rect 41230 24188 41236 24200
rect 40166 24160 41236 24188
rect 40166 24157 40178 24160
rect 40120 24151 40178 24157
rect 41230 24148 41236 24160
rect 41288 24148 41294 24200
rect 41960 24191 42018 24197
rect 41960 24157 41972 24191
rect 42006 24188 42018 24191
rect 43806 24188 43812 24200
rect 42006 24160 43812 24188
rect 42006 24157 42018 24160
rect 41960 24151 42018 24157
rect 43806 24148 43812 24160
rect 43864 24148 43870 24200
rect 47578 24188 47584 24200
rect 47539 24160 47584 24188
rect 47578 24148 47584 24160
rect 47636 24148 47642 24200
rect 48314 24148 48320 24200
rect 48372 24188 48378 24200
rect 49605 24191 49663 24197
rect 49605 24188 49617 24191
rect 48372 24160 49617 24188
rect 48372 24148 48378 24160
rect 49605 24157 49617 24160
rect 49651 24157 49663 24191
rect 50154 24188 50160 24200
rect 50115 24160 50160 24188
rect 49605 24151 49663 24157
rect 50154 24148 50160 24160
rect 50212 24148 50218 24200
rect 55576 24191 55634 24197
rect 55576 24157 55588 24191
rect 55622 24188 55634 24191
rect 57072 24188 57100 24364
rect 59541 24361 59553 24364
rect 59587 24361 59599 24395
rect 59541 24355 59599 24361
rect 55622 24160 57100 24188
rect 57149 24191 57207 24197
rect 55622 24157 55634 24160
rect 55576 24151 55634 24157
rect 57149 24157 57161 24191
rect 57195 24157 57207 24191
rect 57149 24151 57207 24157
rect 35400 24092 36584 24120
rect 39868 24120 39896 24148
rect 41414 24120 41420 24132
rect 39868 24092 41420 24120
rect 35400 24080 35406 24092
rect 41414 24080 41420 24092
rect 41472 24080 41478 24132
rect 45272 24123 45330 24129
rect 45272 24089 45284 24123
rect 45318 24120 45330 24123
rect 46842 24120 46848 24132
rect 45318 24092 46848 24120
rect 45318 24089 45330 24092
rect 45272 24083 45330 24089
rect 46842 24080 46848 24092
rect 46900 24080 46906 24132
rect 47848 24123 47906 24129
rect 47848 24089 47860 24123
rect 47894 24120 47906 24123
rect 48866 24120 48872 24132
rect 47894 24092 48872 24120
rect 47894 24089 47906 24092
rect 47848 24083 47906 24089
rect 48866 24080 48872 24092
rect 48924 24080 48930 24132
rect 50424 24123 50482 24129
rect 50424 24089 50436 24123
rect 50470 24120 50482 24123
rect 50798 24120 50804 24132
rect 50470 24092 50804 24120
rect 50470 24089 50482 24092
rect 50424 24083 50482 24089
rect 50798 24080 50804 24092
rect 50856 24080 50862 24132
rect 53368 24123 53426 24129
rect 53368 24089 53380 24123
rect 53414 24120 53426 24123
rect 53414 24092 55214 24120
rect 53414 24089 53426 24092
rect 53368 24083 53426 24089
rect 14090 24052 14096 24064
rect 11624 24024 14096 24052
rect 14090 24012 14096 24024
rect 14148 24012 14154 24064
rect 16850 24052 16856 24064
rect 16811 24024 16856 24052
rect 16850 24012 16856 24024
rect 16908 24012 16914 24064
rect 18690 24052 18696 24064
rect 18651 24024 18696 24052
rect 18690 24012 18696 24024
rect 18748 24012 18754 24064
rect 20806 24052 20812 24064
rect 20767 24024 20812 24052
rect 20806 24012 20812 24024
rect 20864 24012 20870 24064
rect 22646 24052 22652 24064
rect 22607 24024 22652 24052
rect 22646 24012 22652 24024
rect 22704 24012 22710 24064
rect 27614 24052 27620 24064
rect 27575 24024 27620 24052
rect 27614 24012 27620 24024
rect 27672 24012 27678 24064
rect 36078 24052 36084 24064
rect 36039 24024 36084 24052
rect 36078 24012 36084 24024
rect 36136 24012 36142 24064
rect 46382 24052 46388 24064
rect 46343 24024 46388 24052
rect 46382 24012 46388 24024
rect 46440 24012 46446 24064
rect 49418 24052 49424 24064
rect 49331 24024 49424 24052
rect 49418 24012 49424 24024
rect 49476 24052 49482 24064
rect 49970 24052 49976 24064
rect 49476 24024 49976 24052
rect 49476 24012 49482 24024
rect 49970 24012 49976 24024
rect 50028 24012 50034 24064
rect 51534 24052 51540 24064
rect 51495 24024 51540 24052
rect 51534 24012 51540 24024
rect 51592 24012 51598 24064
rect 54478 24052 54484 24064
rect 54439 24024 54484 24052
rect 54478 24012 54484 24024
rect 54536 24012 54542 24064
rect 55186 24052 55214 24092
rect 56778 24080 56784 24132
rect 56836 24120 56842 24132
rect 57164 24120 57192 24151
rect 56836 24092 57192 24120
rect 56836 24080 56842 24092
rect 57238 24080 57244 24132
rect 57296 24120 57302 24132
rect 57394 24123 57452 24129
rect 57394 24120 57406 24123
rect 57296 24092 57406 24120
rect 57296 24080 57302 24092
rect 57394 24089 57406 24092
rect 57440 24089 57452 24123
rect 59449 24123 59507 24129
rect 59449 24120 59461 24123
rect 57394 24083 57452 24089
rect 57532 24092 59461 24120
rect 57532 24052 57560 24092
rect 59449 24089 59461 24092
rect 59495 24089 59507 24123
rect 59449 24083 59507 24089
rect 58526 24052 58532 24064
rect 55186 24024 57560 24052
rect 58487 24024 58532 24052
rect 58526 24012 58532 24024
rect 58584 24012 58590 24064
rect 1104 23962 59340 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 59340 23962
rect 1104 23888 59340 23910
rect 5813 23851 5871 23857
rect 5813 23817 5825 23851
rect 5859 23848 5871 23851
rect 6086 23848 6092 23860
rect 5859 23820 6092 23848
rect 5859 23817 5871 23820
rect 5813 23811 5871 23817
rect 6086 23808 6092 23820
rect 6144 23808 6150 23860
rect 13262 23848 13268 23860
rect 13223 23820 13268 23848
rect 13262 23808 13268 23820
rect 13320 23808 13326 23860
rect 14090 23808 14096 23860
rect 14148 23848 14154 23860
rect 14148 23820 19196 23848
rect 14148 23808 14154 23820
rect 2584 23783 2642 23789
rect 2584 23749 2596 23783
rect 2630 23780 2642 23783
rect 3234 23780 3240 23792
rect 2630 23752 3240 23780
rect 2630 23749 2642 23752
rect 2584 23743 2642 23749
rect 3234 23740 3240 23752
rect 3292 23740 3298 23792
rect 9668 23783 9726 23789
rect 9668 23749 9680 23783
rect 9714 23780 9726 23783
rect 10686 23780 10692 23792
rect 9714 23752 10692 23780
rect 9714 23749 9726 23752
rect 9668 23743 9726 23749
rect 10686 23740 10692 23752
rect 10744 23740 10750 23792
rect 17672 23783 17730 23789
rect 17672 23749 17684 23783
rect 17718 23780 17730 23783
rect 18690 23780 18696 23792
rect 17718 23752 18696 23780
rect 17718 23749 17730 23752
rect 17672 23743 17730 23749
rect 18690 23740 18696 23752
rect 18748 23740 18754 23792
rect 19168 23780 19196 23820
rect 19242 23808 19248 23860
rect 19300 23848 19306 23860
rect 20625 23851 20683 23857
rect 20625 23848 20637 23851
rect 19300 23820 20637 23848
rect 19300 23808 19306 23820
rect 20625 23817 20637 23820
rect 20671 23817 20683 23851
rect 23198 23848 23204 23860
rect 23159 23820 23204 23848
rect 20625 23811 20683 23817
rect 23198 23808 23204 23820
rect 23256 23808 23262 23860
rect 25498 23848 25504 23860
rect 25459 23820 25504 23848
rect 25498 23808 25504 23820
rect 25556 23808 25562 23860
rect 28350 23848 28356 23860
rect 28311 23820 28356 23848
rect 28350 23808 28356 23820
rect 28408 23808 28414 23860
rect 33505 23851 33563 23857
rect 33505 23817 33517 23851
rect 33551 23848 33563 23851
rect 34514 23848 34520 23860
rect 33551 23820 34520 23848
rect 33551 23817 33563 23820
rect 33505 23811 33563 23817
rect 34514 23808 34520 23820
rect 34572 23808 34578 23860
rect 35345 23851 35403 23857
rect 35345 23817 35357 23851
rect 35391 23848 35403 23851
rect 36170 23848 36176 23860
rect 35391 23820 36176 23848
rect 35391 23817 35403 23820
rect 35345 23811 35403 23817
rect 36170 23808 36176 23820
rect 36228 23808 36234 23860
rect 41877 23851 41935 23857
rect 41877 23817 41889 23851
rect 41923 23817 41935 23851
rect 41877 23811 41935 23817
rect 19512 23783 19570 23789
rect 19168 23752 19472 23780
rect 2222 23672 2228 23724
rect 2280 23712 2286 23724
rect 2317 23715 2375 23721
rect 2317 23712 2329 23715
rect 2280 23684 2329 23712
rect 2280 23672 2286 23684
rect 2317 23681 2329 23684
rect 2363 23712 2375 23715
rect 4700 23715 4758 23721
rect 2363 23684 4476 23712
rect 2363 23681 2375 23684
rect 2317 23675 2375 23681
rect 4448 23653 4476 23684
rect 4700 23681 4712 23715
rect 4746 23712 4758 23715
rect 6546 23712 6552 23724
rect 4746 23684 6552 23712
rect 4746 23681 4758 23684
rect 4700 23675 4758 23681
rect 6546 23672 6552 23684
rect 6604 23672 6610 23724
rect 7828 23715 7886 23721
rect 7828 23681 7840 23715
rect 7874 23712 7886 23715
rect 9306 23712 9312 23724
rect 7874 23684 9312 23712
rect 7874 23681 7886 23684
rect 7828 23675 7886 23681
rect 9306 23672 9312 23684
rect 9364 23672 9370 23724
rect 12152 23715 12210 23721
rect 12152 23681 12164 23715
rect 12198 23712 12210 23715
rect 13078 23712 13084 23724
rect 12198 23684 13084 23712
rect 12198 23681 12210 23684
rect 12152 23675 12210 23681
rect 13078 23672 13084 23684
rect 13136 23672 13142 23724
rect 15004 23715 15062 23721
rect 15004 23681 15016 23715
rect 15050 23712 15062 23715
rect 15746 23712 15752 23724
rect 15050 23684 15752 23712
rect 15050 23681 15062 23684
rect 15004 23675 15062 23681
rect 15746 23672 15752 23684
rect 15804 23672 15810 23724
rect 19245 23715 19303 23721
rect 19245 23681 19257 23715
rect 19291 23712 19303 23715
rect 19334 23712 19340 23724
rect 19291 23684 19340 23712
rect 19291 23681 19303 23684
rect 19245 23675 19303 23681
rect 19334 23672 19340 23684
rect 19392 23672 19398 23724
rect 19444 23712 19472 23752
rect 19512 23749 19524 23783
rect 19558 23780 19570 23783
rect 20806 23780 20812 23792
rect 19558 23752 20812 23780
rect 19558 23749 19570 23752
rect 19512 23743 19570 23749
rect 20806 23740 20812 23752
rect 20864 23740 20870 23792
rect 22088 23783 22146 23789
rect 22088 23749 22100 23783
rect 22134 23780 22146 23783
rect 22646 23780 22652 23792
rect 22134 23752 22652 23780
rect 22134 23749 22146 23752
rect 22088 23743 22146 23749
rect 22646 23740 22652 23752
rect 22704 23740 22710 23792
rect 27240 23783 27298 23789
rect 27240 23749 27252 23783
rect 27286 23780 27298 23783
rect 27614 23780 27620 23792
rect 27286 23752 27620 23780
rect 27286 23749 27298 23752
rect 27240 23743 27298 23749
rect 27614 23740 27620 23752
rect 27672 23740 27678 23792
rect 29086 23789 29092 23792
rect 29080 23780 29092 23789
rect 29047 23752 29092 23780
rect 29080 23743 29092 23752
rect 29086 23740 29092 23743
rect 29144 23740 29150 23792
rect 32398 23789 32404 23792
rect 32392 23780 32404 23789
rect 32359 23752 32404 23780
rect 32392 23743 32404 23752
rect 32398 23740 32404 23743
rect 32456 23740 32462 23792
rect 34232 23783 34290 23789
rect 34232 23749 34244 23783
rect 34278 23780 34290 23783
rect 36078 23780 36084 23792
rect 34278 23752 36084 23780
rect 34278 23749 34290 23752
rect 34232 23743 34290 23749
rect 36078 23740 36084 23752
rect 36136 23740 36142 23792
rect 41892 23780 41920 23811
rect 48866 23808 48872 23860
rect 48924 23848 48930 23860
rect 48961 23851 49019 23857
rect 48961 23848 48973 23851
rect 48924 23820 48973 23848
rect 48924 23808 48930 23820
rect 48961 23817 48973 23820
rect 49007 23817 49019 23851
rect 50798 23848 50804 23860
rect 50759 23820 50804 23848
rect 48961 23811 49019 23817
rect 50798 23808 50804 23820
rect 50856 23808 50862 23860
rect 54754 23848 54760 23860
rect 54715 23820 54760 23848
rect 54754 23808 54760 23820
rect 54812 23808 54818 23860
rect 57330 23848 57336 23860
rect 57291 23820 57336 23848
rect 57330 23808 57336 23820
rect 57388 23808 57394 23860
rect 45922 23789 45928 23792
rect 45916 23780 45928 23789
rect 38764 23752 41920 23780
rect 45883 23752 45928 23780
rect 20990 23712 20996 23724
rect 19444 23684 20996 23712
rect 20990 23672 20996 23684
rect 21048 23672 21054 23724
rect 21818 23712 21824 23724
rect 21779 23684 21824 23712
rect 21818 23672 21824 23684
rect 21876 23672 21882 23724
rect 24388 23715 24446 23721
rect 24388 23681 24400 23715
rect 24434 23712 24446 23715
rect 25774 23712 25780 23724
rect 24434 23684 25780 23712
rect 24434 23681 24446 23684
rect 24388 23675 24446 23681
rect 25774 23672 25780 23684
rect 25832 23672 25838 23724
rect 31386 23672 31392 23724
rect 31444 23712 31450 23724
rect 32125 23715 32183 23721
rect 32125 23712 32137 23715
rect 31444 23684 32137 23712
rect 31444 23672 31450 23684
rect 32125 23681 32137 23684
rect 32171 23712 32183 23715
rect 32171 23684 33180 23712
rect 32171 23681 32183 23684
rect 32125 23675 32183 23681
rect 4433 23647 4491 23653
rect 4433 23613 4445 23647
rect 4479 23613 4491 23647
rect 4433 23607 4491 23613
rect 3694 23508 3700 23520
rect 3655 23480 3700 23508
rect 3694 23468 3700 23480
rect 3752 23468 3758 23520
rect 4448 23508 4476 23607
rect 7006 23604 7012 23656
rect 7064 23644 7070 23656
rect 7561 23647 7619 23653
rect 7561 23644 7573 23647
rect 7064 23616 7573 23644
rect 7064 23604 7070 23616
rect 7561 23613 7573 23616
rect 7607 23613 7619 23647
rect 7561 23607 7619 23613
rect 9214 23604 9220 23656
rect 9272 23644 9278 23656
rect 9401 23647 9459 23653
rect 9401 23644 9413 23647
rect 9272 23616 9413 23644
rect 9272 23604 9278 23616
rect 9401 23613 9413 23616
rect 9447 23613 9459 23647
rect 9401 23607 9459 23613
rect 11885 23647 11943 23653
rect 11885 23613 11897 23647
rect 11931 23613 11943 23647
rect 11885 23607 11943 23613
rect 5166 23508 5172 23520
rect 4448 23480 5172 23508
rect 5166 23468 5172 23480
rect 5224 23468 5230 23520
rect 8938 23508 8944 23520
rect 8899 23480 8944 23508
rect 8938 23468 8944 23480
rect 8996 23468 9002 23520
rect 10778 23508 10784 23520
rect 10739 23480 10784 23508
rect 10778 23468 10784 23480
rect 10836 23468 10842 23520
rect 11900 23508 11928 23607
rect 13814 23604 13820 23656
rect 13872 23644 13878 23656
rect 14734 23644 14740 23656
rect 13872 23616 14740 23644
rect 13872 23604 13878 23616
rect 14734 23604 14740 23616
rect 14792 23604 14798 23656
rect 17405 23647 17463 23653
rect 17405 23644 17417 23647
rect 16546 23616 17417 23644
rect 16546 23576 16574 23616
rect 17405 23613 17417 23616
rect 17451 23613 17463 23647
rect 24118 23644 24124 23656
rect 24079 23616 24124 23644
rect 17405 23607 17463 23613
rect 15672 23548 16574 23576
rect 12066 23508 12072 23520
rect 11900 23480 12072 23508
rect 12066 23468 12072 23480
rect 12124 23508 12130 23520
rect 12250 23508 12256 23520
rect 12124 23480 12256 23508
rect 12124 23468 12130 23480
rect 12250 23468 12256 23480
rect 12308 23468 12314 23520
rect 15470 23468 15476 23520
rect 15528 23508 15534 23520
rect 15672 23508 15700 23548
rect 15528 23480 15700 23508
rect 15528 23468 15534 23480
rect 16022 23468 16028 23520
rect 16080 23508 16086 23520
rect 16117 23511 16175 23517
rect 16117 23508 16129 23511
rect 16080 23480 16129 23508
rect 16080 23468 16086 23480
rect 16117 23477 16129 23480
rect 16163 23477 16175 23511
rect 17420 23508 17448 23607
rect 24118 23604 24124 23616
rect 24176 23604 24182 23656
rect 26234 23604 26240 23656
rect 26292 23644 26298 23656
rect 26973 23647 27031 23653
rect 26973 23644 26985 23647
rect 26292 23616 26985 23644
rect 26292 23604 26298 23616
rect 26973 23613 26985 23616
rect 27019 23613 27031 23647
rect 26973 23607 27031 23613
rect 28813 23647 28871 23653
rect 28813 23613 28825 23647
rect 28859 23613 28871 23647
rect 33152 23644 33180 23684
rect 33594 23672 33600 23724
rect 33652 23712 33658 23724
rect 38764 23712 38792 23752
rect 45916 23743 45928 23752
rect 45922 23740 45928 23743
rect 45980 23740 45986 23792
rect 49694 23789 49700 23792
rect 49688 23780 49700 23789
rect 49655 23752 49700 23780
rect 49688 23743 49700 23752
rect 49694 23740 49700 23743
rect 49752 23740 49758 23792
rect 53644 23783 53702 23789
rect 53644 23749 53656 23783
rect 53690 23780 53702 23783
rect 54478 23780 54484 23792
rect 53690 23752 54484 23780
rect 53690 23749 53702 23752
rect 53644 23743 53702 23749
rect 54478 23740 54484 23752
rect 54536 23740 54542 23792
rect 56220 23783 56278 23789
rect 56220 23749 56232 23783
rect 56266 23780 56278 23783
rect 58526 23780 58532 23792
rect 56266 23752 58532 23780
rect 56266 23749 56278 23752
rect 56220 23743 56278 23749
rect 58526 23740 58532 23752
rect 58584 23740 58590 23792
rect 33652 23684 38792 23712
rect 38832 23715 38890 23721
rect 33652 23672 33658 23684
rect 38832 23681 38844 23715
rect 38878 23712 38890 23715
rect 40034 23712 40040 23724
rect 38878 23684 40040 23712
rect 38878 23681 38890 23684
rect 38832 23675 38890 23681
rect 40034 23672 40040 23684
rect 40092 23672 40098 23724
rect 40764 23715 40822 23721
rect 40764 23681 40776 23715
rect 40810 23712 40822 23715
rect 41690 23712 41696 23724
rect 40810 23684 41696 23712
rect 40810 23681 40822 23684
rect 40764 23675 40822 23681
rect 41690 23672 41696 23684
rect 41748 23672 41754 23724
rect 44076 23715 44134 23721
rect 44076 23681 44088 23715
rect 44122 23712 44134 23715
rect 44818 23712 44824 23724
rect 44122 23684 44824 23712
rect 44122 23681 44134 23684
rect 44076 23675 44134 23681
rect 44818 23672 44824 23684
rect 44876 23672 44882 23724
rect 47578 23712 47584 23724
rect 45664 23684 47584 23712
rect 33962 23644 33968 23656
rect 33152 23616 33968 23644
rect 28813 23607 28871 23613
rect 18046 23508 18052 23520
rect 17420 23480 18052 23508
rect 16117 23471 16175 23477
rect 18046 23468 18052 23480
rect 18104 23468 18110 23520
rect 18782 23508 18788 23520
rect 18743 23480 18788 23508
rect 18782 23468 18788 23480
rect 18840 23468 18846 23520
rect 26988 23508 27016 23607
rect 27614 23508 27620 23520
rect 26988 23480 27620 23508
rect 27614 23468 27620 23480
rect 27672 23508 27678 23520
rect 28828 23508 28856 23607
rect 33962 23604 33968 23616
rect 34020 23604 34026 23656
rect 37642 23604 37648 23656
rect 37700 23644 37706 23656
rect 38565 23647 38623 23653
rect 38565 23644 38577 23647
rect 37700 23616 38577 23644
rect 37700 23604 37706 23616
rect 38565 23613 38577 23616
rect 38611 23613 38623 23647
rect 38565 23607 38623 23613
rect 40497 23647 40555 23653
rect 40497 23613 40509 23647
rect 40543 23613 40555 23647
rect 40497 23607 40555 23613
rect 30190 23508 30196 23520
rect 27672 23480 28856 23508
rect 30151 23480 30196 23508
rect 27672 23468 27678 23480
rect 30190 23468 30196 23480
rect 30248 23468 30254 23520
rect 38194 23468 38200 23520
rect 38252 23508 38258 23520
rect 39945 23511 40003 23517
rect 39945 23508 39957 23511
rect 38252 23480 39957 23508
rect 38252 23468 38258 23480
rect 39945 23477 39957 23480
rect 39991 23477 40003 23511
rect 40512 23508 40540 23607
rect 43070 23604 43076 23656
rect 43128 23644 43134 23656
rect 43809 23647 43867 23653
rect 43809 23644 43821 23647
rect 43128 23616 43821 23644
rect 43128 23604 43134 23616
rect 43809 23613 43821 23616
rect 43855 23613 43867 23647
rect 43809 23607 43867 23613
rect 45554 23604 45560 23656
rect 45612 23644 45618 23656
rect 45664 23653 45692 23684
rect 47578 23672 47584 23684
rect 47636 23672 47642 23724
rect 47848 23715 47906 23721
rect 47848 23681 47860 23715
rect 47894 23712 47906 23715
rect 49326 23712 49332 23724
rect 47894 23684 49332 23712
rect 47894 23681 47906 23684
rect 47848 23675 47906 23681
rect 49326 23672 49332 23684
rect 49384 23672 49390 23724
rect 49421 23715 49479 23721
rect 49421 23681 49433 23715
rect 49467 23712 49479 23715
rect 49510 23712 49516 23724
rect 49467 23684 49516 23712
rect 49467 23681 49479 23684
rect 49421 23675 49479 23681
rect 49510 23672 49516 23684
rect 49568 23712 49574 23724
rect 50154 23712 50160 23724
rect 49568 23684 50160 23712
rect 49568 23672 49574 23684
rect 50154 23672 50160 23684
rect 50212 23672 50218 23724
rect 53374 23712 53380 23724
rect 53287 23684 53380 23712
rect 53374 23672 53380 23684
rect 53432 23712 53438 23724
rect 55953 23715 56011 23721
rect 55953 23712 55965 23715
rect 53432 23684 55965 23712
rect 53432 23672 53438 23684
rect 55953 23681 55965 23684
rect 55999 23712 56011 23715
rect 56778 23712 56784 23724
rect 55999 23684 56784 23712
rect 55999 23681 56011 23684
rect 55953 23675 56011 23681
rect 56778 23672 56784 23684
rect 56836 23672 56842 23724
rect 45649 23647 45707 23653
rect 45649 23644 45661 23647
rect 45612 23616 45661 23644
rect 45612 23604 45618 23616
rect 45649 23613 45661 23616
rect 45695 23613 45707 23647
rect 45649 23607 45707 23613
rect 41414 23508 41420 23520
rect 40512 23480 41420 23508
rect 39945 23471 40003 23477
rect 41414 23468 41420 23480
rect 41472 23468 41478 23520
rect 45186 23508 45192 23520
rect 45147 23480 45192 23508
rect 45186 23468 45192 23480
rect 45244 23468 45250 23520
rect 47026 23508 47032 23520
rect 46987 23480 47032 23508
rect 47026 23468 47032 23480
rect 47084 23468 47090 23520
rect 1104 23418 59340 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 59340 23418
rect 1104 23344 59340 23366
rect 6546 23304 6552 23316
rect 6507 23276 6552 23304
rect 6546 23264 6552 23276
rect 6604 23264 6610 23316
rect 8018 23264 8024 23316
rect 8076 23304 8082 23316
rect 8389 23307 8447 23313
rect 8389 23304 8401 23307
rect 8076 23276 8401 23304
rect 8076 23264 8082 23276
rect 8389 23273 8401 23276
rect 8435 23273 8447 23307
rect 8389 23267 8447 23273
rect 15746 23264 15752 23316
rect 15804 23304 15810 23316
rect 16853 23307 16911 23313
rect 16853 23304 16865 23307
rect 15804 23276 16865 23304
rect 15804 23264 15810 23276
rect 16853 23273 16865 23276
rect 16899 23273 16911 23307
rect 16853 23267 16911 23273
rect 18506 23264 18512 23316
rect 18564 23304 18570 23316
rect 18693 23307 18751 23313
rect 18693 23304 18705 23307
rect 18564 23276 18705 23304
rect 18564 23264 18570 23276
rect 18693 23273 18705 23276
rect 18739 23273 18751 23307
rect 25774 23304 25780 23316
rect 25735 23276 25780 23304
rect 18693 23267 18751 23273
rect 25774 23264 25780 23276
rect 25832 23264 25838 23316
rect 27617 23307 27675 23313
rect 27617 23273 27629 23307
rect 27663 23304 27675 23307
rect 27706 23304 27712 23316
rect 27663 23276 27712 23304
rect 27663 23273 27675 23276
rect 27617 23267 27675 23273
rect 27706 23264 27712 23276
rect 27764 23264 27770 23316
rect 40586 23264 40592 23316
rect 40644 23304 40650 23316
rect 40644 23276 46796 23304
rect 40644 23264 40650 23276
rect 46768 23236 46796 23276
rect 46842 23264 46848 23316
rect 46900 23304 46906 23316
rect 46937 23307 46995 23313
rect 46937 23304 46949 23307
rect 46900 23276 46949 23304
rect 46900 23264 46906 23276
rect 46937 23273 46949 23276
rect 46983 23273 46995 23307
rect 48314 23304 48320 23316
rect 46937 23267 46995 23273
rect 47044 23276 48320 23304
rect 47044 23236 47072 23276
rect 48314 23264 48320 23276
rect 48372 23264 48378 23316
rect 49326 23304 49332 23316
rect 49287 23276 49332 23304
rect 49326 23264 49332 23276
rect 49384 23264 49390 23316
rect 46768 23208 47072 23236
rect 5166 23168 5172 23180
rect 5127 23140 5172 23168
rect 5166 23128 5172 23140
rect 5224 23128 5230 23180
rect 12250 23128 12256 23180
rect 12308 23168 12314 23180
rect 13541 23171 13599 23177
rect 13541 23168 13553 23171
rect 12308 23140 13553 23168
rect 12308 23128 12314 23140
rect 13541 23137 13553 23140
rect 13587 23168 13599 23171
rect 13722 23168 13728 23180
rect 13587 23140 13728 23168
rect 13587 23137 13599 23140
rect 13541 23131 13599 23137
rect 13722 23128 13728 23140
rect 13780 23128 13786 23180
rect 15470 23168 15476 23180
rect 15431 23140 15476 23168
rect 15470 23128 15476 23140
rect 15528 23128 15534 23180
rect 17310 23168 17316 23180
rect 17271 23140 17316 23168
rect 17310 23128 17316 23140
rect 17368 23128 17374 23180
rect 30374 23128 30380 23180
rect 30432 23168 30438 23180
rect 30834 23168 30840 23180
rect 30432 23140 30840 23168
rect 30432 23128 30438 23140
rect 30834 23128 30840 23140
rect 30892 23168 30898 23180
rect 30929 23171 30987 23177
rect 30929 23168 30941 23171
rect 30892 23140 30941 23168
rect 30892 23128 30898 23140
rect 30929 23137 30941 23140
rect 30975 23137 30987 23171
rect 30929 23131 30987 23137
rect 1857 23103 1915 23109
rect 1857 23069 1869 23103
rect 1903 23069 1915 23103
rect 1857 23063 1915 23069
rect 2124 23103 2182 23109
rect 2124 23069 2136 23103
rect 2170 23100 2182 23103
rect 3694 23100 3700 23112
rect 2170 23072 3700 23100
rect 2170 23069 2182 23072
rect 2124 23063 2182 23069
rect 1872 23032 1900 23063
rect 3694 23060 3700 23072
rect 3752 23060 3758 23112
rect 5436 23103 5494 23109
rect 5436 23069 5448 23103
rect 5482 23100 5494 23103
rect 6178 23100 6184 23112
rect 5482 23072 6184 23100
rect 5482 23069 5494 23072
rect 5436 23063 5494 23069
rect 6178 23060 6184 23072
rect 6236 23060 6242 23112
rect 7006 23100 7012 23112
rect 6967 23072 7012 23100
rect 7006 23060 7012 23072
rect 7064 23060 7070 23112
rect 7276 23103 7334 23109
rect 7276 23069 7288 23103
rect 7322 23100 7334 23103
rect 8938 23100 8944 23112
rect 7322 23072 8944 23100
rect 7322 23069 7334 23072
rect 7276 23063 7334 23069
rect 8938 23060 8944 23072
rect 8996 23060 9002 23112
rect 9214 23060 9220 23112
rect 9272 23100 9278 23112
rect 9309 23103 9367 23109
rect 9309 23100 9321 23103
rect 9272 23072 9321 23100
rect 9272 23060 9278 23072
rect 9309 23069 9321 23072
rect 9355 23069 9367 23103
rect 9309 23063 9367 23069
rect 9576 23103 9634 23109
rect 9576 23069 9588 23103
rect 9622 23100 9634 23103
rect 10778 23100 10784 23112
rect 9622 23072 10784 23100
rect 9622 23069 9634 23072
rect 9576 23063 9634 23069
rect 10778 23060 10784 23072
rect 10836 23060 10842 23112
rect 15740 23103 15798 23109
rect 15740 23069 15752 23103
rect 15786 23100 15798 23103
rect 16850 23100 16856 23112
rect 15786 23072 16856 23100
rect 15786 23069 15798 23072
rect 15740 23063 15798 23069
rect 16850 23060 16856 23072
rect 16908 23060 16914 23112
rect 17580 23103 17638 23109
rect 17580 23069 17592 23103
rect 17626 23100 17638 23103
rect 18782 23100 18788 23112
rect 17626 23072 18788 23100
rect 17626 23069 17638 23072
rect 17580 23063 17638 23069
rect 18782 23060 18788 23072
rect 18840 23060 18846 23112
rect 19245 23103 19303 23109
rect 19245 23069 19257 23103
rect 19291 23069 19303 23103
rect 21082 23100 21088 23112
rect 21043 23072 21088 23100
rect 19245 23063 19303 23069
rect 2222 23032 2228 23044
rect 1872 23004 2228 23032
rect 2222 22992 2228 23004
rect 2280 22992 2286 23044
rect 11514 22992 11520 23044
rect 11572 23032 11578 23044
rect 11793 23035 11851 23041
rect 11793 23032 11805 23035
rect 11572 23004 11805 23032
rect 11572 22992 11578 23004
rect 11793 23001 11805 23004
rect 11839 23001 11851 23035
rect 11793 22995 11851 23001
rect 18046 22992 18052 23044
rect 18104 23032 18110 23044
rect 19260 23032 19288 23063
rect 21082 23060 21088 23072
rect 21140 23060 21146 23112
rect 24118 23060 24124 23112
rect 24176 23100 24182 23112
rect 24397 23103 24455 23109
rect 24397 23100 24409 23103
rect 24176 23072 24409 23100
rect 24176 23060 24182 23072
rect 24397 23069 24409 23072
rect 24443 23100 24455 23103
rect 26237 23103 26295 23109
rect 26237 23100 26249 23103
rect 24443 23072 26249 23100
rect 24443 23069 24455 23072
rect 24397 23063 24455 23069
rect 26237 23069 26249 23072
rect 26283 23069 26295 23103
rect 26237 23063 26295 23069
rect 26504 23103 26562 23109
rect 26504 23069 26516 23103
rect 26550 23100 26562 23103
rect 27890 23100 27896 23112
rect 26550 23072 27896 23100
rect 26550 23069 26562 23072
rect 26504 23063 26562 23069
rect 18104 23004 19288 23032
rect 19512 23035 19570 23041
rect 18104 22992 18110 23004
rect 19512 23001 19524 23035
rect 19558 23032 19570 23035
rect 21174 23032 21180 23044
rect 19558 23004 21180 23032
rect 19558 23001 19570 23004
rect 19512 22995 19570 23001
rect 21174 22992 21180 23004
rect 21232 22992 21238 23044
rect 21352 23035 21410 23041
rect 21352 23001 21364 23035
rect 21398 23032 21410 23035
rect 22830 23032 22836 23044
rect 21398 23004 22836 23032
rect 21398 23001 21410 23004
rect 21352 22995 21410 23001
rect 22830 22992 22836 23004
rect 22888 22992 22894 23044
rect 24664 23035 24722 23041
rect 24664 23001 24676 23035
rect 24710 23032 24722 23035
rect 25130 23032 25136 23044
rect 24710 23004 25136 23032
rect 24710 23001 24722 23004
rect 24664 22995 24722 23001
rect 25130 22992 25136 23004
rect 25188 22992 25194 23044
rect 26252 23032 26280 23063
rect 27890 23060 27896 23072
rect 27948 23060 27954 23112
rect 30944 23100 30972 23131
rect 47578 23128 47584 23180
rect 47636 23168 47642 23180
rect 47949 23171 48007 23177
rect 47949 23168 47961 23171
rect 47636 23140 47961 23168
rect 47636 23128 47642 23140
rect 47949 23137 47961 23140
rect 47995 23137 48007 23171
rect 47949 23131 48007 23137
rect 32766 23100 32772 23112
rect 30944 23072 32772 23100
rect 32766 23060 32772 23072
rect 32824 23060 32830 23112
rect 35253 23103 35311 23109
rect 35253 23069 35265 23103
rect 35299 23100 35311 23103
rect 36078 23100 36084 23112
rect 35299 23072 36084 23100
rect 35299 23069 35311 23072
rect 35253 23063 35311 23069
rect 36078 23060 36084 23072
rect 36136 23060 36142 23112
rect 37642 23100 37648 23112
rect 37603 23072 37648 23100
rect 37642 23060 37648 23072
rect 37700 23060 37706 23112
rect 40402 23060 40408 23112
rect 40460 23100 40466 23112
rect 40586 23100 40592 23112
rect 40460 23072 40592 23100
rect 40460 23060 40466 23072
rect 40586 23060 40592 23072
rect 40644 23060 40650 23112
rect 41233 23103 41291 23109
rect 41233 23069 41245 23103
rect 41279 23069 41291 23103
rect 43070 23100 43076 23112
rect 43031 23072 43076 23100
rect 41233 23063 41291 23069
rect 27614 23032 27620 23044
rect 26252 23004 27620 23032
rect 27614 22992 27620 23004
rect 27672 22992 27678 23044
rect 31196 23035 31254 23041
rect 31196 23001 31208 23035
rect 31242 23032 31254 23035
rect 31846 23032 31852 23044
rect 31242 23004 31852 23032
rect 31242 23001 31254 23004
rect 31196 22995 31254 23001
rect 31846 22992 31852 23004
rect 31904 22992 31910 23044
rect 33036 23035 33094 23041
rect 33036 23001 33048 23035
rect 33082 23032 33094 23035
rect 34790 23032 34796 23044
rect 33082 23004 34796 23032
rect 33082 23001 33094 23004
rect 33036 22995 33094 23001
rect 34790 22992 34796 23004
rect 34848 22992 34854 23044
rect 35520 23035 35578 23041
rect 35520 23001 35532 23035
rect 35566 23032 35578 23035
rect 36538 23032 36544 23044
rect 35566 23004 36544 23032
rect 35566 23001 35578 23004
rect 35520 22995 35578 23001
rect 36538 22992 36544 23004
rect 36596 22992 36602 23044
rect 37912 23035 37970 23041
rect 37912 23001 37924 23035
rect 37958 23032 37970 23035
rect 39298 23032 39304 23044
rect 37958 23004 39304 23032
rect 37958 23001 37970 23004
rect 37912 22995 37970 23001
rect 39298 22992 39304 23004
rect 39356 22992 39362 23044
rect 40310 22992 40316 23044
rect 40368 23032 40374 23044
rect 41248 23032 41276 23063
rect 43070 23060 43076 23072
rect 43128 23060 43134 23112
rect 45554 23060 45560 23112
rect 45612 23100 45618 23112
rect 45824 23103 45882 23109
rect 45612 23072 45657 23100
rect 45612 23060 45618 23072
rect 45824 23069 45836 23103
rect 45870 23100 45882 23103
rect 47026 23100 47032 23112
rect 45870 23072 47032 23100
rect 45870 23069 45882 23072
rect 45824 23063 45882 23069
rect 47026 23060 47032 23072
rect 47084 23060 47090 23112
rect 50157 23103 50215 23109
rect 50157 23069 50169 23103
rect 50203 23069 50215 23103
rect 50157 23063 50215 23069
rect 50424 23103 50482 23109
rect 50424 23069 50436 23103
rect 50470 23100 50482 23103
rect 51534 23100 51540 23112
rect 50470 23072 51540 23100
rect 50470 23069 50482 23072
rect 50424 23063 50482 23069
rect 40368 23004 41276 23032
rect 41500 23035 41558 23041
rect 40368 22992 40374 23004
rect 41500 23001 41512 23035
rect 41546 23032 41558 23035
rect 42426 23032 42432 23044
rect 41546 23004 42432 23032
rect 41546 23001 41558 23004
rect 41500 22995 41558 23001
rect 42426 22992 42432 23004
rect 42484 22992 42490 23044
rect 43340 23035 43398 23041
rect 43340 23001 43352 23035
rect 43386 23032 43398 23035
rect 44174 23032 44180 23044
rect 43386 23004 44180 23032
rect 43386 23001 43398 23004
rect 43340 22995 43398 23001
rect 44174 22992 44180 23004
rect 44232 22992 44238 23044
rect 48216 23035 48274 23041
rect 48216 23001 48228 23035
rect 48262 23032 48274 23035
rect 49602 23032 49608 23044
rect 48262 23004 49608 23032
rect 48262 23001 48274 23004
rect 48216 22995 48274 23001
rect 49602 22992 49608 23004
rect 49660 22992 49666 23044
rect 50172 23032 50200 23063
rect 51534 23060 51540 23072
rect 51592 23060 51598 23112
rect 51997 23103 52055 23109
rect 51997 23069 52009 23103
rect 52043 23100 52055 23103
rect 53374 23100 53380 23112
rect 52043 23072 53380 23100
rect 52043 23069 52055 23072
rect 51997 23063 52055 23069
rect 53374 23060 53380 23072
rect 53432 23060 53438 23112
rect 56778 23060 56784 23112
rect 56836 23100 56842 23112
rect 57149 23103 57207 23109
rect 57149 23100 57161 23103
rect 56836 23072 57161 23100
rect 56836 23060 56842 23072
rect 57149 23069 57161 23072
rect 57195 23069 57207 23103
rect 57149 23063 57207 23069
rect 50614 23032 50620 23044
rect 50172 23004 50620 23032
rect 50614 22992 50620 23004
rect 50672 22992 50678 23044
rect 52086 22992 52092 23044
rect 52144 23032 52150 23044
rect 52242 23035 52300 23041
rect 52242 23032 52254 23035
rect 52144 23004 52254 23032
rect 52144 22992 52150 23004
rect 52242 23001 52254 23004
rect 52288 23001 52300 23035
rect 52242 22995 52300 23001
rect 57416 23035 57474 23041
rect 57416 23001 57428 23035
rect 57462 23032 57474 23035
rect 58434 23032 58440 23044
rect 57462 23004 58440 23032
rect 57462 23001 57474 23004
rect 57416 22995 57474 23001
rect 58434 22992 58440 23004
rect 58492 22992 58498 23044
rect 3234 22964 3240 22976
rect 3195 22936 3240 22964
rect 3234 22924 3240 22936
rect 3292 22924 3298 22976
rect 10686 22964 10692 22976
rect 10647 22936 10692 22964
rect 10686 22924 10692 22936
rect 10744 22924 10750 22976
rect 20625 22967 20683 22973
rect 20625 22933 20637 22967
rect 20671 22964 20683 22967
rect 22094 22964 22100 22976
rect 20671 22936 22100 22964
rect 20671 22933 20683 22936
rect 20625 22927 20683 22933
rect 22094 22924 22100 22936
rect 22152 22924 22158 22976
rect 22462 22964 22468 22976
rect 22423 22936 22468 22964
rect 22462 22924 22468 22936
rect 22520 22924 22526 22976
rect 32306 22964 32312 22976
rect 32267 22936 32312 22964
rect 32306 22924 32312 22936
rect 32364 22924 32370 22976
rect 33502 22924 33508 22976
rect 33560 22964 33566 22976
rect 34149 22967 34207 22973
rect 34149 22964 34161 22967
rect 33560 22936 34161 22964
rect 33560 22924 33566 22936
rect 34149 22933 34161 22936
rect 34195 22933 34207 22967
rect 36630 22964 36636 22976
rect 36591 22936 36636 22964
rect 34149 22927 34207 22933
rect 36630 22924 36636 22936
rect 36688 22924 36694 22976
rect 37366 22924 37372 22976
rect 37424 22964 37430 22976
rect 39025 22967 39083 22973
rect 39025 22964 39037 22967
rect 37424 22936 39037 22964
rect 37424 22924 37430 22936
rect 39025 22933 39037 22936
rect 39071 22933 39083 22967
rect 39025 22927 39083 22933
rect 40126 22924 40132 22976
rect 40184 22964 40190 22976
rect 40405 22967 40463 22973
rect 40405 22964 40417 22967
rect 40184 22936 40417 22964
rect 40184 22924 40190 22936
rect 40405 22933 40417 22936
rect 40451 22964 40463 22967
rect 42058 22964 42064 22976
rect 40451 22936 42064 22964
rect 40451 22933 40463 22936
rect 40405 22927 40463 22933
rect 42058 22924 42064 22936
rect 42116 22924 42122 22976
rect 42610 22964 42616 22976
rect 42571 22936 42616 22964
rect 42610 22924 42616 22936
rect 42668 22924 42674 22976
rect 44450 22964 44456 22976
rect 44411 22936 44456 22964
rect 44450 22924 44456 22936
rect 44508 22924 44514 22976
rect 51534 22964 51540 22976
rect 51495 22936 51540 22964
rect 51534 22924 51540 22936
rect 51592 22924 51598 22976
rect 52730 22924 52736 22976
rect 52788 22964 52794 22976
rect 53377 22967 53435 22973
rect 53377 22964 53389 22967
rect 52788 22936 53389 22964
rect 52788 22924 52794 22936
rect 53377 22933 53389 22936
rect 53423 22933 53435 22967
rect 58526 22964 58532 22976
rect 58487 22936 58532 22964
rect 53377 22927 53435 22933
rect 58526 22924 58532 22936
rect 58584 22924 58590 22976
rect 1104 22874 59340 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 59340 22874
rect 1104 22800 59340 22822
rect 9306 22720 9312 22772
rect 9364 22760 9370 22772
rect 10597 22763 10655 22769
rect 10597 22760 10609 22763
rect 9364 22732 10609 22760
rect 9364 22720 9370 22732
rect 10597 22729 10609 22732
rect 10643 22729 10655 22763
rect 13078 22760 13084 22772
rect 13039 22732 13084 22760
rect 10597 22723 10655 22729
rect 13078 22720 13084 22732
rect 13136 22720 13142 22772
rect 21100 22732 22600 22760
rect 2492 22695 2550 22701
rect 2492 22661 2504 22695
rect 2538 22692 2550 22695
rect 3234 22692 3240 22704
rect 2538 22664 3240 22692
rect 2538 22661 2550 22664
rect 2492 22655 2550 22661
rect 3234 22652 3240 22664
rect 3292 22652 3298 22704
rect 9484 22695 9542 22701
rect 9484 22661 9496 22695
rect 9530 22692 9542 22695
rect 10686 22692 10692 22704
rect 9530 22664 10692 22692
rect 9530 22661 9542 22664
rect 9484 22655 9542 22661
rect 10686 22652 10692 22664
rect 10744 22652 10750 22704
rect 12250 22692 12256 22704
rect 11716 22664 12256 22692
rect 2222 22624 2228 22636
rect 2183 22596 2228 22624
rect 2222 22584 2228 22596
rect 2280 22584 2286 22636
rect 9214 22624 9220 22636
rect 9127 22596 9220 22624
rect 9214 22584 9220 22596
rect 9272 22624 9278 22636
rect 11716 22633 11744 22664
rect 12250 22652 12256 22664
rect 12308 22652 12314 22704
rect 15470 22692 15476 22704
rect 14752 22664 15476 22692
rect 11701 22627 11759 22633
rect 11701 22624 11713 22627
rect 9272 22596 11713 22624
rect 9272 22584 9278 22596
rect 11701 22593 11713 22596
rect 11747 22593 11759 22627
rect 11701 22587 11759 22593
rect 11968 22627 12026 22633
rect 11968 22593 11980 22627
rect 12014 22624 12026 22627
rect 12894 22624 12900 22636
rect 12014 22596 12900 22624
rect 12014 22593 12026 22596
rect 11968 22587 12026 22593
rect 12894 22584 12900 22596
rect 12952 22584 12958 22636
rect 14752 22633 14780 22664
rect 15470 22652 15476 22664
rect 15528 22652 15534 22704
rect 14737 22627 14795 22633
rect 14737 22593 14749 22627
rect 14783 22593 14795 22627
rect 14737 22587 14795 22593
rect 15004 22627 15062 22633
rect 15004 22593 15016 22627
rect 15050 22624 15062 22627
rect 15746 22624 15752 22636
rect 15050 22596 15752 22624
rect 15050 22593 15062 22596
rect 15004 22587 15062 22593
rect 15746 22584 15752 22596
rect 15804 22584 15810 22636
rect 18046 22584 18052 22636
rect 18104 22624 18110 22636
rect 18141 22627 18199 22633
rect 18141 22624 18153 22627
rect 18104 22596 18153 22624
rect 18104 22584 18110 22596
rect 18141 22593 18153 22596
rect 18187 22593 18199 22627
rect 18141 22587 18199 22593
rect 18408 22627 18466 22633
rect 18408 22593 18420 22627
rect 18454 22624 18466 22627
rect 20622 22624 20628 22636
rect 18454 22596 20628 22624
rect 18454 22593 18466 22596
rect 18408 22587 18466 22593
rect 20622 22584 20628 22596
rect 20680 22584 20686 22636
rect 20990 22584 20996 22636
rect 21048 22624 21054 22636
rect 21100 22633 21128 22732
rect 22088 22695 22146 22701
rect 22088 22661 22100 22695
rect 22134 22692 22146 22695
rect 22462 22692 22468 22704
rect 22134 22664 22468 22692
rect 22134 22661 22146 22664
rect 22088 22655 22146 22661
rect 22462 22652 22468 22664
rect 22520 22652 22526 22704
rect 22572 22692 22600 22732
rect 23106 22720 23112 22772
rect 23164 22760 23170 22772
rect 23201 22763 23259 22769
rect 23201 22760 23213 22763
rect 23164 22732 23213 22760
rect 23164 22720 23170 22732
rect 23201 22729 23213 22732
rect 23247 22729 23259 22763
rect 25130 22760 25136 22772
rect 23201 22723 23259 22729
rect 23676 22732 24256 22760
rect 25091 22732 25136 22760
rect 23676 22692 23704 22732
rect 24118 22692 24124 22704
rect 22572 22664 23704 22692
rect 23768 22664 24124 22692
rect 21085 22627 21143 22633
rect 21085 22624 21097 22627
rect 21048 22596 21097 22624
rect 21048 22584 21054 22596
rect 21085 22593 21097 22596
rect 21131 22593 21143 22627
rect 21085 22587 21143 22593
rect 21726 22584 21732 22636
rect 21784 22624 21790 22636
rect 23768 22633 23796 22664
rect 24118 22652 24124 22664
rect 24176 22652 24182 22704
rect 24228 22692 24256 22732
rect 25130 22720 25136 22732
rect 25188 22720 25194 22772
rect 30926 22760 30932 22772
rect 26206 22732 30328 22760
rect 30887 22732 30932 22760
rect 26206 22692 26234 22732
rect 24228 22664 26234 22692
rect 27341 22695 27399 22701
rect 27341 22661 27353 22695
rect 27387 22692 27399 22695
rect 27798 22692 27804 22704
rect 27387 22664 27804 22692
rect 27387 22661 27399 22664
rect 27341 22655 27399 22661
rect 21821 22627 21879 22633
rect 21821 22624 21833 22627
rect 21784 22596 21833 22624
rect 21784 22584 21790 22596
rect 21821 22593 21833 22596
rect 21867 22593 21879 22627
rect 21821 22587 21879 22593
rect 23753 22627 23811 22633
rect 23753 22593 23765 22627
rect 23799 22593 23811 22627
rect 23753 22587 23811 22593
rect 24020 22627 24078 22633
rect 24020 22593 24032 22627
rect 24066 22624 24078 22627
rect 25774 22624 25780 22636
rect 24066 22596 25780 22624
rect 24066 22593 24078 22596
rect 24020 22587 24078 22593
rect 25774 22584 25780 22596
rect 25832 22584 25838 22636
rect 25958 22516 25964 22568
rect 26016 22556 26022 22568
rect 27356 22556 27384 22655
rect 27798 22652 27804 22664
rect 27856 22652 27862 22704
rect 29816 22695 29874 22701
rect 29816 22661 29828 22695
rect 29862 22692 29874 22695
rect 30190 22692 30196 22704
rect 29862 22664 30196 22692
rect 29862 22661 29874 22664
rect 29816 22655 29874 22661
rect 30190 22652 30196 22664
rect 30248 22652 30254 22704
rect 30300 22692 30328 22732
rect 30926 22720 30932 22732
rect 30984 22720 30990 22772
rect 44818 22720 44824 22772
rect 44876 22760 44882 22772
rect 46201 22763 46259 22769
rect 46201 22760 46213 22763
rect 44876 22732 46213 22760
rect 44876 22720 44882 22732
rect 46201 22729 46213 22732
rect 46247 22729 46259 22763
rect 49602 22760 49608 22772
rect 49563 22732 49608 22760
rect 46201 22723 46259 22729
rect 49602 22720 49608 22732
rect 49660 22720 49666 22772
rect 50614 22760 50620 22772
rect 49712 22732 50620 22760
rect 31110 22692 31116 22704
rect 30300 22664 31116 22692
rect 31110 22652 31116 22664
rect 31168 22652 31174 22704
rect 43248 22695 43306 22701
rect 38488 22664 40356 22692
rect 32766 22584 32772 22636
rect 32824 22624 32830 22636
rect 33505 22627 33563 22633
rect 33505 22624 33517 22627
rect 32824 22596 33517 22624
rect 32824 22584 32830 22596
rect 33505 22593 33517 22596
rect 33551 22593 33563 22627
rect 33505 22587 33563 22593
rect 33772 22627 33830 22633
rect 33772 22593 33784 22627
rect 33818 22624 33830 22627
rect 34146 22624 34152 22636
rect 33818 22596 34152 22624
rect 33818 22593 33830 22596
rect 33772 22587 33830 22593
rect 34146 22584 34152 22596
rect 34204 22584 34210 22636
rect 35342 22624 35348 22636
rect 35303 22596 35348 22624
rect 35342 22584 35348 22596
rect 35400 22584 35406 22636
rect 35612 22627 35670 22633
rect 35612 22593 35624 22627
rect 35658 22624 35670 22627
rect 37458 22624 37464 22636
rect 35658 22596 37464 22624
rect 35658 22593 35670 22596
rect 35612 22587 35670 22593
rect 37458 22584 37464 22596
rect 37516 22584 37522 22636
rect 29549 22559 29607 22565
rect 29549 22556 29561 22559
rect 26016 22528 27384 22556
rect 28644 22528 29561 22556
rect 26016 22516 26022 22528
rect 3602 22420 3608 22432
rect 3563 22392 3608 22420
rect 3602 22380 3608 22392
rect 3660 22380 3666 22432
rect 16114 22420 16120 22432
rect 16075 22392 16120 22420
rect 16114 22380 16120 22392
rect 16172 22380 16178 22432
rect 19521 22423 19579 22429
rect 19521 22389 19533 22423
rect 19567 22420 19579 22423
rect 20806 22420 20812 22432
rect 19567 22392 20812 22420
rect 19567 22389 19579 22392
rect 19521 22383 19579 22389
rect 20806 22380 20812 22392
rect 20864 22380 20870 22432
rect 20898 22380 20904 22432
rect 20956 22420 20962 22432
rect 20956 22392 21001 22420
rect 20956 22380 20962 22392
rect 27614 22380 27620 22432
rect 27672 22420 27678 22432
rect 28644 22429 28672 22528
rect 29549 22525 29561 22528
rect 29595 22525 29607 22559
rect 29549 22519 29607 22525
rect 37642 22516 37648 22568
rect 37700 22556 37706 22568
rect 38488 22565 38516 22664
rect 40328 22636 40356 22664
rect 43248 22661 43260 22695
rect 43294 22692 43306 22695
rect 45186 22692 45192 22704
rect 43294 22664 45192 22692
rect 43294 22661 43306 22664
rect 43248 22655 43306 22661
rect 45186 22652 45192 22664
rect 45244 22652 45250 22704
rect 49712 22692 49740 22732
rect 50614 22720 50620 22732
rect 50672 22720 50678 22772
rect 57238 22760 57244 22772
rect 57199 22732 57244 22760
rect 57238 22720 57244 22732
rect 57296 22720 57302 22772
rect 48240 22664 49740 22692
rect 50424 22695 50482 22701
rect 38740 22627 38798 22633
rect 38740 22593 38752 22627
rect 38786 22624 38798 22627
rect 40218 22624 40224 22636
rect 38786 22596 40224 22624
rect 38786 22593 38798 22596
rect 38740 22587 38798 22593
rect 40218 22584 40224 22596
rect 40276 22584 40282 22636
rect 40310 22584 40316 22636
rect 40368 22624 40374 22636
rect 40580 22627 40638 22633
rect 40368 22596 40461 22624
rect 40368 22584 40374 22596
rect 40580 22593 40592 22627
rect 40626 22624 40638 22627
rect 41874 22624 41880 22636
rect 40626 22596 41880 22624
rect 40626 22593 40638 22596
rect 40580 22587 40638 22593
rect 41874 22584 41880 22596
rect 41932 22584 41938 22636
rect 42981 22627 43039 22633
rect 42981 22593 42993 22627
rect 43027 22624 43039 22627
rect 43070 22624 43076 22636
rect 43027 22596 43076 22624
rect 43027 22593 43039 22596
rect 42981 22587 43039 22593
rect 43070 22584 43076 22596
rect 43128 22624 43134 22636
rect 45088 22627 45146 22633
rect 43128 22596 44864 22624
rect 43128 22584 43134 22596
rect 44836 22565 44864 22596
rect 45088 22593 45100 22627
rect 45134 22624 45146 22627
rect 46382 22624 46388 22636
rect 45134 22596 46388 22624
rect 45134 22593 45146 22596
rect 45088 22587 45146 22593
rect 46382 22584 46388 22596
rect 46440 22584 46446 22636
rect 48240 22633 48268 22664
rect 50424 22661 50436 22695
rect 50470 22692 50482 22695
rect 51534 22692 51540 22704
rect 50470 22664 51540 22692
rect 50470 22661 50482 22664
rect 50424 22655 50482 22661
rect 51534 22652 51540 22664
rect 51592 22652 51598 22704
rect 56128 22695 56186 22701
rect 56128 22661 56140 22695
rect 56174 22692 56186 22695
rect 58526 22692 58532 22704
rect 56174 22664 58532 22692
rect 56174 22661 56186 22664
rect 56128 22655 56186 22661
rect 58526 22652 58532 22664
rect 58584 22652 58590 22704
rect 48225 22627 48283 22633
rect 48225 22593 48237 22627
rect 48271 22593 48283 22627
rect 48225 22587 48283 22593
rect 48492 22627 48550 22633
rect 48492 22593 48504 22627
rect 48538 22624 48550 22627
rect 49694 22624 49700 22636
rect 48538 22596 49700 22624
rect 48538 22593 48550 22596
rect 48492 22587 48550 22593
rect 49694 22584 49700 22596
rect 49752 22584 49758 22636
rect 50154 22624 50160 22636
rect 50115 22596 50160 22624
rect 50154 22584 50160 22596
rect 50212 22584 50218 22636
rect 53000 22627 53058 22633
rect 53000 22593 53012 22627
rect 53046 22624 53058 22627
rect 55950 22624 55956 22636
rect 53046 22596 55956 22624
rect 53046 22593 53058 22596
rect 53000 22587 53058 22593
rect 55950 22584 55956 22596
rect 56008 22584 56014 22636
rect 38473 22559 38531 22565
rect 38473 22556 38485 22559
rect 37700 22528 38485 22556
rect 37700 22516 37706 22528
rect 38473 22525 38485 22528
rect 38519 22525 38531 22559
rect 38473 22519 38531 22525
rect 44821 22559 44879 22565
rect 44821 22525 44833 22559
rect 44867 22525 44879 22559
rect 44821 22519 44879 22525
rect 28629 22423 28687 22429
rect 28629 22420 28641 22423
rect 27672 22392 28641 22420
rect 27672 22380 27678 22392
rect 28629 22389 28641 22392
rect 28675 22389 28687 22423
rect 28629 22383 28687 22389
rect 34514 22380 34520 22432
rect 34572 22420 34578 22432
rect 34885 22423 34943 22429
rect 34885 22420 34897 22423
rect 34572 22392 34897 22420
rect 34572 22380 34578 22392
rect 34885 22389 34897 22392
rect 34931 22389 34943 22423
rect 36722 22420 36728 22432
rect 36683 22392 36728 22420
rect 34885 22383 34943 22389
rect 36722 22380 36728 22392
rect 36780 22380 36786 22432
rect 39850 22420 39856 22432
rect 39811 22392 39856 22420
rect 39850 22380 39856 22392
rect 39908 22380 39914 22432
rect 41690 22420 41696 22432
rect 41651 22392 41696 22420
rect 41690 22380 41696 22392
rect 41748 22380 41754 22432
rect 42058 22380 42064 22432
rect 42116 22420 42122 22432
rect 42794 22420 42800 22432
rect 42116 22392 42800 22420
rect 42116 22380 42122 22392
rect 42794 22380 42800 22392
rect 42852 22380 42858 22432
rect 44358 22420 44364 22432
rect 44319 22392 44364 22420
rect 44358 22380 44364 22392
rect 44416 22380 44422 22432
rect 44836 22420 44864 22519
rect 51994 22516 52000 22568
rect 52052 22556 52058 22568
rect 52733 22559 52791 22565
rect 52733 22556 52745 22559
rect 52052 22528 52745 22556
rect 52052 22516 52058 22528
rect 52733 22525 52745 22528
rect 52779 22525 52791 22559
rect 52733 22519 52791 22525
rect 55861 22559 55919 22565
rect 55861 22525 55873 22559
rect 55907 22525 55919 22559
rect 55861 22519 55919 22525
rect 55122 22448 55128 22500
rect 55180 22488 55186 22500
rect 55876 22488 55904 22519
rect 55180 22460 55904 22488
rect 55180 22448 55186 22460
rect 45554 22420 45560 22432
rect 44836 22392 45560 22420
rect 45554 22380 45560 22392
rect 45612 22380 45618 22432
rect 51166 22380 51172 22432
rect 51224 22420 51230 22432
rect 51537 22423 51595 22429
rect 51537 22420 51549 22423
rect 51224 22392 51549 22420
rect 51224 22380 51230 22392
rect 51537 22389 51549 22392
rect 51583 22389 51595 22423
rect 51537 22383 51595 22389
rect 54113 22423 54171 22429
rect 54113 22389 54125 22423
rect 54159 22420 54171 22423
rect 55398 22420 55404 22432
rect 54159 22392 55404 22420
rect 54159 22389 54171 22392
rect 54113 22383 54171 22389
rect 55398 22380 55404 22392
rect 55456 22380 55462 22432
rect 55876 22420 55904 22460
rect 56778 22420 56784 22432
rect 55876 22392 56784 22420
rect 56778 22380 56784 22392
rect 56836 22380 56842 22432
rect 1104 22330 59340 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 59340 22330
rect 1104 22256 59340 22278
rect 20622 22216 20628 22228
rect 20583 22188 20628 22216
rect 20622 22176 20628 22188
rect 20680 22176 20686 22228
rect 25774 22216 25780 22228
rect 25735 22188 25780 22216
rect 25774 22176 25780 22188
rect 25832 22176 25838 22228
rect 31846 22176 31852 22228
rect 31904 22216 31910 22228
rect 32309 22219 32367 22225
rect 32309 22216 32321 22219
rect 31904 22188 32321 22216
rect 31904 22176 31910 22188
rect 32309 22185 32321 22188
rect 32355 22185 32367 22219
rect 34146 22216 34152 22228
rect 34107 22188 34152 22216
rect 32309 22179 32367 22185
rect 34146 22176 34152 22188
rect 34204 22176 34210 22228
rect 37458 22216 37464 22228
rect 37419 22188 37464 22216
rect 37458 22176 37464 22188
rect 37516 22176 37522 22228
rect 39298 22216 39304 22228
rect 39259 22188 39304 22216
rect 39298 22176 39304 22188
rect 39356 22176 39362 22228
rect 42426 22176 42432 22228
rect 42484 22216 42490 22228
rect 42613 22219 42671 22225
rect 42613 22216 42625 22219
rect 42484 22188 42625 22216
rect 42484 22176 42490 22188
rect 42613 22185 42625 22188
rect 42659 22185 42671 22219
rect 42613 22179 42671 22185
rect 44174 22176 44180 22228
rect 44232 22216 44238 22228
rect 44453 22219 44511 22225
rect 44453 22216 44465 22219
rect 44232 22188 44465 22216
rect 44232 22176 44238 22188
rect 44453 22185 44465 22188
rect 44499 22185 44511 22219
rect 44453 22179 44511 22185
rect 51997 22219 52055 22225
rect 51997 22185 52009 22219
rect 52043 22216 52055 22219
rect 52086 22216 52092 22228
rect 52043 22188 52092 22216
rect 52043 22185 52055 22188
rect 51997 22179 52055 22185
rect 52086 22176 52092 22188
rect 52144 22176 52150 22228
rect 15470 22040 15476 22092
rect 15528 22080 15534 22092
rect 15749 22083 15807 22089
rect 15749 22080 15761 22083
rect 15528 22052 15761 22080
rect 15528 22040 15534 22052
rect 15749 22049 15761 22052
rect 15795 22049 15807 22083
rect 15749 22043 15807 22049
rect 1857 22015 1915 22021
rect 1857 21981 1869 22015
rect 1903 21981 1915 22015
rect 1857 21975 1915 21981
rect 2124 22015 2182 22021
rect 2124 21981 2136 22015
rect 2170 22012 2182 22015
rect 3602 22012 3608 22024
rect 2170 21984 3608 22012
rect 2170 21981 2182 21984
rect 2124 21975 2182 21981
rect 1872 21944 1900 21975
rect 3602 21972 3608 21984
rect 3660 21972 3666 22024
rect 3789 22015 3847 22021
rect 3789 21981 3801 22015
rect 3835 22012 3847 22015
rect 4430 22012 4436 22024
rect 3835 21984 4436 22012
rect 3835 21981 3847 21984
rect 3789 21975 3847 21981
rect 4430 21972 4436 21984
rect 4488 22012 4494 22024
rect 5166 22012 5172 22024
rect 4488 21984 5172 22012
rect 4488 21972 4494 21984
rect 5166 21972 5172 21984
rect 5224 22012 5230 22024
rect 5442 22012 5448 22024
rect 5224 21984 5448 22012
rect 5224 21972 5230 21984
rect 5442 21972 5448 21984
rect 5500 21972 5506 22024
rect 11609 22015 11667 22021
rect 11609 21981 11621 22015
rect 11655 22012 11667 22015
rect 12250 22012 12256 22024
rect 11655 21984 12256 22012
rect 11655 21981 11667 21984
rect 11609 21975 11667 21981
rect 12250 21972 12256 21984
rect 12308 21972 12314 22024
rect 15764 22012 15792 22043
rect 30834 22040 30840 22092
rect 30892 22080 30898 22092
rect 30929 22083 30987 22089
rect 30929 22080 30941 22083
rect 30892 22052 30941 22080
rect 30892 22040 30898 22052
rect 30929 22049 30941 22052
rect 30975 22049 30987 22083
rect 30929 22043 30987 22049
rect 15838 22012 15844 22024
rect 15764 21984 15844 22012
rect 15838 21972 15844 21984
rect 15896 21972 15902 22024
rect 16022 22021 16028 22024
rect 16016 22012 16028 22021
rect 15983 21984 16028 22012
rect 16016 21975 16028 21984
rect 16022 21972 16028 21975
rect 16080 21972 16086 22024
rect 19150 21972 19156 22024
rect 19208 22012 19214 22024
rect 19245 22015 19303 22021
rect 19245 22012 19257 22015
rect 19208 21984 19257 22012
rect 19208 21972 19214 21984
rect 19245 21981 19257 21984
rect 19291 21981 19303 22015
rect 21082 22012 21088 22024
rect 21043 21984 21088 22012
rect 19245 21975 19303 21981
rect 21082 21972 21088 21984
rect 21140 21972 21146 22024
rect 21726 21972 21732 22024
rect 21784 22012 21790 22024
rect 24397 22015 24455 22021
rect 24397 22012 24409 22015
rect 21784 21984 24409 22012
rect 21784 21972 21790 21984
rect 24397 21981 24409 21984
rect 24443 21981 24455 22015
rect 27614 22012 27620 22024
rect 27575 21984 27620 22012
rect 24397 21975 24455 21981
rect 27614 21972 27620 21984
rect 27672 21972 27678 22024
rect 30944 22012 30972 22043
rect 37642 22040 37648 22092
rect 37700 22080 37706 22092
rect 37921 22083 37979 22089
rect 37921 22080 37933 22083
rect 37700 22052 37933 22080
rect 37700 22040 37706 22052
rect 37921 22049 37933 22052
rect 37967 22049 37979 22083
rect 37921 22043 37979 22049
rect 32769 22015 32827 22021
rect 32769 22012 32781 22015
rect 30944 21984 32781 22012
rect 32769 21981 32781 21984
rect 32815 21981 32827 22015
rect 36078 22012 36084 22024
rect 36039 21984 36084 22012
rect 32769 21975 32827 21981
rect 36078 21972 36084 21984
rect 36136 21972 36142 22024
rect 36348 22015 36406 22021
rect 36348 21981 36360 22015
rect 36394 22012 36406 22015
rect 37366 22012 37372 22024
rect 36394 21984 37372 22012
rect 36394 21981 36406 21984
rect 36348 21975 36406 21981
rect 37366 21972 37372 21984
rect 37424 21972 37430 22024
rect 38194 22021 38200 22024
rect 38188 22012 38200 22021
rect 38155 21984 38200 22012
rect 38188 21975 38200 21984
rect 38194 21972 38200 21975
rect 38252 21972 38258 22024
rect 40310 21972 40316 22024
rect 40368 22012 40374 22024
rect 41233 22015 41291 22021
rect 41233 22012 41245 22015
rect 40368 21984 41245 22012
rect 40368 21972 40374 21984
rect 41233 21981 41245 21984
rect 41279 22012 41291 22015
rect 43073 22015 43131 22021
rect 43073 22012 43085 22015
rect 41279 21984 43085 22012
rect 41279 21981 41291 21984
rect 41233 21975 41291 21981
rect 43073 21981 43085 21984
rect 43119 21981 43131 22015
rect 43073 21975 43131 21981
rect 43340 22015 43398 22021
rect 43340 21981 43352 22015
rect 43386 22012 43398 22015
rect 44358 22012 44364 22024
rect 43386 21984 44364 22012
rect 43386 21981 43398 21984
rect 43340 21975 43398 21981
rect 44358 21972 44364 21984
rect 44416 21972 44422 22024
rect 46293 22015 46351 22021
rect 46293 21981 46305 22015
rect 46339 22012 46351 22015
rect 49970 22012 49976 22024
rect 46339 21984 49976 22012
rect 46339 21981 46351 21984
rect 46293 21975 46351 21981
rect 49970 21972 49976 21984
rect 50028 21972 50034 22024
rect 50614 22012 50620 22024
rect 50527 21984 50620 22012
rect 50614 21972 50620 21984
rect 50672 21972 50678 22024
rect 50884 22015 50942 22021
rect 50884 21981 50896 22015
rect 50930 22012 50942 22015
rect 51166 22012 51172 22024
rect 50930 21984 51172 22012
rect 50930 21981 50942 21984
rect 50884 21975 50942 21981
rect 51166 21972 51172 21984
rect 51224 21972 51230 22024
rect 52730 22021 52736 22024
rect 52457 22015 52515 22021
rect 52457 21981 52469 22015
rect 52503 21981 52515 22015
rect 52724 22012 52736 22021
rect 52691 21984 52736 22012
rect 52457 21975 52515 21981
rect 52724 21975 52736 21984
rect 2222 21944 2228 21956
rect 1872 21916 2228 21944
rect 2222 21904 2228 21916
rect 2280 21904 2286 21956
rect 3418 21904 3424 21956
rect 3476 21944 3482 21956
rect 4034 21947 4092 21953
rect 4034 21944 4046 21947
rect 3476 21916 4046 21944
rect 3476 21904 3482 21916
rect 4034 21913 4046 21916
rect 4080 21913 4092 21947
rect 4034 21907 4092 21913
rect 11876 21947 11934 21953
rect 11876 21913 11888 21947
rect 11922 21944 11934 21947
rect 13262 21944 13268 21956
rect 11922 21916 13268 21944
rect 11922 21913 11934 21916
rect 11876 21907 11934 21913
rect 13262 21904 13268 21916
rect 13320 21904 13326 21956
rect 19512 21947 19570 21953
rect 19512 21913 19524 21947
rect 19558 21944 19570 21947
rect 20530 21944 20536 21956
rect 19558 21916 20536 21944
rect 19558 21913 19570 21916
rect 19512 21907 19570 21913
rect 20530 21904 20536 21916
rect 20588 21904 20594 21956
rect 21352 21947 21410 21953
rect 21352 21913 21364 21947
rect 21398 21944 21410 21947
rect 23198 21944 23204 21956
rect 21398 21916 23204 21944
rect 21398 21913 21410 21916
rect 21352 21907 21410 21913
rect 23198 21904 23204 21916
rect 23256 21904 23262 21956
rect 24664 21947 24722 21953
rect 24664 21913 24676 21947
rect 24710 21944 24722 21947
rect 25130 21944 25136 21956
rect 24710 21916 25136 21944
rect 24710 21913 24722 21916
rect 24664 21907 24722 21913
rect 25130 21904 25136 21916
rect 25188 21904 25194 21956
rect 27884 21947 27942 21953
rect 27884 21913 27896 21947
rect 27930 21944 27942 21947
rect 28902 21944 28908 21956
rect 27930 21916 28908 21944
rect 27930 21913 27942 21916
rect 27884 21907 27942 21913
rect 28902 21904 28908 21916
rect 28960 21904 28966 21956
rect 31196 21947 31254 21953
rect 31196 21913 31208 21947
rect 31242 21944 31254 21947
rect 33036 21947 33094 21953
rect 31242 21916 32996 21944
rect 31242 21913 31254 21916
rect 31196 21907 31254 21913
rect 3234 21876 3240 21888
rect 3195 21848 3240 21876
rect 3234 21836 3240 21848
rect 3292 21836 3298 21888
rect 5166 21876 5172 21888
rect 5127 21848 5172 21876
rect 5166 21836 5172 21848
rect 5224 21836 5230 21888
rect 12986 21876 12992 21888
rect 12947 21848 12992 21876
rect 12986 21836 12992 21848
rect 13044 21836 13050 21888
rect 15746 21836 15752 21888
rect 15804 21876 15810 21888
rect 17129 21879 17187 21885
rect 17129 21876 17141 21879
rect 15804 21848 17141 21876
rect 15804 21836 15810 21848
rect 17129 21845 17141 21848
rect 17175 21845 17187 21879
rect 17129 21839 17187 21845
rect 21174 21836 21180 21888
rect 21232 21876 21238 21888
rect 22465 21879 22523 21885
rect 22465 21876 22477 21879
rect 21232 21848 22477 21876
rect 21232 21836 21238 21848
rect 22465 21845 22477 21848
rect 22511 21845 22523 21879
rect 28994 21876 29000 21888
rect 28955 21848 29000 21876
rect 22465 21839 22523 21845
rect 28994 21836 29000 21848
rect 29052 21836 29058 21888
rect 32968 21876 32996 21916
rect 33036 21913 33048 21947
rect 33082 21944 33094 21947
rect 36262 21944 36268 21956
rect 33082 21916 36268 21944
rect 33082 21913 33094 21916
rect 33036 21907 33094 21913
rect 36262 21904 36268 21916
rect 36320 21904 36326 21956
rect 41500 21947 41558 21953
rect 41500 21913 41512 21947
rect 41546 21944 41558 21947
rect 44082 21944 44088 21956
rect 41546 21916 44088 21944
rect 41546 21913 41558 21916
rect 41500 21907 41558 21913
rect 44082 21904 44088 21916
rect 44140 21904 44146 21956
rect 50632 21944 50660 21972
rect 50982 21944 50988 21956
rect 50632 21916 50988 21944
rect 50982 21904 50988 21916
rect 51040 21944 51046 21956
rect 52472 21944 52500 21975
rect 52730 21972 52736 21975
rect 52788 21972 52794 22024
rect 55674 21972 55680 22024
rect 55732 22012 55738 22024
rect 56137 22015 56195 22021
rect 56137 22012 56149 22015
rect 55732 21984 56149 22012
rect 55732 21972 55738 21984
rect 56137 21981 56149 21984
rect 56183 22012 56195 22015
rect 56410 22012 56416 22024
rect 56183 21984 56416 22012
rect 56183 21981 56195 21984
rect 56137 21975 56195 21981
rect 56410 21972 56416 21984
rect 56468 21972 56474 22024
rect 51040 21916 52500 21944
rect 51040 21904 51046 21916
rect 33870 21876 33876 21888
rect 32968 21848 33876 21876
rect 33870 21836 33876 21848
rect 33928 21836 33934 21888
rect 47578 21876 47584 21888
rect 47539 21848 47584 21876
rect 47578 21836 47584 21848
rect 47636 21836 47642 21888
rect 53834 21876 53840 21888
rect 53795 21848 53840 21876
rect 53834 21836 53840 21848
rect 53892 21836 53898 21888
rect 56778 21836 56784 21888
rect 56836 21876 56842 21888
rect 57425 21879 57483 21885
rect 57425 21876 57437 21879
rect 56836 21848 57437 21876
rect 56836 21836 56842 21848
rect 57425 21845 57437 21848
rect 57471 21845 57483 21879
rect 57425 21839 57483 21845
rect 1104 21786 59340 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 59340 21786
rect 1104 21712 59340 21734
rect 3418 21672 3424 21684
rect 3379 21644 3424 21672
rect 3418 21632 3424 21644
rect 3476 21632 3482 21684
rect 16117 21675 16175 21681
rect 16117 21641 16129 21675
rect 16163 21672 16175 21675
rect 16163 21644 16574 21672
rect 16163 21641 16175 21644
rect 16117 21635 16175 21641
rect 2308 21607 2366 21613
rect 2308 21573 2320 21607
rect 2354 21604 2366 21607
rect 3234 21604 3240 21616
rect 2354 21576 3240 21604
rect 2354 21573 2366 21576
rect 2308 21567 2366 21573
rect 3234 21564 3240 21576
rect 3292 21564 3298 21616
rect 4148 21607 4206 21613
rect 4148 21573 4160 21607
rect 4194 21604 4206 21607
rect 5166 21604 5172 21616
rect 4194 21576 5172 21604
rect 4194 21573 4206 21576
rect 4148 21567 4206 21573
rect 5166 21564 5172 21576
rect 5224 21564 5230 21616
rect 16546 21604 16574 21644
rect 22830 21632 22836 21684
rect 22888 21672 22894 21684
rect 23201 21675 23259 21681
rect 23201 21672 23213 21675
rect 22888 21644 23213 21672
rect 22888 21632 22894 21644
rect 23201 21641 23213 21644
rect 23247 21641 23259 21675
rect 25130 21672 25136 21684
rect 25091 21644 25136 21672
rect 23201 21635 23259 21641
rect 25130 21632 25136 21644
rect 25188 21632 25194 21684
rect 28902 21632 28908 21684
rect 28960 21672 28966 21684
rect 28997 21675 29055 21681
rect 28997 21672 29009 21675
rect 28960 21644 29009 21672
rect 28960 21632 28966 21644
rect 28997 21641 29009 21644
rect 29043 21641 29055 21675
rect 28997 21635 29055 21641
rect 34790 21632 34796 21684
rect 34848 21672 34854 21684
rect 34885 21675 34943 21681
rect 34885 21672 34897 21675
rect 34848 21644 34897 21672
rect 34848 21632 34854 21644
rect 34885 21641 34897 21644
rect 34931 21641 34943 21675
rect 34885 21635 34943 21641
rect 36538 21632 36544 21684
rect 36596 21672 36602 21684
rect 36725 21675 36783 21681
rect 36725 21672 36737 21675
rect 36596 21644 36737 21672
rect 36596 21632 36602 21644
rect 36725 21641 36737 21644
rect 36771 21641 36783 21675
rect 40034 21672 40040 21684
rect 39995 21644 40040 21672
rect 36725 21635 36783 21641
rect 40034 21632 40040 21644
rect 40092 21632 40098 21684
rect 41874 21672 41880 21684
rect 41835 21644 41880 21672
rect 41874 21632 41880 21644
rect 41932 21632 41938 21684
rect 49694 21672 49700 21684
rect 49655 21644 49700 21672
rect 49694 21632 49700 21644
rect 49752 21632 49758 21684
rect 51537 21675 51595 21681
rect 51537 21641 51549 21675
rect 51583 21641 51595 21675
rect 51537 21635 51595 21641
rect 22094 21613 22100 21616
rect 16914 21607 16972 21613
rect 16914 21604 16926 21607
rect 16546 21576 16926 21604
rect 16914 21573 16926 21576
rect 16960 21573 16972 21607
rect 22088 21604 22100 21613
rect 22055 21576 22100 21604
rect 16914 21567 16972 21573
rect 22088 21567 22100 21576
rect 22094 21564 22100 21567
rect 22152 21564 22158 21616
rect 30460 21607 30518 21613
rect 30460 21573 30472 21607
rect 30506 21604 30518 21607
rect 32306 21604 32312 21616
rect 30506 21576 32312 21604
rect 30506 21573 30518 21576
rect 30460 21567 30518 21573
rect 32306 21564 32312 21576
rect 32364 21564 32370 21616
rect 33772 21607 33830 21613
rect 33772 21573 33784 21607
rect 33818 21604 33830 21607
rect 34514 21604 34520 21616
rect 33818 21576 34520 21604
rect 33818 21573 33830 21576
rect 33772 21567 33830 21573
rect 34514 21564 34520 21576
rect 34572 21564 34578 21616
rect 36078 21604 36084 21616
rect 35360 21576 36084 21604
rect 2041 21539 2099 21545
rect 2041 21505 2053 21539
rect 2087 21536 2099 21539
rect 2130 21536 2136 21548
rect 2087 21508 2136 21536
rect 2087 21505 2099 21508
rect 2041 21499 2099 21505
rect 2130 21496 2136 21508
rect 2188 21496 2194 21548
rect 3881 21539 3939 21545
rect 3881 21505 3893 21539
rect 3927 21536 3939 21539
rect 4430 21536 4436 21548
rect 3927 21508 4436 21536
rect 3927 21505 3939 21508
rect 3881 21499 3939 21505
rect 4430 21496 4436 21508
rect 4488 21496 4494 21548
rect 7276 21539 7334 21545
rect 7276 21505 7288 21539
rect 7322 21536 7334 21539
rect 9582 21536 9588 21548
rect 7322 21508 9588 21536
rect 7322 21505 7334 21508
rect 7276 21499 7334 21505
rect 9582 21496 9588 21508
rect 9640 21496 9646 21548
rect 12250 21536 12256 21548
rect 12211 21508 12256 21536
rect 12250 21496 12256 21508
rect 12308 21496 12314 21548
rect 12520 21539 12578 21545
rect 12520 21505 12532 21539
rect 12566 21536 12578 21539
rect 14458 21536 14464 21548
rect 12566 21508 14464 21536
rect 12566 21505 12578 21508
rect 12520 21499 12578 21505
rect 14458 21496 14464 21508
rect 14516 21496 14522 21548
rect 14734 21536 14740 21548
rect 14695 21508 14740 21536
rect 14734 21496 14740 21508
rect 14792 21496 14798 21548
rect 15004 21539 15062 21545
rect 15004 21505 15016 21539
rect 15050 21536 15062 21539
rect 16482 21536 16488 21548
rect 15050 21508 16488 21536
rect 15050 21505 15062 21508
rect 15004 21499 15062 21505
rect 16482 21496 16488 21508
rect 16540 21496 16546 21548
rect 18046 21496 18052 21548
rect 18104 21536 18110 21548
rect 18414 21536 18420 21548
rect 18104 21508 18420 21536
rect 18104 21496 18110 21508
rect 18414 21496 18420 21508
rect 18472 21536 18478 21548
rect 18509 21539 18567 21545
rect 18509 21536 18521 21539
rect 18472 21508 18521 21536
rect 18472 21496 18478 21508
rect 18509 21505 18521 21508
rect 18555 21505 18567 21539
rect 18509 21499 18567 21505
rect 18776 21539 18834 21545
rect 18776 21505 18788 21539
rect 18822 21536 18834 21539
rect 20622 21536 20628 21548
rect 18822 21508 20628 21536
rect 18822 21505 18834 21508
rect 18776 21499 18834 21505
rect 20622 21496 20628 21508
rect 20680 21496 20686 21548
rect 21726 21496 21732 21548
rect 21784 21536 21790 21548
rect 21821 21539 21879 21545
rect 21821 21536 21833 21539
rect 21784 21508 21833 21536
rect 21784 21496 21790 21508
rect 21821 21505 21833 21508
rect 21867 21505 21879 21539
rect 21821 21499 21879 21505
rect 24020 21539 24078 21545
rect 24020 21505 24032 21539
rect 24066 21536 24078 21539
rect 25774 21536 25780 21548
rect 24066 21508 25780 21536
rect 24066 21505 24078 21508
rect 24020 21499 24078 21505
rect 25774 21496 25780 21508
rect 25832 21496 25838 21548
rect 27884 21539 27942 21545
rect 27884 21505 27896 21539
rect 27930 21536 27942 21539
rect 28810 21536 28816 21548
rect 27930 21508 28816 21536
rect 27930 21505 27942 21508
rect 27884 21499 27942 21505
rect 28810 21496 28816 21508
rect 28868 21496 28874 21548
rect 30006 21496 30012 21548
rect 30064 21536 30070 21548
rect 30193 21539 30251 21545
rect 30193 21536 30205 21539
rect 30064 21508 30205 21536
rect 30064 21496 30070 21508
rect 30193 21505 30205 21508
rect 30239 21536 30251 21539
rect 30834 21536 30840 21548
rect 30239 21508 30840 21536
rect 30239 21505 30251 21508
rect 30193 21499 30251 21505
rect 30834 21496 30840 21508
rect 30892 21496 30898 21548
rect 35360 21545 35388 21576
rect 36078 21564 36084 21576
rect 36136 21604 36142 21616
rect 38924 21607 38982 21613
rect 36136 21576 38700 21604
rect 36136 21564 36142 21576
rect 33505 21539 33563 21545
rect 33505 21505 33517 21539
rect 33551 21536 33563 21539
rect 35345 21539 35403 21545
rect 35345 21536 35357 21539
rect 33551 21508 35357 21536
rect 33551 21505 33563 21508
rect 33505 21499 33563 21505
rect 35345 21505 35357 21508
rect 35391 21505 35403 21539
rect 35345 21499 35403 21505
rect 35612 21539 35670 21545
rect 35612 21505 35624 21539
rect 35658 21536 35670 21539
rect 37550 21536 37556 21548
rect 35658 21508 37556 21536
rect 35658 21505 35670 21508
rect 35612 21499 35670 21505
rect 37550 21496 37556 21508
rect 37608 21496 37614 21548
rect 38672 21545 38700 21576
rect 38924 21573 38936 21607
rect 38970 21604 38982 21607
rect 39850 21604 39856 21616
rect 38970 21576 39856 21604
rect 38970 21573 38982 21576
rect 38924 21567 38982 21573
rect 39850 21564 39856 21576
rect 39908 21564 39914 21616
rect 40764 21607 40822 21613
rect 40764 21573 40776 21607
rect 40810 21604 40822 21607
rect 42610 21604 42616 21616
rect 40810 21576 42616 21604
rect 40810 21573 40822 21576
rect 40764 21567 40822 21573
rect 42610 21564 42616 21576
rect 42668 21564 42674 21616
rect 42794 21604 42800 21616
rect 42755 21576 42800 21604
rect 42794 21564 42800 21576
rect 42852 21564 42858 21616
rect 48584 21607 48642 21613
rect 48584 21573 48596 21607
rect 48630 21604 48642 21607
rect 51552 21604 51580 21635
rect 48630 21576 51580 21604
rect 53460 21607 53518 21613
rect 48630 21573 48642 21576
rect 48584 21567 48642 21573
rect 53460 21573 53472 21607
rect 53506 21604 53518 21607
rect 53834 21604 53840 21616
rect 53506 21576 53840 21604
rect 53506 21573 53518 21576
rect 53460 21567 53518 21573
rect 53834 21564 53840 21576
rect 53892 21564 53898 21616
rect 38657 21539 38715 21545
rect 38657 21505 38669 21539
rect 38703 21505 38715 21539
rect 38657 21499 38715 21505
rect 40310 21496 40316 21548
rect 40368 21536 40374 21548
rect 40497 21539 40555 21545
rect 40497 21536 40509 21539
rect 40368 21508 40509 21536
rect 40368 21496 40374 21508
rect 40497 21505 40509 21508
rect 40543 21505 40555 21539
rect 40497 21499 40555 21505
rect 44174 21496 44180 21548
rect 44232 21536 44238 21548
rect 45261 21539 45319 21545
rect 45261 21536 45273 21539
rect 44232 21508 45273 21536
rect 44232 21496 44238 21508
rect 45261 21505 45273 21508
rect 45307 21505 45319 21539
rect 45261 21499 45319 21505
rect 48317 21539 48375 21545
rect 48317 21505 48329 21539
rect 48363 21536 48375 21539
rect 50062 21536 50068 21548
rect 48363 21508 50068 21536
rect 48363 21505 48375 21508
rect 48317 21499 48375 21505
rect 50062 21496 50068 21508
rect 50120 21496 50126 21548
rect 50424 21539 50482 21545
rect 50424 21505 50436 21539
rect 50470 21536 50482 21539
rect 51534 21536 51540 21548
rect 50470 21508 51540 21536
rect 50470 21505 50482 21508
rect 50424 21499 50482 21505
rect 51534 21496 51540 21508
rect 51592 21496 51598 21548
rect 53193 21539 53251 21545
rect 53193 21505 53205 21539
rect 53239 21536 53251 21539
rect 55033 21539 55091 21545
rect 55033 21536 55045 21539
rect 53239 21508 55045 21536
rect 53239 21505 53251 21508
rect 53193 21499 53251 21505
rect 55033 21505 55045 21508
rect 55079 21536 55091 21539
rect 55122 21536 55128 21548
rect 55079 21508 55128 21536
rect 55079 21505 55091 21508
rect 55033 21499 55091 21505
rect 55122 21496 55128 21508
rect 55180 21496 55186 21548
rect 55300 21539 55358 21545
rect 55300 21505 55312 21539
rect 55346 21536 55358 21539
rect 56686 21536 56692 21548
rect 55346 21508 56692 21536
rect 55346 21505 55358 21508
rect 55300 21499 55358 21505
rect 56686 21496 56692 21508
rect 56744 21496 56750 21548
rect 7006 21468 7012 21480
rect 6967 21440 7012 21468
rect 7006 21428 7012 21440
rect 7064 21428 7070 21480
rect 15838 21428 15844 21480
rect 15896 21468 15902 21480
rect 16669 21471 16727 21477
rect 16669 21468 16681 21471
rect 15896 21440 16681 21468
rect 15896 21428 15902 21440
rect 16669 21437 16681 21440
rect 16715 21437 16727 21471
rect 16669 21431 16727 21437
rect 23753 21471 23811 21477
rect 23753 21437 23765 21471
rect 23799 21437 23811 21471
rect 27614 21468 27620 21480
rect 27575 21440 27620 21468
rect 23753 21431 23811 21437
rect 4890 21292 4896 21344
rect 4948 21332 4954 21344
rect 5261 21335 5319 21341
rect 5261 21332 5273 21335
rect 4948 21304 5273 21332
rect 4948 21292 4954 21304
rect 5261 21301 5273 21304
rect 5307 21301 5319 21335
rect 5261 21295 5319 21301
rect 8389 21335 8447 21341
rect 8389 21301 8401 21335
rect 8435 21332 8447 21335
rect 8478 21332 8484 21344
rect 8435 21304 8484 21332
rect 8435 21301 8447 21304
rect 8389 21295 8447 21301
rect 8478 21292 8484 21304
rect 8536 21292 8542 21344
rect 13630 21332 13636 21344
rect 13591 21304 13636 21332
rect 13630 21292 13636 21304
rect 13688 21292 13694 21344
rect 18046 21332 18052 21344
rect 18007 21304 18052 21332
rect 18046 21292 18052 21304
rect 18104 21292 18110 21344
rect 19886 21332 19892 21344
rect 19847 21304 19892 21332
rect 19886 21292 19892 21304
rect 19944 21292 19950 21344
rect 23768 21332 23796 21431
rect 27614 21428 27620 21440
rect 27672 21428 27678 21480
rect 45005 21471 45063 21477
rect 45005 21468 45017 21471
rect 44100 21440 45017 21468
rect 24486 21332 24492 21344
rect 23768 21304 24492 21332
rect 24486 21292 24492 21304
rect 24544 21292 24550 21344
rect 31570 21332 31576 21344
rect 31531 21304 31576 21332
rect 31570 21292 31576 21304
rect 31628 21292 31634 21344
rect 42426 21292 42432 21344
rect 42484 21332 42490 21344
rect 44100 21341 44128 21440
rect 45005 21437 45017 21440
rect 45051 21437 45063 21471
rect 45005 21431 45063 21437
rect 50157 21471 50215 21477
rect 50157 21437 50169 21471
rect 50203 21437 50215 21471
rect 50157 21431 50215 21437
rect 44085 21335 44143 21341
rect 44085 21332 44097 21335
rect 42484 21304 44097 21332
rect 42484 21292 42490 21304
rect 44085 21301 44097 21304
rect 44131 21301 44143 21335
rect 46382 21332 46388 21344
rect 46343 21304 46388 21332
rect 44085 21295 44143 21301
rect 46382 21292 46388 21304
rect 46440 21292 46446 21344
rect 50172 21332 50200 21431
rect 51994 21332 52000 21344
rect 50172 21304 52000 21332
rect 51994 21292 52000 21304
rect 52052 21292 52058 21344
rect 54570 21332 54576 21344
rect 54531 21304 54576 21332
rect 54570 21292 54576 21304
rect 54628 21292 54634 21344
rect 56413 21335 56471 21341
rect 56413 21301 56425 21335
rect 56459 21332 56471 21335
rect 57238 21332 57244 21344
rect 56459 21304 57244 21332
rect 56459 21301 56471 21304
rect 56413 21295 56471 21301
rect 57238 21292 57244 21304
rect 57296 21292 57302 21344
rect 1104 21242 59340 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 59340 21242
rect 1104 21168 59340 21190
rect 5442 21128 5448 21140
rect 5403 21100 5448 21128
rect 5442 21088 5448 21100
rect 5500 21088 5506 21140
rect 12250 21128 12256 21140
rect 11900 21100 12256 21128
rect 4338 21020 4344 21072
rect 4396 21060 4402 21072
rect 5460 21060 5488 21088
rect 4396 21032 5488 21060
rect 4396 21020 4402 21032
rect 11900 21001 11928 21100
rect 12250 21088 12256 21100
rect 12308 21088 12314 21140
rect 13262 21128 13268 21140
rect 13223 21100 13268 21128
rect 13262 21088 13268 21100
rect 13320 21088 13326 21140
rect 15838 21128 15844 21140
rect 15120 21100 15844 21128
rect 11885 20995 11943 21001
rect 11885 20961 11897 20995
rect 11931 20961 11943 20995
rect 11885 20955 11943 20961
rect 14734 20952 14740 21004
rect 14792 20992 14798 21004
rect 15120 21001 15148 21100
rect 15838 21088 15844 21100
rect 15896 21088 15902 21140
rect 16482 21128 16488 21140
rect 16443 21100 16488 21128
rect 16482 21088 16488 21100
rect 16540 21088 16546 21140
rect 18414 21128 18420 21140
rect 18375 21100 18420 21128
rect 18414 21088 18420 21100
rect 18472 21088 18478 21140
rect 20530 21088 20536 21140
rect 20588 21128 20594 21140
rect 20625 21131 20683 21137
rect 20625 21128 20637 21131
rect 20588 21100 20637 21128
rect 20588 21088 20594 21100
rect 20625 21097 20637 21100
rect 20671 21097 20683 21131
rect 25774 21128 25780 21140
rect 25735 21100 25780 21128
rect 20625 21091 20683 21097
rect 25774 21088 25780 21100
rect 25832 21088 25838 21140
rect 27614 21128 27620 21140
rect 27448 21100 27620 21128
rect 15105 20995 15163 21001
rect 15105 20992 15117 20995
rect 14792 20964 15117 20992
rect 14792 20952 14798 20964
rect 15105 20961 15117 20964
rect 15151 20961 15163 20995
rect 18432 20992 18460 21088
rect 19242 20992 19248 21004
rect 18432 20964 19248 20992
rect 15105 20955 15163 20961
rect 19242 20952 19248 20964
rect 19300 20952 19306 21004
rect 6362 20924 6368 20936
rect 6323 20896 6368 20924
rect 6362 20884 6368 20896
rect 6420 20924 6426 20936
rect 7006 20924 7012 20936
rect 6420 20896 7012 20924
rect 6420 20884 6426 20896
rect 7006 20884 7012 20896
rect 7064 20924 7070 20936
rect 8202 20924 8208 20936
rect 7064 20896 8208 20924
rect 7064 20884 7070 20896
rect 8202 20884 8208 20896
rect 8260 20884 8266 20936
rect 8938 20924 8944 20936
rect 8899 20896 8944 20924
rect 8938 20884 8944 20896
rect 8996 20884 9002 20936
rect 12152 20927 12210 20933
rect 12152 20893 12164 20927
rect 12198 20924 12210 20927
rect 13630 20924 13636 20936
rect 12198 20896 13636 20924
rect 12198 20893 12210 20896
rect 12152 20887 12210 20893
rect 13630 20884 13636 20896
rect 13688 20884 13694 20936
rect 15372 20927 15430 20933
rect 15372 20893 15384 20927
rect 15418 20924 15430 20927
rect 16114 20924 16120 20936
rect 15418 20896 16120 20924
rect 15418 20893 15430 20896
rect 15372 20887 15430 20893
rect 16114 20884 16120 20896
rect 16172 20884 16178 20936
rect 19512 20927 19570 20933
rect 19512 20893 19524 20927
rect 19558 20924 19570 20927
rect 19886 20924 19892 20936
rect 19558 20896 19892 20924
rect 19558 20893 19570 20896
rect 19512 20887 19570 20893
rect 19886 20884 19892 20896
rect 19944 20884 19950 20936
rect 21082 20924 21088 20936
rect 21043 20896 21088 20924
rect 21082 20884 21088 20896
rect 21140 20884 21146 20936
rect 24397 20927 24455 20933
rect 24397 20893 24409 20927
rect 24443 20924 24455 20927
rect 24486 20924 24492 20936
rect 24443 20896 24492 20924
rect 24443 20893 24455 20896
rect 24397 20887 24455 20893
rect 24486 20884 24492 20896
rect 24544 20884 24550 20936
rect 26970 20884 26976 20936
rect 27028 20924 27034 20936
rect 27448 20933 27476 21100
rect 27614 21088 27620 21100
rect 27672 21088 27678 21140
rect 28810 21128 28816 21140
rect 28771 21100 28816 21128
rect 28810 21088 28816 21100
rect 28868 21088 28874 21140
rect 37550 21128 37556 21140
rect 37511 21100 37556 21128
rect 37550 21088 37556 21100
rect 37608 21088 37614 21140
rect 40218 21088 40224 21140
rect 40276 21128 40282 21140
rect 41233 21131 41291 21137
rect 41233 21128 41245 21131
rect 40276 21100 41245 21128
rect 40276 21088 40282 21100
rect 41233 21097 41245 21100
rect 41279 21097 41291 21131
rect 44082 21128 44088 21140
rect 44043 21100 44088 21128
rect 41233 21091 41291 21097
rect 44082 21088 44088 21100
rect 44140 21088 44146 21140
rect 51534 21128 51540 21140
rect 51495 21100 51540 21128
rect 51534 21088 51540 21100
rect 51592 21088 51598 21140
rect 56686 21128 56692 21140
rect 56647 21100 56692 21128
rect 56686 21088 56692 21100
rect 56744 21088 56750 21140
rect 58434 21088 58440 21140
rect 58492 21128 58498 21140
rect 58529 21131 58587 21137
rect 58529 21128 58541 21131
rect 58492 21100 58541 21128
rect 58492 21088 58498 21100
rect 58529 21097 58541 21100
rect 58575 21097 58587 21131
rect 58529 21091 58587 21097
rect 30006 20992 30012 21004
rect 29967 20964 30012 20992
rect 30006 20952 30012 20964
rect 30064 20952 30070 21004
rect 51994 20992 52000 21004
rect 51955 20964 52000 20992
rect 51994 20952 52000 20964
rect 52052 20952 52058 21004
rect 27433 20927 27491 20933
rect 27433 20924 27445 20927
rect 27028 20896 27445 20924
rect 27028 20884 27034 20896
rect 27433 20893 27445 20896
rect 27479 20893 27491 20927
rect 27433 20887 27491 20893
rect 30276 20927 30334 20933
rect 30276 20893 30288 20927
rect 30322 20924 30334 20927
rect 31570 20924 31576 20936
rect 30322 20896 31576 20924
rect 30322 20893 30334 20896
rect 30276 20887 30334 20893
rect 31570 20884 31576 20896
rect 31628 20884 31634 20936
rect 31849 20927 31907 20933
rect 31849 20893 31861 20927
rect 31895 20924 31907 20927
rect 32950 20924 32956 20936
rect 31895 20896 32956 20924
rect 31895 20893 31907 20896
rect 31849 20887 31907 20893
rect 32950 20884 32956 20896
rect 33008 20924 33014 20936
rect 34974 20924 34980 20936
rect 33008 20896 34980 20924
rect 33008 20884 33014 20896
rect 34974 20884 34980 20896
rect 35032 20884 35038 20936
rect 36078 20884 36084 20936
rect 36136 20924 36142 20936
rect 36173 20927 36231 20933
rect 36173 20924 36185 20927
rect 36136 20896 36185 20924
rect 36136 20884 36142 20896
rect 36173 20893 36185 20896
rect 36219 20893 36231 20927
rect 36173 20887 36231 20893
rect 36440 20927 36498 20933
rect 36440 20893 36452 20927
rect 36486 20924 36498 20927
rect 36722 20924 36728 20936
rect 36486 20896 36728 20924
rect 36486 20893 36498 20896
rect 36440 20887 36498 20893
rect 36722 20884 36728 20896
rect 36780 20884 36786 20936
rect 39853 20927 39911 20933
rect 39853 20893 39865 20927
rect 39899 20893 39911 20927
rect 39853 20887 39911 20893
rect 40120 20927 40178 20933
rect 40120 20893 40132 20927
rect 40166 20924 40178 20927
rect 41690 20924 41696 20936
rect 40166 20896 41696 20924
rect 40166 20893 40178 20896
rect 40120 20887 40178 20893
rect 4157 20859 4215 20865
rect 4157 20825 4169 20859
rect 4203 20856 4215 20859
rect 5258 20856 5264 20868
rect 4203 20828 5264 20856
rect 4203 20825 4215 20828
rect 4157 20819 4215 20825
rect 5258 20816 5264 20828
rect 5316 20856 5322 20868
rect 5810 20856 5816 20868
rect 5316 20828 5816 20856
rect 5316 20816 5322 20828
rect 5810 20816 5816 20828
rect 5868 20816 5874 20868
rect 6632 20859 6690 20865
rect 6632 20825 6644 20859
rect 6678 20856 6690 20859
rect 7650 20856 7656 20868
rect 6678 20828 7656 20856
rect 6678 20825 6690 20828
rect 6632 20819 6690 20825
rect 7650 20816 7656 20828
rect 7708 20816 7714 20868
rect 9208 20859 9266 20865
rect 9208 20825 9220 20859
rect 9254 20856 9266 20859
rect 10226 20856 10232 20868
rect 9254 20828 10232 20856
rect 9254 20825 9266 20828
rect 9208 20819 9266 20825
rect 10226 20816 10232 20828
rect 10284 20816 10290 20868
rect 16945 20859 17003 20865
rect 16945 20825 16957 20859
rect 16991 20825 17003 20859
rect 16945 20819 17003 20825
rect 7742 20788 7748 20800
rect 7703 20760 7748 20788
rect 7742 20748 7748 20760
rect 7800 20748 7806 20800
rect 9674 20748 9680 20800
rect 9732 20788 9738 20800
rect 10321 20791 10379 20797
rect 10321 20788 10333 20791
rect 9732 20760 10333 20788
rect 9732 20748 9738 20760
rect 10321 20757 10333 20760
rect 10367 20757 10379 20791
rect 16960 20788 16988 20819
rect 20806 20816 20812 20868
rect 20864 20856 20870 20868
rect 21330 20859 21388 20865
rect 21330 20856 21342 20859
rect 20864 20828 21342 20856
rect 20864 20816 20870 20828
rect 21330 20825 21342 20828
rect 21376 20825 21388 20859
rect 21330 20819 21388 20825
rect 24664 20859 24722 20865
rect 24664 20825 24676 20859
rect 24710 20856 24722 20859
rect 25682 20856 25688 20868
rect 24710 20828 25688 20856
rect 24710 20825 24722 20828
rect 24664 20819 24722 20825
rect 25682 20816 25688 20828
rect 25740 20816 25746 20868
rect 27700 20859 27758 20865
rect 27700 20825 27712 20859
rect 27746 20856 27758 20859
rect 28902 20856 28908 20868
rect 27746 20828 28908 20856
rect 27746 20825 27758 20828
rect 27700 20819 27758 20825
rect 28902 20816 28908 20828
rect 28960 20816 28966 20868
rect 39868 20856 39896 20887
rect 41690 20884 41696 20896
rect 41748 20884 41754 20936
rect 42426 20884 42432 20936
rect 42484 20924 42490 20936
rect 42705 20927 42763 20933
rect 42705 20924 42717 20927
rect 42484 20896 42717 20924
rect 42484 20884 42490 20896
rect 42705 20893 42717 20896
rect 42751 20893 42763 20927
rect 42705 20887 42763 20893
rect 42972 20927 43030 20933
rect 42972 20893 42984 20927
rect 43018 20924 43030 20927
rect 44450 20924 44456 20936
rect 43018 20896 44456 20924
rect 43018 20893 43030 20896
rect 42972 20887 43030 20893
rect 44450 20884 44456 20896
rect 44508 20884 44514 20936
rect 45554 20884 45560 20936
rect 45612 20924 45618 20936
rect 45649 20927 45707 20933
rect 45649 20924 45661 20927
rect 45612 20896 45661 20924
rect 45612 20884 45618 20896
rect 45649 20893 45661 20896
rect 45695 20924 45707 20927
rect 47489 20927 47547 20933
rect 47489 20924 47501 20927
rect 45695 20896 47501 20924
rect 45695 20893 45707 20896
rect 45649 20887 45707 20893
rect 47489 20893 47501 20896
rect 47535 20924 47547 20927
rect 47578 20924 47584 20936
rect 47535 20896 47584 20924
rect 47535 20893 47547 20896
rect 47489 20887 47547 20893
rect 47578 20884 47584 20896
rect 47636 20884 47642 20936
rect 50154 20924 50160 20936
rect 50067 20896 50160 20924
rect 50154 20884 50160 20896
rect 50212 20924 50218 20936
rect 50982 20924 50988 20936
rect 50212 20896 50988 20924
rect 50212 20884 50218 20896
rect 50982 20884 50988 20896
rect 51040 20884 51046 20936
rect 52264 20927 52322 20933
rect 52264 20893 52276 20927
rect 52310 20924 52322 20927
rect 54570 20924 54576 20936
rect 52310 20896 54576 20924
rect 52310 20893 52322 20896
rect 52264 20887 52322 20893
rect 54570 20884 54576 20896
rect 54628 20884 54634 20936
rect 55306 20924 55312 20936
rect 55267 20896 55312 20924
rect 55306 20884 55312 20896
rect 55364 20884 55370 20936
rect 56778 20884 56784 20936
rect 56836 20924 56842 20936
rect 57149 20927 57207 20933
rect 57149 20924 57161 20927
rect 56836 20896 57161 20924
rect 56836 20884 56842 20896
rect 57149 20893 57161 20896
rect 57195 20893 57207 20927
rect 57149 20887 57207 20893
rect 40310 20856 40316 20868
rect 39868 20828 40316 20856
rect 40310 20816 40316 20828
rect 40368 20816 40374 20868
rect 45916 20859 45974 20865
rect 45916 20825 45928 20859
rect 45962 20856 45974 20859
rect 46750 20856 46756 20868
rect 45962 20828 46756 20856
rect 45962 20825 45974 20828
rect 45916 20819 45974 20825
rect 46750 20816 46756 20828
rect 46808 20816 46814 20868
rect 47756 20859 47814 20865
rect 47756 20825 47768 20859
rect 47802 20856 47814 20859
rect 48590 20856 48596 20868
rect 47802 20828 48596 20856
rect 47802 20825 47814 20828
rect 47756 20819 47814 20825
rect 48590 20816 48596 20828
rect 48648 20816 48654 20868
rect 50424 20859 50482 20865
rect 50424 20825 50436 20859
rect 50470 20856 50482 20859
rect 50798 20856 50804 20868
rect 50470 20828 50804 20856
rect 50470 20825 50482 20828
rect 50424 20819 50482 20825
rect 50798 20816 50804 20828
rect 50856 20816 50862 20868
rect 55576 20859 55634 20865
rect 55576 20825 55588 20859
rect 55622 20856 55634 20859
rect 56686 20856 56692 20868
rect 55622 20828 56692 20856
rect 55622 20825 55634 20828
rect 55576 20819 55634 20825
rect 56686 20816 56692 20828
rect 56744 20816 56750 20868
rect 57416 20859 57474 20865
rect 57416 20825 57428 20859
rect 57462 20856 57474 20859
rect 58434 20856 58440 20868
rect 57462 20828 58440 20856
rect 57462 20825 57474 20828
rect 57416 20819 57474 20825
rect 58434 20816 58440 20828
rect 58492 20816 58498 20868
rect 20898 20788 20904 20800
rect 16960 20760 20904 20788
rect 10321 20751 10379 20757
rect 20898 20748 20904 20760
rect 20956 20748 20962 20800
rect 22462 20788 22468 20800
rect 22423 20760 22468 20788
rect 22462 20748 22468 20760
rect 22520 20748 22526 20800
rect 31386 20788 31392 20800
rect 31347 20760 31392 20788
rect 31386 20748 31392 20760
rect 31444 20748 31450 20800
rect 32490 20748 32496 20800
rect 32548 20788 32554 20800
rect 33137 20791 33195 20797
rect 33137 20788 33149 20791
rect 32548 20760 33149 20788
rect 32548 20748 32554 20760
rect 33137 20757 33149 20760
rect 33183 20757 33195 20791
rect 33137 20751 33195 20757
rect 47029 20791 47087 20797
rect 47029 20757 47041 20791
rect 47075 20788 47087 20791
rect 47302 20788 47308 20800
rect 47075 20760 47308 20788
rect 47075 20757 47087 20760
rect 47029 20751 47087 20757
rect 47302 20748 47308 20760
rect 47360 20748 47366 20800
rect 48866 20788 48872 20800
rect 48827 20760 48872 20788
rect 48866 20748 48872 20760
rect 48924 20748 48930 20800
rect 52546 20748 52552 20800
rect 52604 20788 52610 20800
rect 53377 20791 53435 20797
rect 53377 20788 53389 20791
rect 52604 20760 53389 20788
rect 52604 20748 52610 20760
rect 53377 20757 53389 20760
rect 53423 20757 53435 20791
rect 53377 20751 53435 20757
rect 1104 20698 59340 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 59340 20698
rect 1104 20624 59340 20646
rect 3881 20587 3939 20593
rect 3881 20553 3893 20587
rect 3927 20553 3939 20587
rect 3881 20547 3939 20553
rect 3896 20516 3924 20547
rect 7650 20544 7656 20596
rect 7708 20584 7714 20596
rect 7745 20587 7803 20593
rect 7745 20584 7757 20587
rect 7708 20556 7757 20584
rect 7708 20544 7714 20556
rect 7745 20553 7757 20556
rect 7791 20553 7803 20587
rect 9582 20584 9588 20596
rect 9543 20556 9588 20584
rect 7745 20547 7803 20553
rect 9582 20544 9588 20556
rect 9640 20544 9646 20596
rect 20622 20544 20628 20596
rect 20680 20584 20686 20596
rect 20901 20587 20959 20593
rect 20901 20584 20913 20587
rect 20680 20556 20913 20584
rect 20680 20544 20686 20556
rect 20901 20553 20913 20556
rect 20947 20553 20959 20587
rect 23198 20584 23204 20596
rect 23159 20556 23204 20584
rect 20901 20547 20959 20553
rect 23198 20544 23204 20556
rect 23256 20544 23262 20596
rect 33870 20584 33876 20596
rect 33831 20556 33876 20584
rect 33870 20544 33876 20556
rect 33928 20544 33934 20596
rect 40126 20584 40132 20596
rect 35866 20556 40132 20584
rect 4586 20519 4644 20525
rect 4586 20516 4598 20519
rect 3896 20488 4598 20516
rect 4586 20485 4598 20488
rect 4632 20485 4644 20519
rect 8938 20516 8944 20528
rect 4586 20479 4644 20485
rect 8220 20488 8944 20516
rect 2768 20451 2826 20457
rect 2768 20417 2780 20451
rect 2814 20448 2826 20451
rect 4890 20448 4896 20460
rect 2814 20420 4896 20448
rect 2814 20417 2826 20420
rect 2768 20411 2826 20417
rect 4890 20408 4896 20420
rect 4948 20408 4954 20460
rect 5534 20408 5540 20460
rect 5592 20448 5598 20460
rect 8220 20457 8248 20488
rect 8938 20476 8944 20488
rect 8996 20476 9002 20528
rect 11876 20519 11934 20525
rect 11876 20485 11888 20519
rect 11922 20516 11934 20519
rect 12986 20516 12992 20528
rect 11922 20488 12992 20516
rect 11922 20485 11934 20488
rect 11876 20479 11934 20485
rect 12986 20476 12992 20488
rect 13044 20476 13050 20528
rect 15004 20519 15062 20525
rect 15004 20485 15016 20519
rect 15050 20516 15062 20519
rect 18046 20516 18052 20528
rect 15050 20488 18052 20516
rect 15050 20485 15062 20488
rect 15004 20479 15062 20485
rect 18046 20476 18052 20488
rect 18104 20476 18110 20528
rect 21082 20516 21088 20528
rect 19536 20488 21088 20516
rect 6621 20451 6679 20457
rect 6621 20448 6633 20451
rect 5592 20420 6633 20448
rect 5592 20408 5598 20420
rect 6621 20417 6633 20420
rect 6667 20417 6679 20451
rect 6621 20411 6679 20417
rect 8205 20451 8263 20457
rect 8205 20417 8217 20451
rect 8251 20417 8263 20451
rect 8205 20411 8263 20417
rect 8294 20408 8300 20460
rect 8352 20448 8358 20460
rect 8461 20451 8519 20457
rect 8461 20448 8473 20451
rect 8352 20420 8473 20448
rect 8352 20408 8358 20420
rect 8461 20417 8473 20420
rect 8507 20417 8519 20451
rect 14734 20448 14740 20460
rect 14695 20420 14740 20448
rect 8461 20411 8519 20417
rect 14734 20408 14740 20420
rect 14792 20408 14798 20460
rect 17948 20451 18006 20457
rect 17948 20417 17960 20451
rect 17994 20448 18006 20451
rect 18690 20448 18696 20460
rect 17994 20420 18696 20448
rect 17994 20417 18006 20420
rect 17948 20411 18006 20417
rect 18690 20408 18696 20420
rect 18748 20408 18754 20460
rect 19334 20408 19340 20460
rect 19392 20448 19398 20460
rect 19536 20457 19564 20488
rect 21082 20476 21088 20488
rect 21140 20476 21146 20528
rect 22088 20519 22146 20525
rect 22088 20485 22100 20519
rect 22134 20516 22146 20519
rect 22462 20516 22468 20528
rect 22134 20488 22468 20516
rect 22134 20485 22146 20488
rect 22088 20479 22146 20485
rect 22462 20476 22468 20488
rect 22520 20476 22526 20528
rect 24756 20519 24814 20525
rect 24756 20485 24768 20519
rect 24802 20516 24814 20519
rect 28994 20516 29000 20528
rect 24802 20488 29000 20516
rect 24802 20485 24814 20488
rect 24756 20479 24814 20485
rect 28994 20476 29000 20488
rect 29052 20476 29058 20528
rect 32760 20519 32818 20525
rect 30208 20488 32260 20516
rect 19521 20451 19579 20457
rect 19521 20448 19533 20451
rect 19392 20420 19533 20448
rect 19392 20408 19398 20420
rect 19521 20417 19533 20420
rect 19567 20417 19579 20451
rect 19521 20411 19579 20417
rect 19788 20451 19846 20457
rect 19788 20417 19800 20451
rect 19834 20448 19846 20451
rect 20622 20448 20628 20460
rect 19834 20420 20628 20448
rect 19834 20417 19846 20420
rect 19788 20411 19846 20417
rect 20622 20408 20628 20420
rect 20680 20408 20686 20460
rect 21726 20408 21732 20460
rect 21784 20448 21790 20460
rect 21821 20451 21879 20457
rect 21821 20448 21833 20451
rect 21784 20420 21833 20448
rect 21784 20408 21790 20420
rect 21821 20417 21833 20420
rect 21867 20417 21879 20451
rect 21821 20411 21879 20417
rect 27608 20451 27666 20457
rect 27608 20417 27620 20451
rect 27654 20448 27666 20451
rect 28534 20448 28540 20460
rect 27654 20420 28540 20448
rect 27654 20417 27666 20420
rect 27608 20411 27666 20417
rect 28534 20408 28540 20420
rect 28592 20408 28598 20460
rect 30006 20408 30012 20460
rect 30064 20448 30070 20460
rect 30208 20457 30236 20488
rect 30193 20451 30251 20457
rect 30193 20448 30205 20451
rect 30064 20420 30205 20448
rect 30064 20408 30070 20420
rect 30193 20417 30205 20420
rect 30239 20417 30251 20451
rect 30193 20411 30251 20417
rect 30460 20451 30518 20457
rect 30460 20417 30472 20451
rect 30506 20448 30518 20451
rect 32122 20448 32128 20460
rect 30506 20420 32128 20448
rect 30506 20417 30518 20420
rect 30460 20411 30518 20417
rect 32122 20408 32128 20420
rect 32180 20408 32186 20460
rect 2501 20383 2559 20389
rect 2501 20349 2513 20383
rect 2547 20349 2559 20383
rect 2501 20343 2559 20349
rect 2516 20244 2544 20343
rect 4062 20340 4068 20392
rect 4120 20380 4126 20392
rect 4338 20380 4344 20392
rect 4120 20352 4344 20380
rect 4120 20340 4126 20352
rect 4338 20340 4344 20352
rect 4396 20340 4402 20392
rect 6362 20380 6368 20392
rect 6323 20352 6368 20380
rect 6362 20340 6368 20352
rect 6420 20340 6426 20392
rect 11606 20380 11612 20392
rect 11567 20352 11612 20380
rect 11606 20340 11612 20352
rect 11664 20340 11670 20392
rect 17681 20383 17739 20389
rect 17681 20349 17693 20383
rect 17727 20349 17739 20383
rect 24486 20380 24492 20392
rect 24447 20352 24492 20380
rect 17681 20343 17739 20349
rect 12894 20272 12900 20324
rect 12952 20312 12958 20324
rect 12989 20315 13047 20321
rect 12989 20312 13001 20315
rect 12952 20284 13001 20312
rect 12952 20272 12958 20284
rect 12989 20281 13001 20284
rect 13035 20281 13047 20315
rect 12989 20275 13047 20281
rect 4062 20244 4068 20256
rect 2516 20216 4068 20244
rect 4062 20204 4068 20216
rect 4120 20204 4126 20256
rect 5718 20244 5724 20256
rect 5679 20216 5724 20244
rect 5718 20204 5724 20216
rect 5776 20204 5782 20256
rect 16114 20244 16120 20256
rect 16075 20216 16120 20244
rect 16114 20204 16120 20216
rect 16172 20204 16178 20256
rect 17696 20244 17724 20343
rect 24486 20340 24492 20352
rect 24544 20340 24550 20392
rect 26970 20340 26976 20392
rect 27028 20380 27034 20392
rect 27341 20383 27399 20389
rect 27341 20380 27353 20383
rect 27028 20352 27353 20380
rect 27028 20340 27034 20352
rect 27341 20349 27353 20352
rect 27387 20349 27399 20383
rect 32232 20380 32260 20488
rect 32760 20485 32772 20519
rect 32806 20516 32818 20519
rect 33502 20516 33508 20528
rect 32806 20488 33508 20516
rect 32806 20485 32818 20488
rect 32760 20479 32818 20485
rect 33502 20476 33508 20488
rect 33560 20476 33566 20528
rect 34974 20516 34980 20528
rect 34935 20488 34980 20516
rect 34974 20476 34980 20488
rect 35032 20516 35038 20528
rect 35866 20516 35894 20556
rect 40126 20544 40132 20556
rect 40184 20544 40190 20596
rect 43809 20587 43867 20593
rect 43809 20553 43821 20587
rect 43855 20584 43867 20587
rect 44174 20584 44180 20596
rect 43855 20556 44180 20584
rect 43855 20553 43867 20556
rect 43809 20547 43867 20553
rect 44174 20544 44180 20556
rect 44232 20544 44238 20596
rect 46750 20584 46756 20596
rect 46711 20556 46756 20584
rect 46750 20544 46756 20556
rect 46808 20544 46814 20596
rect 50982 20544 50988 20596
rect 51040 20584 51046 20596
rect 51261 20587 51319 20593
rect 51261 20584 51273 20587
rect 51040 20556 51273 20584
rect 51040 20544 51046 20556
rect 51261 20553 51273 20556
rect 51307 20553 51319 20587
rect 51261 20547 51319 20553
rect 54113 20587 54171 20593
rect 54113 20553 54125 20587
rect 54159 20553 54171 20587
rect 55950 20584 55956 20596
rect 55911 20556 55956 20584
rect 54113 20547 54171 20553
rect 38654 20516 38660 20528
rect 35032 20488 35894 20516
rect 37292 20488 38660 20516
rect 35032 20476 35038 20488
rect 37292 20457 37320 20488
rect 38654 20476 38660 20488
rect 38712 20476 38718 20528
rect 49970 20516 49976 20528
rect 49931 20488 49976 20516
rect 49970 20476 49976 20488
rect 50028 20476 50034 20528
rect 54128 20516 54156 20547
rect 55950 20544 55956 20556
rect 56008 20544 56014 20596
rect 54818 20519 54876 20525
rect 54818 20516 54830 20519
rect 52748 20488 53512 20516
rect 54128 20488 54830 20516
rect 37277 20451 37335 20457
rect 37277 20417 37289 20451
rect 37323 20417 37335 20451
rect 37277 20411 37335 20417
rect 37544 20451 37602 20457
rect 37544 20417 37556 20451
rect 37590 20448 37602 20451
rect 38746 20448 38752 20460
rect 37590 20420 38752 20448
rect 37590 20417 37602 20420
rect 37544 20411 37602 20417
rect 38746 20408 38752 20420
rect 38804 20408 38810 20460
rect 40310 20408 40316 20460
rect 40368 20448 40374 20460
rect 40497 20451 40555 20457
rect 40497 20448 40509 20451
rect 40368 20420 40509 20448
rect 40368 20408 40374 20420
rect 40497 20417 40509 20420
rect 40543 20417 40555 20451
rect 40497 20411 40555 20417
rect 40764 20451 40822 20457
rect 40764 20417 40776 20451
rect 40810 20448 40822 20451
rect 41782 20448 41788 20460
rect 40810 20420 41788 20448
rect 40810 20417 40822 20420
rect 40764 20411 40822 20417
rect 41782 20408 41788 20420
rect 41840 20408 41846 20460
rect 42696 20451 42754 20457
rect 42696 20417 42708 20451
rect 42742 20448 42754 20451
rect 43714 20448 43720 20460
rect 42742 20420 43720 20448
rect 42742 20417 42754 20420
rect 42696 20411 42754 20417
rect 43714 20408 43720 20420
rect 43772 20408 43778 20460
rect 45462 20448 45468 20460
rect 45388 20420 45468 20448
rect 32490 20380 32496 20392
rect 32232 20352 32496 20380
rect 27341 20343 27399 20349
rect 32490 20340 32496 20352
rect 32548 20340 32554 20392
rect 42426 20380 42432 20392
rect 42387 20352 42432 20380
rect 42426 20340 42432 20352
rect 42484 20340 42490 20392
rect 45094 20340 45100 20392
rect 45152 20380 45158 20392
rect 45388 20389 45416 20420
rect 45462 20408 45468 20420
rect 45520 20408 45526 20460
rect 45640 20451 45698 20457
rect 45640 20417 45652 20451
rect 45686 20448 45698 20451
rect 46566 20448 46572 20460
rect 45686 20420 46572 20448
rect 45686 20417 45698 20420
rect 45640 20411 45698 20417
rect 46566 20408 46572 20420
rect 46624 20408 46630 20460
rect 47578 20408 47584 20460
rect 47636 20448 47642 20460
rect 47765 20451 47823 20457
rect 47765 20448 47777 20451
rect 47636 20420 47777 20448
rect 47636 20408 47642 20420
rect 47765 20417 47777 20420
rect 47811 20417 47823 20451
rect 47765 20411 47823 20417
rect 48032 20451 48090 20457
rect 48032 20417 48044 20451
rect 48078 20448 48090 20451
rect 48958 20448 48964 20460
rect 48078 20420 48964 20448
rect 48078 20417 48090 20420
rect 48032 20411 48090 20417
rect 48958 20408 48964 20420
rect 49016 20408 49022 20460
rect 45373 20383 45431 20389
rect 45373 20380 45385 20383
rect 45152 20352 45385 20380
rect 45152 20340 45158 20352
rect 45373 20349 45385 20352
rect 45419 20349 45431 20383
rect 45373 20343 45431 20349
rect 51994 20340 52000 20392
rect 52052 20380 52058 20392
rect 52748 20389 52776 20488
rect 53000 20451 53058 20457
rect 53000 20417 53012 20451
rect 53046 20448 53058 20451
rect 53374 20448 53380 20460
rect 53046 20420 53380 20448
rect 53046 20417 53058 20420
rect 53000 20411 53058 20417
rect 53374 20408 53380 20420
rect 53432 20408 53438 20460
rect 53484 20448 53512 20488
rect 54818 20485 54830 20488
rect 54864 20485 54876 20519
rect 54818 20479 54876 20485
rect 54570 20448 54576 20460
rect 53484 20420 54576 20448
rect 54570 20408 54576 20420
rect 54628 20408 54634 20460
rect 52733 20383 52791 20389
rect 52733 20380 52745 20383
rect 52052 20352 52745 20380
rect 52052 20340 52058 20352
rect 52733 20349 52745 20352
rect 52779 20349 52791 20383
rect 52733 20343 52791 20349
rect 19150 20312 19156 20324
rect 18616 20284 19156 20312
rect 18616 20244 18644 20284
rect 19150 20272 19156 20284
rect 19208 20272 19214 20324
rect 17696 20216 18644 20244
rect 19061 20247 19119 20253
rect 19061 20213 19073 20247
rect 19107 20244 19119 20247
rect 19334 20244 19340 20256
rect 19107 20216 19340 20244
rect 19107 20213 19119 20216
rect 19061 20207 19119 20213
rect 19334 20204 19340 20216
rect 19392 20204 19398 20256
rect 25866 20244 25872 20256
rect 25827 20216 25872 20244
rect 25866 20204 25872 20216
rect 25924 20204 25930 20256
rect 28718 20244 28724 20256
rect 28679 20216 28724 20244
rect 28718 20204 28724 20216
rect 28776 20204 28782 20256
rect 31573 20247 31631 20253
rect 31573 20213 31585 20247
rect 31619 20244 31631 20247
rect 32674 20244 32680 20256
rect 31619 20216 32680 20244
rect 31619 20213 31631 20216
rect 31573 20207 31631 20213
rect 32674 20204 32680 20216
rect 32732 20204 32738 20256
rect 36078 20204 36084 20256
rect 36136 20244 36142 20256
rect 36265 20247 36323 20253
rect 36265 20244 36277 20247
rect 36136 20216 36277 20244
rect 36136 20204 36142 20216
rect 36265 20213 36277 20216
rect 36311 20213 36323 20247
rect 36265 20207 36323 20213
rect 38657 20247 38715 20253
rect 38657 20213 38669 20247
rect 38703 20244 38715 20247
rect 38838 20244 38844 20256
rect 38703 20216 38844 20244
rect 38703 20213 38715 20216
rect 38657 20207 38715 20213
rect 38838 20204 38844 20216
rect 38896 20204 38902 20256
rect 41414 20204 41420 20256
rect 41472 20244 41478 20256
rect 41877 20247 41935 20253
rect 41877 20244 41889 20247
rect 41472 20216 41889 20244
rect 41472 20204 41478 20216
rect 41877 20213 41889 20216
rect 41923 20213 41935 20247
rect 41877 20207 41935 20213
rect 49145 20247 49203 20253
rect 49145 20213 49157 20247
rect 49191 20244 49203 20247
rect 50246 20244 50252 20256
rect 49191 20216 50252 20244
rect 49191 20213 49203 20216
rect 49145 20207 49203 20213
rect 50246 20204 50252 20216
rect 50304 20204 50310 20256
rect 1104 20154 59340 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 59340 20154
rect 1104 20080 59340 20102
rect 14458 20000 14464 20052
rect 14516 20040 14522 20052
rect 16301 20043 16359 20049
rect 16301 20040 16313 20043
rect 14516 20012 16313 20040
rect 14516 20000 14522 20012
rect 16301 20009 16313 20012
rect 16347 20009 16359 20043
rect 18690 20040 18696 20052
rect 18651 20012 18696 20040
rect 16301 20003 16359 20009
rect 18690 20000 18696 20012
rect 18748 20000 18754 20052
rect 20622 20040 20628 20052
rect 20583 20012 20628 20040
rect 20622 20000 20628 20012
rect 20680 20000 20686 20052
rect 21726 20000 21732 20052
rect 21784 20040 21790 20052
rect 22741 20043 22799 20049
rect 22741 20040 22753 20043
rect 21784 20012 22753 20040
rect 21784 20000 21790 20012
rect 22741 20009 22753 20012
rect 22787 20009 22799 20043
rect 22741 20003 22799 20009
rect 25682 20000 25688 20052
rect 25740 20040 25746 20052
rect 25777 20043 25835 20049
rect 25777 20040 25789 20043
rect 25740 20012 25789 20040
rect 25740 20000 25746 20012
rect 25777 20009 25789 20012
rect 25823 20009 25835 20043
rect 28534 20040 28540 20052
rect 28495 20012 28540 20040
rect 25777 20003 25835 20009
rect 28534 20000 28540 20012
rect 28592 20000 28598 20052
rect 32122 20040 32128 20052
rect 32083 20012 32128 20040
rect 32122 20000 32128 20012
rect 32180 20000 32186 20052
rect 36078 20040 36084 20052
rect 32600 20012 36084 20040
rect 14090 19864 14096 19916
rect 14148 19904 14154 19916
rect 14734 19904 14740 19916
rect 14148 19876 14740 19904
rect 14148 19864 14154 19876
rect 14734 19864 14740 19876
rect 14792 19904 14798 19916
rect 14921 19907 14979 19913
rect 14921 19904 14933 19907
rect 14792 19876 14933 19904
rect 14792 19864 14798 19876
rect 14921 19873 14933 19876
rect 14967 19873 14979 19907
rect 14921 19867 14979 19873
rect 30006 19864 30012 19916
rect 30064 19904 30070 19916
rect 30745 19907 30803 19913
rect 30745 19904 30757 19907
rect 30064 19876 30757 19904
rect 30064 19864 30070 19876
rect 30745 19873 30757 19876
rect 30791 19873 30803 19907
rect 30745 19867 30803 19873
rect 32122 19864 32128 19916
rect 32180 19904 32186 19916
rect 32600 19913 32628 20012
rect 34900 19913 34928 20012
rect 36078 20000 36084 20012
rect 36136 20000 36142 20052
rect 36262 20040 36268 20052
rect 36223 20012 36268 20040
rect 36262 20000 36268 20012
rect 36320 20000 36326 20052
rect 43714 20040 43720 20052
rect 43675 20012 43720 20040
rect 43714 20000 43720 20012
rect 43772 20000 43778 20052
rect 46566 20040 46572 20052
rect 46527 20012 46572 20040
rect 46566 20000 46572 20012
rect 46624 20000 46630 20052
rect 48590 20040 48596 20052
rect 48551 20012 48596 20040
rect 48590 20000 48596 20012
rect 48648 20000 48654 20052
rect 53374 20040 53380 20052
rect 53335 20012 53380 20040
rect 53374 20000 53380 20012
rect 53432 20000 53438 20052
rect 56686 20040 56692 20052
rect 56647 20012 56692 20040
rect 56686 20000 56692 20012
rect 56744 20000 56750 20052
rect 58434 20000 58440 20052
rect 58492 20040 58498 20052
rect 58529 20043 58587 20049
rect 58529 20040 58541 20043
rect 58492 20012 58541 20040
rect 58492 20000 58498 20012
rect 58529 20009 58541 20012
rect 58575 20009 58587 20043
rect 58529 20003 58587 20009
rect 32585 19907 32643 19913
rect 32585 19904 32597 19907
rect 32180 19876 32597 19904
rect 32180 19864 32186 19876
rect 32585 19873 32597 19876
rect 32631 19873 32643 19907
rect 32585 19867 32643 19873
rect 34885 19907 34943 19913
rect 34885 19873 34897 19907
rect 34931 19873 34943 19907
rect 34885 19867 34943 19873
rect 40310 19864 40316 19916
rect 40368 19904 40374 19916
rect 40497 19907 40555 19913
rect 40497 19904 40509 19907
rect 40368 19876 40509 19904
rect 40368 19864 40374 19876
rect 40497 19873 40509 19876
rect 40543 19873 40555 19907
rect 50154 19904 50160 19916
rect 50115 19876 50160 19904
rect 40497 19867 40555 19873
rect 4341 19839 4399 19845
rect 4341 19805 4353 19839
rect 4387 19805 4399 19839
rect 4341 19799 4399 19805
rect 4608 19839 4666 19845
rect 4608 19805 4620 19839
rect 4654 19836 4666 19839
rect 5718 19836 5724 19848
rect 4654 19808 5724 19836
rect 4654 19805 4666 19808
rect 4608 19799 4666 19805
rect 4356 19768 4384 19799
rect 5718 19796 5724 19808
rect 5776 19796 5782 19848
rect 5810 19796 5816 19848
rect 5868 19836 5874 19848
rect 6641 19839 6699 19845
rect 6641 19836 6653 19839
rect 5868 19808 6653 19836
rect 5868 19796 5874 19808
rect 6641 19805 6653 19808
rect 6687 19805 6699 19839
rect 8938 19836 8944 19848
rect 8899 19808 8944 19836
rect 6641 19799 6699 19805
rect 8938 19796 8944 19808
rect 8996 19796 9002 19848
rect 11517 19839 11575 19845
rect 11517 19805 11529 19839
rect 11563 19836 11575 19839
rect 11606 19836 11612 19848
rect 11563 19808 11612 19836
rect 11563 19805 11575 19808
rect 11517 19799 11575 19805
rect 11606 19796 11612 19808
rect 11664 19796 11670 19848
rect 15188 19839 15246 19845
rect 15188 19805 15200 19839
rect 15234 19836 15246 19839
rect 16114 19836 16120 19848
rect 15234 19808 16120 19836
rect 15234 19805 15246 19808
rect 15188 19799 15246 19805
rect 16114 19796 16120 19808
rect 16172 19796 16178 19848
rect 17310 19836 17316 19848
rect 17271 19808 17316 19836
rect 17310 19796 17316 19808
rect 17368 19796 17374 19848
rect 19242 19836 19248 19848
rect 19203 19808 19248 19836
rect 19242 19796 19248 19808
rect 19300 19796 19306 19848
rect 19334 19796 19340 19848
rect 19392 19836 19398 19848
rect 19501 19839 19559 19845
rect 19501 19836 19513 19839
rect 19392 19808 19513 19836
rect 19392 19796 19398 19808
rect 19501 19805 19513 19808
rect 19547 19805 19559 19839
rect 19501 19799 19559 19805
rect 23658 19796 23664 19848
rect 23716 19836 23722 19848
rect 24397 19839 24455 19845
rect 24397 19836 24409 19839
rect 23716 19808 24409 19836
rect 23716 19796 23722 19808
rect 24397 19805 24409 19808
rect 24443 19836 24455 19839
rect 24486 19836 24492 19848
rect 24443 19808 24492 19836
rect 24443 19805 24455 19808
rect 24397 19799 24455 19805
rect 24486 19796 24492 19808
rect 24544 19796 24550 19848
rect 24664 19839 24722 19845
rect 24664 19805 24676 19839
rect 24710 19836 24722 19839
rect 25866 19836 25872 19848
rect 24710 19808 25872 19836
rect 24710 19805 24722 19808
rect 24664 19799 24722 19805
rect 25866 19796 25872 19808
rect 25924 19796 25930 19848
rect 26970 19796 26976 19848
rect 27028 19836 27034 19848
rect 27157 19839 27215 19845
rect 27157 19836 27169 19839
rect 27028 19808 27169 19836
rect 27028 19796 27034 19808
rect 27157 19805 27169 19808
rect 27203 19805 27215 19839
rect 27157 19799 27215 19805
rect 31012 19839 31070 19845
rect 31012 19805 31024 19839
rect 31058 19836 31070 19839
rect 31386 19836 31392 19848
rect 31058 19808 31392 19836
rect 31058 19805 31070 19808
rect 31012 19799 31070 19805
rect 31386 19796 31392 19808
rect 31444 19796 31450 19848
rect 32674 19796 32680 19848
rect 32732 19836 32738 19848
rect 32841 19839 32899 19845
rect 32841 19836 32853 19839
rect 32732 19808 32853 19836
rect 32732 19796 32738 19808
rect 32841 19805 32853 19808
rect 32887 19805 32899 19839
rect 32841 19799 32899 19805
rect 35152 19839 35210 19845
rect 35152 19805 35164 19839
rect 35198 19836 35210 19839
rect 36630 19836 36636 19848
rect 35198 19808 36636 19836
rect 35198 19805 35210 19808
rect 35152 19799 35210 19805
rect 36630 19796 36636 19808
rect 36688 19796 36694 19848
rect 37829 19839 37887 19845
rect 37829 19805 37841 19839
rect 37875 19836 37887 19839
rect 38654 19836 38660 19848
rect 37875 19808 38660 19836
rect 37875 19805 37887 19808
rect 37829 19799 37887 19805
rect 38654 19796 38660 19808
rect 38712 19796 38718 19848
rect 40512 19836 40540 19867
rect 50154 19864 50160 19876
rect 50212 19864 50218 19916
rect 51994 19904 52000 19916
rect 51955 19876 52000 19904
rect 51994 19864 52000 19876
rect 52052 19864 52058 19916
rect 42337 19839 42395 19845
rect 42337 19836 42349 19839
rect 40512 19808 42349 19836
rect 42337 19805 42349 19808
rect 42383 19836 42395 19839
rect 42426 19836 42432 19848
rect 42383 19808 42432 19836
rect 42383 19805 42395 19808
rect 42337 19799 42395 19805
rect 42426 19796 42432 19808
rect 42484 19796 42490 19848
rect 45094 19796 45100 19848
rect 45152 19836 45158 19848
rect 45189 19839 45247 19845
rect 45189 19836 45201 19839
rect 45152 19808 45201 19836
rect 45152 19796 45158 19808
rect 45189 19805 45201 19808
rect 45235 19805 45247 19839
rect 47210 19836 47216 19848
rect 47171 19808 47216 19836
rect 45189 19799 45247 19805
rect 47210 19796 47216 19808
rect 47268 19796 47274 19848
rect 47302 19796 47308 19848
rect 47360 19836 47366 19848
rect 47469 19839 47527 19845
rect 47469 19836 47481 19839
rect 47360 19808 47481 19836
rect 47360 19796 47366 19808
rect 47469 19805 47481 19808
rect 47515 19805 47527 19839
rect 47469 19799 47527 19805
rect 50246 19796 50252 19848
rect 50304 19836 50310 19848
rect 50413 19839 50471 19845
rect 50413 19836 50425 19839
rect 50304 19808 50425 19836
rect 50304 19796 50310 19808
rect 50413 19805 50425 19808
rect 50459 19805 50471 19839
rect 50413 19799 50471 19805
rect 52264 19839 52322 19845
rect 52264 19805 52276 19839
rect 52310 19836 52322 19839
rect 52546 19836 52552 19848
rect 52310 19808 52552 19836
rect 52310 19805 52322 19808
rect 52264 19799 52322 19805
rect 52546 19796 52552 19808
rect 52604 19796 52610 19848
rect 54570 19796 54576 19848
rect 54628 19836 54634 19848
rect 55306 19836 55312 19848
rect 54628 19808 55312 19836
rect 54628 19796 54634 19808
rect 55306 19796 55312 19808
rect 55364 19796 55370 19848
rect 55398 19796 55404 19848
rect 55456 19836 55462 19848
rect 55565 19839 55623 19845
rect 55565 19836 55577 19839
rect 55456 19808 55577 19836
rect 55456 19796 55462 19808
rect 55565 19805 55577 19808
rect 55611 19805 55623 19839
rect 55565 19799 55623 19805
rect 55858 19796 55864 19848
rect 55916 19836 55922 19848
rect 57149 19839 57207 19845
rect 57149 19836 57161 19839
rect 55916 19808 57161 19836
rect 55916 19796 55922 19808
rect 57149 19805 57161 19808
rect 57195 19805 57207 19839
rect 57149 19799 57207 19805
rect 57238 19796 57244 19848
rect 57296 19836 57302 19848
rect 57405 19839 57463 19845
rect 57405 19836 57417 19839
rect 57296 19808 57417 19836
rect 57296 19796 57302 19808
rect 57405 19805 57417 19808
rect 57451 19805 57463 19839
rect 57405 19799 57463 19805
rect 8202 19768 8208 19780
rect 4356 19740 4660 19768
rect 8163 19740 8208 19768
rect 4632 19712 4660 19740
rect 8202 19728 8208 19740
rect 8260 19728 8266 19780
rect 9208 19771 9266 19777
rect 9208 19737 9220 19771
rect 9254 19768 9266 19771
rect 9582 19768 9588 19780
rect 9254 19740 9588 19768
rect 9254 19737 9266 19740
rect 9208 19731 9266 19737
rect 9582 19728 9588 19740
rect 9640 19728 9646 19780
rect 11784 19771 11842 19777
rect 11784 19737 11796 19771
rect 11830 19768 11842 19771
rect 12802 19768 12808 19780
rect 11830 19740 12808 19768
rect 11830 19737 11842 19740
rect 11784 19731 11842 19737
rect 12802 19728 12808 19740
rect 12860 19728 12866 19780
rect 17580 19771 17638 19777
rect 17580 19737 17592 19771
rect 17626 19768 17638 19771
rect 18690 19768 18696 19780
rect 17626 19740 18696 19768
rect 17626 19737 17638 19740
rect 17580 19731 17638 19737
rect 18690 19728 18696 19740
rect 18748 19728 18754 19780
rect 20898 19728 20904 19780
rect 20956 19768 20962 19780
rect 21453 19771 21511 19777
rect 21453 19768 21465 19771
rect 20956 19740 21465 19768
rect 20956 19728 20962 19740
rect 21453 19737 21465 19740
rect 21499 19768 21511 19771
rect 25958 19768 25964 19780
rect 21499 19740 25964 19768
rect 21499 19737 21511 19740
rect 21453 19731 21511 19737
rect 25958 19728 25964 19740
rect 26016 19728 26022 19780
rect 27424 19771 27482 19777
rect 27424 19737 27436 19771
rect 27470 19768 27482 19771
rect 28350 19768 28356 19780
rect 27470 19740 28356 19768
rect 27470 19737 27482 19740
rect 27424 19731 27482 19737
rect 28350 19728 28356 19740
rect 28408 19728 28414 19780
rect 38096 19771 38154 19777
rect 38096 19737 38108 19771
rect 38142 19768 38154 19771
rect 39114 19768 39120 19780
rect 38142 19740 39120 19768
rect 38142 19737 38154 19740
rect 38096 19731 38154 19737
rect 39114 19728 39120 19740
rect 39172 19728 39178 19780
rect 40764 19771 40822 19777
rect 40764 19737 40776 19771
rect 40810 19768 40822 19771
rect 42604 19771 42662 19777
rect 40810 19740 42564 19768
rect 40810 19737 40822 19740
rect 40764 19731 40822 19737
rect 4614 19660 4620 19712
rect 4672 19660 4678 19712
rect 5718 19700 5724 19712
rect 5679 19672 5724 19700
rect 5718 19660 5724 19672
rect 5776 19660 5782 19712
rect 10318 19700 10324 19712
rect 10279 19672 10324 19700
rect 10318 19660 10324 19672
rect 10376 19660 10382 19712
rect 12894 19700 12900 19712
rect 12855 19672 12900 19700
rect 12894 19660 12900 19672
rect 12952 19660 12958 19712
rect 31754 19660 31760 19712
rect 31812 19700 31818 19712
rect 33965 19703 34023 19709
rect 33965 19700 33977 19703
rect 31812 19672 33977 19700
rect 31812 19660 31818 19672
rect 33965 19669 33977 19672
rect 34011 19669 34023 19703
rect 33965 19663 34023 19669
rect 37826 19660 37832 19712
rect 37884 19700 37890 19712
rect 39209 19703 39267 19709
rect 39209 19700 39221 19703
rect 37884 19672 39221 19700
rect 37884 19660 37890 19672
rect 39209 19669 39221 19672
rect 39255 19669 39267 19703
rect 41874 19700 41880 19712
rect 41835 19672 41880 19700
rect 39209 19663 39267 19669
rect 41874 19660 41880 19672
rect 41932 19660 41938 19712
rect 42536 19700 42564 19740
rect 42604 19737 42616 19771
rect 42650 19768 42662 19771
rect 43806 19768 43812 19780
rect 42650 19740 43812 19768
rect 42650 19737 42662 19740
rect 42604 19731 42662 19737
rect 43806 19728 43812 19740
rect 43864 19728 43870 19780
rect 45456 19771 45514 19777
rect 45456 19737 45468 19771
rect 45502 19768 45514 19771
rect 46566 19768 46572 19780
rect 45502 19740 46572 19768
rect 45502 19737 45514 19740
rect 45456 19731 45514 19737
rect 46566 19728 46572 19740
rect 46624 19728 46630 19780
rect 55324 19768 55352 19796
rect 55876 19768 55904 19796
rect 55324 19740 55904 19768
rect 46382 19700 46388 19712
rect 42536 19672 46388 19700
rect 46382 19660 46388 19672
rect 46440 19660 46446 19712
rect 51534 19700 51540 19712
rect 51495 19672 51540 19700
rect 51534 19660 51540 19672
rect 51592 19660 51598 19712
rect 1104 19610 59340 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 59340 19610
rect 1104 19536 59340 19558
rect 9582 19496 9588 19508
rect 4264 19468 8616 19496
rect 9543 19468 9588 19496
rect 1848 19431 1906 19437
rect 1848 19397 1860 19431
rect 1894 19428 1906 19431
rect 4264 19428 4292 19468
rect 1894 19400 4292 19428
rect 4332 19431 4390 19437
rect 1894 19397 1906 19400
rect 1848 19391 1906 19397
rect 4332 19397 4344 19431
rect 4378 19428 4390 19431
rect 5718 19428 5724 19440
rect 4378 19400 5724 19428
rect 4378 19397 4390 19400
rect 4332 19391 4390 19397
rect 5718 19388 5724 19400
rect 5776 19388 5782 19440
rect 6632 19431 6690 19437
rect 6632 19397 6644 19431
rect 6678 19428 6690 19431
rect 7742 19428 7748 19440
rect 6678 19400 7748 19428
rect 6678 19397 6690 19400
rect 6632 19391 6690 19397
rect 7742 19388 7748 19400
rect 7800 19388 7806 19440
rect 8588 19428 8616 19468
rect 9582 19456 9588 19468
rect 9640 19456 9646 19508
rect 18690 19496 18696 19508
rect 18651 19468 18696 19496
rect 18690 19456 18696 19468
rect 18748 19456 18754 19508
rect 19242 19456 19248 19508
rect 19300 19496 19306 19508
rect 21269 19499 21327 19505
rect 19300 19468 19932 19496
rect 19300 19456 19306 19468
rect 9674 19428 9680 19440
rect 8588 19400 9680 19428
rect 9674 19388 9680 19400
rect 9732 19388 9738 19440
rect 12894 19388 12900 19440
rect 12952 19428 12958 19440
rect 13602 19431 13660 19437
rect 13602 19428 13614 19431
rect 12952 19400 13614 19428
rect 12952 19388 12958 19400
rect 13602 19397 13614 19400
rect 13648 19397 13660 19431
rect 13602 19391 13660 19397
rect 19904 19428 19932 19468
rect 21269 19465 21281 19499
rect 21315 19465 21327 19499
rect 28350 19496 28356 19508
rect 28311 19468 28356 19496
rect 21269 19459 21327 19465
rect 20714 19428 20720 19440
rect 19904 19400 20720 19428
rect 1578 19360 1584 19372
rect 1491 19332 1584 19360
rect 1578 19320 1584 19332
rect 1636 19360 1642 19372
rect 4062 19360 4068 19372
rect 1636 19332 4068 19360
rect 1636 19320 1642 19332
rect 4062 19320 4068 19332
rect 4120 19320 4126 19372
rect 5534 19360 5540 19372
rect 5460 19332 5540 19360
rect 5460 19233 5488 19332
rect 5534 19320 5540 19332
rect 5592 19320 5598 19372
rect 8202 19360 8208 19372
rect 8163 19332 8208 19360
rect 8202 19320 8208 19332
rect 8260 19320 8266 19372
rect 8478 19369 8484 19372
rect 8472 19360 8484 19369
rect 8439 19332 8484 19360
rect 8472 19323 8484 19332
rect 8478 19320 8484 19323
rect 8536 19320 8542 19372
rect 11517 19363 11575 19369
rect 11517 19329 11529 19363
rect 11563 19360 11575 19363
rect 11606 19360 11612 19372
rect 11563 19332 11612 19360
rect 11563 19329 11575 19332
rect 11517 19323 11575 19329
rect 11606 19320 11612 19332
rect 11664 19320 11670 19372
rect 11784 19363 11842 19369
rect 11784 19329 11796 19363
rect 11830 19360 11842 19363
rect 12710 19360 12716 19372
rect 11830 19332 12716 19360
rect 11830 19329 11842 19332
rect 11784 19323 11842 19329
rect 12710 19320 12716 19332
rect 12768 19320 12774 19372
rect 12802 19320 12808 19372
rect 12860 19360 12866 19372
rect 13357 19363 13415 19369
rect 12860 19332 12940 19360
rect 12860 19320 12866 19332
rect 6362 19292 6368 19304
rect 6323 19264 6368 19292
rect 6362 19252 6368 19264
rect 6420 19252 6426 19304
rect 12912 19233 12940 19332
rect 13357 19329 13369 19363
rect 13403 19360 13415 19363
rect 13906 19360 13912 19372
rect 13403 19332 13912 19360
rect 13403 19329 13415 19332
rect 13357 19323 13415 19329
rect 13906 19320 13912 19332
rect 13964 19320 13970 19372
rect 17310 19360 17316 19372
rect 17271 19332 17316 19360
rect 17310 19320 17316 19332
rect 17368 19320 17374 19372
rect 17580 19363 17638 19369
rect 17580 19329 17592 19363
rect 17626 19360 17638 19363
rect 19242 19360 19248 19372
rect 17626 19332 19248 19360
rect 17626 19329 17638 19332
rect 17580 19323 17638 19329
rect 19242 19320 19248 19332
rect 19300 19320 19306 19372
rect 19904 19369 19932 19400
rect 20714 19388 20720 19400
rect 20772 19388 20778 19440
rect 21284 19428 21312 19459
rect 28350 19456 28356 19468
rect 28408 19456 28414 19508
rect 31573 19499 31631 19505
rect 31573 19465 31585 19499
rect 31619 19465 31631 19499
rect 31573 19459 31631 19465
rect 22066 19431 22124 19437
rect 22066 19428 22078 19431
rect 21284 19400 22078 19428
rect 22066 19397 22078 19400
rect 22112 19397 22124 19431
rect 22066 19391 22124 19397
rect 27240 19431 27298 19437
rect 27240 19397 27252 19431
rect 27286 19428 27298 19431
rect 31202 19428 31208 19440
rect 27286 19400 31208 19428
rect 27286 19397 27298 19400
rect 27240 19391 27298 19397
rect 31202 19388 31208 19400
rect 31260 19388 31266 19440
rect 31588 19428 31616 19459
rect 34514 19456 34520 19508
rect 34572 19496 34578 19508
rect 36541 19499 36599 19505
rect 36541 19496 36553 19499
rect 34572 19468 36553 19496
rect 34572 19456 34578 19468
rect 36541 19465 36553 19468
rect 36587 19465 36599 19499
rect 43806 19496 43812 19508
rect 43767 19468 43812 19496
rect 36541 19459 36599 19465
rect 43806 19456 43812 19468
rect 43864 19456 43870 19508
rect 46566 19496 46572 19508
rect 46527 19468 46572 19496
rect 46566 19456 46572 19468
rect 46624 19456 46630 19508
rect 48958 19496 48964 19508
rect 48919 19468 48964 19496
rect 48958 19456 48964 19468
rect 49016 19456 49022 19508
rect 50798 19496 50804 19508
rect 50759 19468 50804 19496
rect 50798 19456 50804 19468
rect 50856 19456 50862 19508
rect 32370 19431 32428 19437
rect 32370 19428 32382 19431
rect 31588 19400 32382 19428
rect 32370 19397 32382 19400
rect 32416 19397 32428 19431
rect 36078 19428 36084 19440
rect 32370 19391 32428 19397
rect 35176 19400 36084 19428
rect 19889 19363 19947 19369
rect 19889 19329 19901 19363
rect 19935 19329 19947 19363
rect 19889 19323 19947 19329
rect 20156 19363 20214 19369
rect 20156 19329 20168 19363
rect 20202 19360 20214 19363
rect 21266 19360 21272 19372
rect 20202 19332 21272 19360
rect 20202 19329 20214 19332
rect 20156 19323 20214 19329
rect 21266 19320 21272 19332
rect 21324 19320 21330 19372
rect 21818 19360 21824 19372
rect 21779 19332 21824 19360
rect 21818 19320 21824 19332
rect 21876 19360 21882 19372
rect 21876 19332 23428 19360
rect 21876 19320 21882 19332
rect 23400 19292 23428 19332
rect 23474 19320 23480 19372
rect 23532 19360 23538 19372
rect 23917 19363 23975 19369
rect 23917 19360 23929 19363
rect 23532 19332 23929 19360
rect 23532 19320 23538 19332
rect 23917 19329 23929 19332
rect 23963 19329 23975 19363
rect 26970 19360 26976 19372
rect 26931 19332 26976 19360
rect 23917 19323 23975 19329
rect 26970 19320 26976 19332
rect 27028 19320 27034 19372
rect 30006 19320 30012 19372
rect 30064 19360 30070 19372
rect 30193 19363 30251 19369
rect 30193 19360 30205 19363
rect 30064 19332 30205 19360
rect 30064 19320 30070 19332
rect 30193 19329 30205 19332
rect 30239 19329 30251 19363
rect 30193 19323 30251 19329
rect 30460 19363 30518 19369
rect 30460 19329 30472 19363
rect 30506 19360 30518 19363
rect 32214 19360 32220 19372
rect 30506 19332 32220 19360
rect 30506 19329 30518 19332
rect 30460 19323 30518 19329
rect 32214 19320 32220 19332
rect 32272 19320 32278 19372
rect 35176 19369 35204 19400
rect 36078 19388 36084 19400
rect 36136 19388 36142 19440
rect 39850 19428 39856 19440
rect 38856 19400 39856 19428
rect 35161 19363 35219 19369
rect 35161 19329 35173 19363
rect 35207 19329 35219 19363
rect 35161 19323 35219 19329
rect 35428 19363 35486 19369
rect 35428 19329 35440 19363
rect 35474 19360 35486 19363
rect 36722 19360 36728 19372
rect 35474 19332 36728 19360
rect 35474 19329 35486 19332
rect 35428 19323 35486 19329
rect 36722 19320 36728 19332
rect 36780 19320 36786 19372
rect 38856 19360 38884 19400
rect 39850 19388 39856 19400
rect 39908 19388 39914 19440
rect 40764 19431 40822 19437
rect 40764 19397 40776 19431
rect 40810 19428 40822 19431
rect 41874 19428 41880 19440
rect 40810 19400 41880 19428
rect 40810 19397 40822 19400
rect 40764 19391 40822 19397
rect 41874 19388 41880 19400
rect 41932 19388 41938 19440
rect 47848 19431 47906 19437
rect 47848 19397 47860 19431
rect 47894 19428 47906 19431
rect 48866 19428 48872 19440
rect 47894 19400 48872 19428
rect 47894 19397 47906 19400
rect 47848 19391 47906 19397
rect 48866 19388 48872 19400
rect 48924 19388 48930 19440
rect 49688 19431 49746 19437
rect 49688 19397 49700 19431
rect 49734 19428 49746 19431
rect 51534 19428 51540 19440
rect 49734 19400 51540 19428
rect 49734 19397 49746 19400
rect 49688 19391 49746 19397
rect 51534 19388 51540 19400
rect 51592 19388 51598 19440
rect 54021 19431 54079 19437
rect 54021 19397 54033 19431
rect 54067 19428 54079 19431
rect 55674 19428 55680 19440
rect 54067 19400 55680 19428
rect 54067 19397 54079 19400
rect 54021 19391 54079 19397
rect 55674 19388 55680 19400
rect 55732 19388 55738 19440
rect 55769 19431 55827 19437
rect 55769 19397 55781 19431
rect 55815 19428 55827 19431
rect 55858 19428 55864 19440
rect 55815 19400 55864 19428
rect 55815 19397 55827 19400
rect 55769 19391 55827 19397
rect 55858 19388 55864 19400
rect 55916 19388 55922 19440
rect 38764 19332 38884 19360
rect 38924 19363 38982 19369
rect 23658 19292 23664 19304
rect 23400 19264 23664 19292
rect 23658 19252 23664 19264
rect 23716 19252 23722 19304
rect 32122 19292 32128 19304
rect 32083 19264 32128 19292
rect 32122 19252 32128 19264
rect 32180 19252 32186 19304
rect 38286 19252 38292 19304
rect 38344 19292 38350 19304
rect 38654 19292 38660 19304
rect 38344 19264 38660 19292
rect 38344 19252 38350 19264
rect 38654 19252 38660 19264
rect 38712 19292 38718 19304
rect 38764 19292 38792 19332
rect 38924 19329 38936 19363
rect 38970 19360 38982 19363
rect 41230 19360 41236 19372
rect 38970 19332 41236 19360
rect 38970 19329 38982 19332
rect 38924 19323 38982 19329
rect 41230 19320 41236 19332
rect 41288 19320 41294 19372
rect 41782 19320 41788 19372
rect 41840 19360 41846 19372
rect 42426 19360 42432 19372
rect 41840 19332 41920 19360
rect 42387 19332 42432 19360
rect 41840 19320 41846 19332
rect 38712 19264 38792 19292
rect 40497 19295 40555 19301
rect 38712 19252 38718 19264
rect 40497 19261 40509 19295
rect 40543 19261 40555 19295
rect 40497 19255 40555 19261
rect 5445 19227 5503 19233
rect 5445 19193 5457 19227
rect 5491 19193 5503 19227
rect 5445 19187 5503 19193
rect 12897 19227 12955 19233
rect 12897 19193 12909 19227
rect 12943 19193 12955 19227
rect 12897 19187 12955 19193
rect 39850 19184 39856 19236
rect 39908 19224 39914 19236
rect 40512 19224 40540 19255
rect 41892 19233 41920 19332
rect 42426 19320 42432 19332
rect 42484 19320 42490 19372
rect 42696 19363 42754 19369
rect 42696 19329 42708 19363
rect 42742 19360 42754 19363
rect 43714 19360 43720 19372
rect 42742 19332 43720 19360
rect 42742 19329 42754 19332
rect 42696 19323 42754 19329
rect 43714 19320 43720 19332
rect 43772 19320 43778 19372
rect 45456 19363 45514 19369
rect 45456 19329 45468 19363
rect 45502 19360 45514 19363
rect 46474 19360 46480 19372
rect 45502 19332 46480 19360
rect 45502 19329 45514 19332
rect 45456 19323 45514 19329
rect 46474 19320 46480 19332
rect 46532 19320 46538 19372
rect 47210 19320 47216 19372
rect 47268 19360 47274 19372
rect 47581 19363 47639 19369
rect 47581 19360 47593 19363
rect 47268 19332 47593 19360
rect 47268 19320 47274 19332
rect 47581 19329 47593 19332
rect 47627 19360 47639 19363
rect 49421 19363 49479 19369
rect 49421 19360 49433 19363
rect 47627 19332 49433 19360
rect 47627 19329 47639 19332
rect 47581 19323 47639 19329
rect 49421 19329 49433 19332
rect 49467 19360 49479 19363
rect 50154 19360 50160 19372
rect 49467 19332 50160 19360
rect 49467 19329 49479 19332
rect 49421 19323 49479 19329
rect 50154 19320 50160 19332
rect 50212 19320 50218 19372
rect 45094 19252 45100 19304
rect 45152 19292 45158 19304
rect 45189 19295 45247 19301
rect 45189 19292 45201 19295
rect 45152 19264 45201 19292
rect 45152 19252 45158 19264
rect 45189 19261 45201 19264
rect 45235 19261 45247 19295
rect 45189 19255 45247 19261
rect 39908 19196 40540 19224
rect 39908 19184 39914 19196
rect 2958 19156 2964 19168
rect 2919 19128 2964 19156
rect 2958 19116 2964 19128
rect 3016 19116 3022 19168
rect 7742 19156 7748 19168
rect 7703 19128 7748 19156
rect 7742 19116 7748 19128
rect 7800 19116 7806 19168
rect 13998 19116 14004 19168
rect 14056 19156 14062 19168
rect 14737 19159 14795 19165
rect 14737 19156 14749 19159
rect 14056 19128 14749 19156
rect 14056 19116 14062 19128
rect 14737 19125 14749 19128
rect 14783 19125 14795 19159
rect 23198 19156 23204 19168
rect 23159 19128 23204 19156
rect 14737 19119 14795 19125
rect 23198 19116 23204 19128
rect 23256 19116 23262 19168
rect 25038 19156 25044 19168
rect 24999 19128 25044 19156
rect 25038 19116 25044 19128
rect 25096 19116 25102 19168
rect 33502 19156 33508 19168
rect 33463 19128 33508 19156
rect 33502 19116 33508 19128
rect 33560 19116 33566 19168
rect 38654 19116 38660 19168
rect 38712 19156 38718 19168
rect 40037 19159 40095 19165
rect 40037 19156 40049 19159
rect 38712 19128 40049 19156
rect 38712 19116 38718 19128
rect 40037 19125 40049 19128
rect 40083 19125 40095 19159
rect 40512 19156 40540 19196
rect 41877 19227 41935 19233
rect 41877 19193 41889 19227
rect 41923 19193 41935 19227
rect 41877 19187 41935 19193
rect 41506 19156 41512 19168
rect 40512 19128 41512 19156
rect 40037 19119 40095 19125
rect 41506 19116 41512 19128
rect 41564 19116 41570 19168
rect 1104 19066 59340 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 59340 19066
rect 1104 18992 59340 19014
rect 10226 18912 10232 18964
rect 10284 18952 10290 18964
rect 10321 18955 10379 18961
rect 10321 18952 10333 18955
rect 10284 18924 10333 18952
rect 10284 18912 10290 18924
rect 10321 18921 10333 18924
rect 10367 18921 10379 18955
rect 10321 18915 10379 18921
rect 32214 18912 32220 18964
rect 32272 18952 32278 18964
rect 32493 18955 32551 18961
rect 32493 18952 32505 18955
rect 32272 18924 32505 18952
rect 32272 18912 32278 18924
rect 32493 18921 32505 18924
rect 32539 18921 32551 18955
rect 41230 18952 41236 18964
rect 41191 18924 41236 18952
rect 32493 18915 32551 18921
rect 41230 18912 41236 18924
rect 41288 18912 41294 18964
rect 43714 18952 43720 18964
rect 43675 18924 43720 18952
rect 43714 18912 43720 18924
rect 43772 18912 43778 18964
rect 46474 18952 46480 18964
rect 46435 18924 46480 18952
rect 46474 18912 46480 18924
rect 46532 18912 46538 18964
rect 1578 18816 1584 18828
rect 1539 18788 1584 18816
rect 1578 18776 1584 18788
rect 1636 18776 1642 18828
rect 39850 18816 39856 18828
rect 39811 18788 39856 18816
rect 39850 18776 39856 18788
rect 39908 18776 39914 18828
rect 1848 18751 1906 18757
rect 1848 18717 1860 18751
rect 1894 18748 1906 18751
rect 2958 18748 2964 18760
rect 1894 18720 2964 18748
rect 1894 18717 1906 18720
rect 1848 18711 1906 18717
rect 2958 18708 2964 18720
rect 3016 18708 3022 18760
rect 6362 18748 6368 18760
rect 6323 18720 6368 18748
rect 6362 18708 6368 18720
rect 6420 18708 6426 18760
rect 6632 18751 6690 18757
rect 6632 18717 6644 18751
rect 6678 18748 6690 18751
rect 7742 18748 7748 18760
rect 6678 18720 7748 18748
rect 6678 18717 6690 18720
rect 6632 18711 6690 18717
rect 7742 18708 7748 18720
rect 7800 18708 7806 18760
rect 8938 18748 8944 18760
rect 8899 18720 8944 18748
rect 8938 18708 8944 18720
rect 8996 18708 9002 18760
rect 9208 18751 9266 18757
rect 9208 18717 9220 18751
rect 9254 18748 9266 18751
rect 10318 18748 10324 18760
rect 9254 18720 10324 18748
rect 9254 18717 9266 18720
rect 9208 18711 9266 18717
rect 10318 18708 10324 18720
rect 10376 18708 10382 18760
rect 11514 18748 11520 18760
rect 11475 18720 11520 18748
rect 11514 18708 11520 18720
rect 11572 18708 11578 18760
rect 11606 18708 11612 18760
rect 11664 18748 11670 18760
rect 13265 18751 13323 18757
rect 13265 18748 13277 18751
rect 11664 18720 13277 18748
rect 11664 18708 11670 18720
rect 13265 18717 13277 18720
rect 13311 18748 13323 18751
rect 13906 18748 13912 18760
rect 13311 18720 13912 18748
rect 13311 18717 13323 18720
rect 13265 18711 13323 18717
rect 13906 18708 13912 18720
rect 13964 18748 13970 18760
rect 14093 18751 14151 18757
rect 14093 18748 14105 18751
rect 13964 18720 14105 18748
rect 13964 18708 13970 18720
rect 14093 18717 14105 18720
rect 14139 18748 14151 18751
rect 15933 18751 15991 18757
rect 15933 18748 15945 18751
rect 14139 18720 15945 18748
rect 14139 18717 14151 18720
rect 14093 18711 14151 18717
rect 15933 18717 15945 18720
rect 15979 18717 15991 18751
rect 20714 18748 20720 18760
rect 20627 18720 20720 18748
rect 15933 18711 15991 18717
rect 20714 18708 20720 18720
rect 20772 18748 20778 18760
rect 21726 18748 21732 18760
rect 20772 18720 21732 18748
rect 20772 18708 20778 18720
rect 21726 18708 21732 18720
rect 21784 18708 21790 18760
rect 25685 18751 25743 18757
rect 25685 18717 25697 18751
rect 25731 18748 25743 18751
rect 25958 18748 25964 18760
rect 25731 18720 25964 18748
rect 25731 18717 25743 18720
rect 25685 18711 25743 18717
rect 25958 18708 25964 18720
rect 26016 18708 26022 18760
rect 31113 18751 31171 18757
rect 31113 18717 31125 18751
rect 31159 18717 31171 18751
rect 31113 18711 31171 18717
rect 31380 18751 31438 18757
rect 31380 18717 31392 18751
rect 31426 18748 31438 18751
rect 31754 18748 31760 18760
rect 31426 18720 31760 18748
rect 31426 18717 31438 18720
rect 31380 18711 31438 18717
rect 14360 18683 14418 18689
rect 14360 18649 14372 18683
rect 14406 18680 14418 18683
rect 14734 18680 14740 18692
rect 14406 18652 14740 18680
rect 14406 18649 14418 18652
rect 14360 18643 14418 18649
rect 14734 18640 14740 18652
rect 14792 18640 14798 18692
rect 16178 18683 16236 18689
rect 16178 18680 16190 18683
rect 15488 18652 16190 18680
rect 2958 18612 2964 18624
rect 2919 18584 2964 18612
rect 2958 18572 2964 18584
rect 3016 18572 3022 18624
rect 7742 18612 7748 18624
rect 7703 18584 7748 18612
rect 7742 18572 7748 18584
rect 7800 18572 7806 18624
rect 15488 18621 15516 18652
rect 16178 18649 16190 18652
rect 16224 18649 16236 18683
rect 16178 18643 16236 18649
rect 20984 18683 21042 18689
rect 20984 18649 20996 18683
rect 21030 18680 21042 18683
rect 22278 18680 22284 18692
rect 21030 18652 22284 18680
rect 21030 18649 21042 18652
rect 20984 18643 21042 18649
rect 22278 18640 22284 18652
rect 22336 18640 22342 18692
rect 27433 18683 27491 18689
rect 27433 18649 27445 18683
rect 27479 18680 27491 18683
rect 27614 18680 27620 18692
rect 27479 18652 27620 18680
rect 27479 18649 27491 18652
rect 27433 18643 27491 18649
rect 27614 18640 27620 18652
rect 27672 18640 27678 18692
rect 31128 18680 31156 18711
rect 31754 18708 31760 18720
rect 31812 18708 31818 18760
rect 36078 18748 36084 18760
rect 36039 18720 36084 18748
rect 36078 18708 36084 18720
rect 36136 18708 36142 18760
rect 36348 18751 36406 18757
rect 36348 18717 36360 18751
rect 36394 18748 36406 18751
rect 37826 18748 37832 18760
rect 36394 18720 37832 18748
rect 36394 18717 36406 18720
rect 36348 18711 36406 18717
rect 37826 18708 37832 18720
rect 37884 18708 37890 18760
rect 37921 18751 37979 18757
rect 37921 18717 37933 18751
rect 37967 18717 37979 18751
rect 37921 18711 37979 18717
rect 40120 18751 40178 18757
rect 40120 18717 40132 18751
rect 40166 18748 40178 18751
rect 41414 18748 41420 18760
rect 40166 18720 41420 18748
rect 40166 18717 40178 18720
rect 40120 18711 40178 18717
rect 32766 18680 32772 18692
rect 31128 18652 32772 18680
rect 32766 18640 32772 18652
rect 32824 18640 32830 18692
rect 15473 18615 15531 18621
rect 15473 18581 15485 18615
rect 15519 18581 15531 18615
rect 15473 18575 15531 18581
rect 15562 18572 15568 18624
rect 15620 18612 15626 18624
rect 17313 18615 17371 18621
rect 17313 18612 17325 18615
rect 15620 18584 17325 18612
rect 15620 18572 15626 18584
rect 17313 18581 17325 18584
rect 17359 18581 17371 18615
rect 17313 18575 17371 18581
rect 20714 18572 20720 18624
rect 20772 18612 20778 18624
rect 22097 18615 22155 18621
rect 22097 18612 22109 18615
rect 20772 18584 22109 18612
rect 20772 18572 20778 18584
rect 22097 18581 22109 18584
rect 22143 18581 22155 18615
rect 37458 18612 37464 18624
rect 37419 18584 37464 18612
rect 22097 18575 22155 18581
rect 37458 18572 37464 18584
rect 37516 18572 37522 18624
rect 37936 18612 37964 18711
rect 41414 18708 41420 18720
rect 41472 18708 41478 18760
rect 42337 18751 42395 18757
rect 42337 18717 42349 18751
rect 42383 18748 42395 18751
rect 42426 18748 42432 18760
rect 42383 18720 42432 18748
rect 42383 18717 42395 18720
rect 42337 18711 42395 18717
rect 42426 18708 42432 18720
rect 42484 18708 42490 18760
rect 45002 18708 45008 18760
rect 45060 18748 45066 18760
rect 45097 18751 45155 18757
rect 45097 18748 45109 18751
rect 45060 18720 45109 18748
rect 45060 18708 45066 18720
rect 45097 18717 45109 18720
rect 45143 18717 45155 18751
rect 45097 18711 45155 18717
rect 51905 18751 51963 18757
rect 51905 18717 51917 18751
rect 51951 18748 51963 18751
rect 51994 18748 52000 18760
rect 51951 18720 52000 18748
rect 51951 18717 51963 18720
rect 51905 18711 51963 18717
rect 51994 18708 52000 18720
rect 52052 18708 52058 18760
rect 56686 18748 56692 18760
rect 56647 18720 56692 18748
rect 56686 18708 56692 18720
rect 56744 18708 56750 18760
rect 38188 18683 38246 18689
rect 38188 18649 38200 18683
rect 38234 18680 38246 18683
rect 39666 18680 39672 18692
rect 38234 18652 39672 18680
rect 38234 18649 38246 18652
rect 38188 18643 38246 18649
rect 39666 18640 39672 18652
rect 39724 18640 39730 18692
rect 42604 18683 42662 18689
rect 42604 18649 42616 18683
rect 42650 18680 42662 18683
rect 43806 18680 43812 18692
rect 42650 18652 43812 18680
rect 42650 18649 42662 18652
rect 42604 18643 42662 18649
rect 43806 18640 43812 18652
rect 43864 18640 43870 18692
rect 45364 18683 45422 18689
rect 45364 18649 45376 18683
rect 45410 18680 45422 18683
rect 46382 18680 46388 18692
rect 45410 18652 46388 18680
rect 45410 18649 45422 18652
rect 45364 18643 45422 18649
rect 46382 18640 46388 18652
rect 46440 18640 46446 18692
rect 52172 18683 52230 18689
rect 52172 18649 52184 18683
rect 52218 18680 52230 18683
rect 52638 18680 52644 18692
rect 52218 18652 52644 18680
rect 52218 18649 52230 18652
rect 52172 18643 52230 18649
rect 52638 18640 52644 18652
rect 52696 18640 52702 18692
rect 56956 18683 57014 18689
rect 56956 18649 56968 18683
rect 57002 18680 57014 18683
rect 57238 18680 57244 18692
rect 57002 18652 57244 18680
rect 57002 18649 57014 18652
rect 56956 18643 57014 18649
rect 57238 18640 57244 18652
rect 57296 18640 57302 18692
rect 38286 18612 38292 18624
rect 37936 18584 38292 18612
rect 38286 18572 38292 18584
rect 38344 18572 38350 18624
rect 39298 18612 39304 18624
rect 39259 18584 39304 18612
rect 39298 18572 39304 18584
rect 39356 18572 39362 18624
rect 51810 18572 51816 18624
rect 51868 18612 51874 18624
rect 53285 18615 53343 18621
rect 53285 18612 53297 18615
rect 51868 18584 53297 18612
rect 51868 18572 51874 18584
rect 53285 18581 53297 18584
rect 53331 18581 53343 18615
rect 58066 18612 58072 18624
rect 58027 18584 58072 18612
rect 53285 18575 53343 18581
rect 58066 18572 58072 18584
rect 58124 18572 58130 18624
rect 1104 18522 59340 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 59340 18522
rect 1104 18448 59340 18470
rect 3145 18411 3203 18417
rect 3145 18377 3157 18411
rect 3191 18377 3203 18411
rect 3145 18371 3203 18377
rect 2032 18343 2090 18349
rect 2032 18309 2044 18343
rect 2078 18340 2090 18343
rect 2958 18340 2964 18352
rect 2078 18312 2964 18340
rect 2078 18309 2090 18312
rect 2032 18303 2090 18309
rect 2958 18300 2964 18312
rect 3016 18300 3022 18352
rect 3160 18340 3188 18371
rect 12710 18368 12716 18420
rect 12768 18408 12774 18420
rect 12897 18411 12955 18417
rect 12897 18408 12909 18411
rect 12768 18380 12909 18408
rect 12768 18368 12774 18380
rect 12897 18377 12909 18380
rect 12943 18377 12955 18411
rect 14734 18408 14740 18420
rect 14695 18380 14740 18408
rect 12897 18371 12955 18377
rect 14734 18368 14740 18380
rect 14792 18368 14798 18420
rect 19242 18368 19248 18420
rect 19300 18408 19306 18420
rect 19429 18411 19487 18417
rect 19429 18408 19441 18411
rect 19300 18380 19441 18408
rect 19300 18368 19306 18380
rect 19429 18377 19441 18380
rect 19475 18377 19487 18411
rect 21266 18408 21272 18420
rect 21227 18380 21272 18408
rect 19429 18371 19487 18377
rect 21266 18368 21272 18380
rect 21324 18368 21330 18420
rect 28902 18408 28908 18420
rect 28863 18380 28908 18408
rect 28902 18368 28908 18380
rect 28960 18368 28966 18420
rect 31202 18408 31208 18420
rect 31163 18380 31208 18408
rect 31202 18368 31208 18380
rect 31260 18368 31266 18420
rect 36722 18408 36728 18420
rect 36683 18380 36728 18408
rect 36722 18368 36728 18380
rect 36780 18368 36786 18420
rect 39666 18408 39672 18420
rect 39627 18380 39672 18408
rect 39666 18368 39672 18380
rect 39724 18368 39730 18420
rect 43806 18408 43812 18420
rect 43767 18380 43812 18408
rect 43806 18368 43812 18380
rect 43864 18368 43870 18420
rect 46382 18408 46388 18420
rect 46343 18380 46388 18408
rect 46382 18368 46388 18380
rect 46440 18368 46446 18420
rect 3850 18343 3908 18349
rect 3850 18340 3862 18343
rect 3160 18312 3862 18340
rect 3850 18309 3862 18312
rect 3896 18309 3908 18343
rect 3850 18303 3908 18309
rect 6632 18343 6690 18349
rect 6632 18309 6644 18343
rect 6678 18340 6690 18343
rect 7742 18340 7748 18352
rect 6678 18312 7748 18340
rect 6678 18309 6690 18312
rect 6632 18303 6690 18309
rect 7742 18300 7748 18312
rect 7800 18300 7806 18352
rect 13624 18343 13682 18349
rect 13624 18309 13636 18343
rect 13670 18340 13682 18343
rect 13998 18340 14004 18352
rect 13670 18312 14004 18340
rect 13670 18309 13682 18312
rect 13624 18303 13682 18309
rect 13998 18300 14004 18312
rect 14056 18300 14062 18352
rect 18316 18343 18374 18349
rect 18316 18309 18328 18343
rect 18362 18340 18374 18343
rect 20530 18340 20536 18352
rect 18362 18312 20536 18340
rect 18362 18309 18374 18312
rect 18316 18303 18374 18309
rect 20530 18300 20536 18312
rect 20588 18300 20594 18352
rect 22088 18343 22146 18349
rect 22088 18309 22100 18343
rect 22134 18340 22146 18343
rect 23198 18340 23204 18352
rect 22134 18312 23204 18340
rect 22134 18309 22146 18312
rect 22088 18303 22146 18309
rect 23198 18300 23204 18312
rect 23256 18300 23262 18352
rect 23928 18343 23986 18349
rect 23928 18309 23940 18343
rect 23974 18340 23986 18343
rect 25038 18340 25044 18352
rect 23974 18312 25044 18340
rect 23974 18309 23986 18312
rect 23928 18303 23986 18309
rect 25038 18300 25044 18312
rect 25096 18300 25102 18352
rect 27792 18343 27850 18349
rect 27792 18309 27804 18343
rect 27838 18340 27850 18343
rect 28718 18340 28724 18352
rect 27838 18312 28724 18340
rect 27838 18309 27850 18312
rect 27792 18303 27850 18309
rect 28718 18300 28724 18312
rect 28776 18300 28782 18352
rect 30092 18343 30150 18349
rect 30092 18309 30104 18343
rect 30138 18340 30150 18343
rect 33502 18340 33508 18352
rect 30138 18312 33508 18340
rect 30138 18309 30150 18312
rect 30092 18303 30150 18309
rect 33502 18300 33508 18312
rect 33560 18300 33566 18352
rect 33772 18343 33830 18349
rect 33772 18309 33784 18343
rect 33818 18340 33830 18343
rect 34514 18340 34520 18352
rect 33818 18312 34520 18340
rect 33818 18309 33830 18312
rect 33772 18303 33830 18309
rect 34514 18300 34520 18312
rect 34572 18300 34578 18352
rect 36078 18340 36084 18352
rect 35360 18312 36084 18340
rect 1578 18232 1584 18284
rect 1636 18272 1642 18284
rect 1765 18275 1823 18281
rect 1765 18272 1777 18275
rect 1636 18244 1777 18272
rect 1636 18232 1642 18244
rect 1765 18241 1777 18244
rect 1811 18241 1823 18275
rect 1765 18235 1823 18241
rect 3605 18275 3663 18281
rect 3605 18241 3617 18275
rect 3651 18272 3663 18275
rect 4614 18272 4620 18284
rect 3651 18244 4620 18272
rect 3651 18241 3663 18244
rect 3605 18235 3663 18241
rect 4614 18232 4620 18244
rect 4672 18272 4678 18284
rect 6362 18272 6368 18284
rect 4672 18244 6368 18272
rect 4672 18232 4678 18244
rect 6362 18232 6368 18244
rect 6420 18272 6426 18284
rect 8205 18275 8263 18281
rect 8205 18272 8217 18275
rect 6420 18244 8217 18272
rect 6420 18232 6426 18244
rect 8205 18241 8217 18244
rect 8251 18241 8263 18275
rect 8205 18235 8263 18241
rect 8294 18232 8300 18284
rect 8352 18232 8358 18284
rect 8472 18275 8530 18281
rect 8472 18241 8484 18275
rect 8518 18272 8530 18275
rect 9398 18272 9404 18284
rect 8518 18244 9404 18272
rect 8518 18241 8530 18244
rect 8472 18235 8530 18241
rect 9398 18232 9404 18244
rect 9456 18232 9462 18284
rect 11517 18275 11575 18281
rect 11517 18241 11529 18275
rect 11563 18272 11575 18275
rect 11606 18272 11612 18284
rect 11563 18244 11612 18272
rect 11563 18241 11575 18244
rect 11517 18235 11575 18241
rect 11606 18232 11612 18244
rect 11664 18232 11670 18284
rect 11784 18275 11842 18281
rect 11784 18241 11796 18275
rect 11830 18272 11842 18275
rect 12894 18272 12900 18284
rect 11830 18244 12900 18272
rect 11830 18241 11842 18244
rect 11784 18235 11842 18241
rect 12894 18232 12900 18244
rect 12952 18232 12958 18284
rect 13357 18275 13415 18281
rect 13357 18241 13369 18275
rect 13403 18272 13415 18275
rect 14090 18272 14096 18284
rect 13403 18244 14096 18272
rect 13403 18241 13415 18244
rect 13357 18235 13415 18241
rect 14090 18232 14096 18244
rect 14148 18232 14154 18284
rect 20156 18275 20214 18281
rect 20156 18241 20168 18275
rect 20202 18272 20214 18275
rect 21266 18272 21272 18284
rect 20202 18244 21272 18272
rect 20202 18241 20214 18244
rect 20156 18235 20214 18241
rect 21266 18232 21272 18244
rect 21324 18232 21330 18284
rect 21726 18232 21732 18284
rect 21784 18272 21790 18284
rect 21821 18275 21879 18281
rect 21821 18272 21833 18275
rect 21784 18244 21833 18272
rect 21784 18232 21790 18244
rect 21821 18241 21833 18244
rect 21867 18241 21879 18275
rect 23658 18272 23664 18284
rect 23619 18244 23664 18272
rect 21821 18235 21879 18241
rect 23658 18232 23664 18244
rect 23716 18232 23722 18284
rect 27525 18275 27583 18281
rect 27525 18241 27537 18275
rect 27571 18272 27583 18275
rect 27614 18272 27620 18284
rect 27571 18244 27620 18272
rect 27571 18241 27583 18244
rect 27525 18235 27583 18241
rect 27614 18232 27620 18244
rect 27672 18232 27678 18284
rect 29825 18275 29883 18281
rect 29825 18241 29837 18275
rect 29871 18272 29883 18275
rect 29914 18272 29920 18284
rect 29871 18244 29920 18272
rect 29871 18241 29883 18244
rect 29825 18235 29883 18241
rect 29914 18232 29920 18244
rect 29972 18232 29978 18284
rect 35360 18281 35388 18312
rect 36078 18300 36084 18312
rect 36136 18300 36142 18352
rect 38556 18343 38614 18349
rect 38556 18309 38568 18343
rect 38602 18340 38614 18343
rect 38654 18340 38660 18352
rect 38602 18312 38660 18340
rect 38602 18309 38614 18312
rect 38556 18303 38614 18309
rect 38654 18300 38660 18312
rect 38712 18300 38718 18352
rect 40126 18340 40132 18352
rect 40087 18312 40132 18340
rect 40126 18300 40132 18312
rect 40184 18300 40190 18352
rect 51258 18340 51264 18352
rect 50724 18312 51264 18340
rect 35345 18275 35403 18281
rect 35345 18272 35357 18275
rect 33520 18244 35357 18272
rect 8312 18204 8340 18232
rect 7760 18176 8340 18204
rect 7760 18145 7788 18176
rect 17310 18164 17316 18216
rect 17368 18204 17374 18216
rect 18049 18207 18107 18213
rect 18049 18204 18061 18207
rect 17368 18176 18061 18204
rect 17368 18164 17374 18176
rect 18049 18173 18061 18176
rect 18095 18173 18107 18207
rect 18049 18167 18107 18173
rect 19889 18207 19947 18213
rect 19889 18173 19901 18207
rect 19935 18173 19947 18207
rect 19889 18167 19947 18173
rect 7745 18139 7803 18145
rect 7745 18105 7757 18139
rect 7791 18105 7803 18139
rect 7745 18099 7803 18105
rect 4982 18068 4988 18080
rect 4943 18040 4988 18068
rect 4982 18028 4988 18040
rect 5040 18028 5046 18080
rect 9582 18068 9588 18080
rect 9543 18040 9588 18068
rect 9582 18028 9588 18040
rect 9640 18028 9646 18080
rect 19904 18068 19932 18167
rect 32766 18164 32772 18216
rect 32824 18204 32830 18216
rect 33520 18213 33548 18244
rect 35345 18241 35357 18244
rect 35391 18241 35403 18275
rect 35345 18235 35403 18241
rect 35612 18275 35670 18281
rect 35612 18241 35624 18275
rect 35658 18272 35670 18275
rect 37090 18272 37096 18284
rect 35658 18244 37096 18272
rect 35658 18241 35670 18244
rect 35612 18235 35670 18241
rect 37090 18232 37096 18244
rect 37148 18232 37154 18284
rect 38286 18272 38292 18284
rect 38247 18244 38292 18272
rect 38286 18232 38292 18244
rect 38344 18232 38350 18284
rect 41506 18232 41512 18284
rect 41564 18272 41570 18284
rect 41877 18275 41935 18281
rect 41877 18272 41889 18275
rect 41564 18244 41889 18272
rect 41564 18232 41570 18244
rect 41877 18241 41889 18244
rect 41923 18272 41935 18275
rect 42429 18275 42487 18281
rect 42429 18272 42441 18275
rect 41923 18244 42441 18272
rect 41923 18241 41935 18244
rect 41877 18235 41935 18241
rect 42429 18241 42441 18244
rect 42475 18241 42487 18275
rect 42429 18235 42487 18241
rect 42696 18275 42754 18281
rect 42696 18241 42708 18275
rect 42742 18272 42754 18275
rect 43530 18272 43536 18284
rect 42742 18244 43536 18272
rect 42742 18241 42754 18244
rect 42696 18235 42754 18241
rect 43530 18232 43536 18244
rect 43588 18232 43594 18284
rect 45005 18275 45063 18281
rect 45005 18241 45017 18275
rect 45051 18272 45063 18275
rect 45094 18272 45100 18284
rect 45051 18244 45100 18272
rect 45051 18241 45063 18244
rect 45005 18235 45063 18241
rect 45094 18232 45100 18244
rect 45152 18232 45158 18284
rect 45272 18275 45330 18281
rect 45272 18241 45284 18275
rect 45318 18272 45330 18275
rect 46382 18272 46388 18284
rect 45318 18244 46388 18272
rect 45318 18241 45330 18244
rect 45272 18235 45330 18241
rect 46382 18232 46388 18244
rect 46440 18232 46446 18284
rect 50724 18281 50752 18312
rect 51258 18300 51264 18312
rect 51316 18340 51322 18352
rect 51994 18340 52000 18352
rect 51316 18312 52000 18340
rect 51316 18300 51322 18312
rect 51994 18300 52000 18312
rect 52052 18300 52058 18352
rect 56220 18343 56278 18349
rect 56220 18309 56232 18343
rect 56266 18340 56278 18343
rect 58066 18340 58072 18352
rect 56266 18312 58072 18340
rect 56266 18309 56278 18312
rect 56220 18303 56278 18309
rect 58066 18300 58072 18312
rect 58124 18300 58130 18352
rect 50709 18275 50767 18281
rect 50709 18241 50721 18275
rect 50755 18241 50767 18275
rect 50709 18235 50767 18241
rect 50976 18275 51034 18281
rect 50976 18241 50988 18275
rect 51022 18272 51034 18275
rect 52178 18272 52184 18284
rect 51022 18244 52184 18272
rect 51022 18241 51034 18244
rect 50976 18235 51034 18241
rect 52178 18232 52184 18244
rect 52236 18232 52242 18284
rect 54196 18275 54254 18281
rect 54196 18241 54208 18275
rect 54242 18272 54254 18275
rect 54754 18272 54760 18284
rect 54242 18244 54760 18272
rect 54242 18241 54254 18244
rect 54196 18235 54254 18241
rect 54754 18232 54760 18244
rect 54812 18232 54818 18284
rect 55953 18275 56011 18281
rect 55953 18241 55965 18275
rect 55999 18272 56011 18275
rect 56686 18272 56692 18284
rect 55999 18244 56692 18272
rect 55999 18241 56011 18244
rect 55953 18235 56011 18241
rect 56686 18232 56692 18244
rect 56744 18232 56750 18284
rect 33505 18207 33563 18213
rect 33505 18204 33517 18207
rect 32824 18176 33517 18204
rect 32824 18164 32830 18176
rect 33505 18173 33517 18176
rect 33551 18173 33563 18207
rect 33505 18167 33563 18173
rect 53834 18164 53840 18216
rect 53892 18204 53898 18216
rect 53929 18207 53987 18213
rect 53929 18204 53941 18207
rect 53892 18176 53941 18204
rect 53892 18164 53898 18176
rect 53929 18173 53941 18176
rect 53975 18173 53987 18207
rect 53929 18167 53987 18173
rect 23201 18139 23259 18145
rect 23201 18105 23213 18139
rect 23247 18136 23259 18139
rect 23474 18136 23480 18148
rect 23247 18108 23480 18136
rect 23247 18105 23259 18108
rect 23201 18099 23259 18105
rect 23474 18096 23480 18108
rect 23532 18096 23538 18148
rect 20898 18068 20904 18080
rect 19904 18040 20904 18068
rect 20898 18028 20904 18040
rect 20956 18028 20962 18080
rect 25041 18071 25099 18077
rect 25041 18037 25053 18071
rect 25087 18068 25099 18071
rect 25222 18068 25228 18080
rect 25087 18040 25228 18068
rect 25087 18037 25099 18040
rect 25041 18031 25099 18037
rect 25222 18028 25228 18040
rect 25280 18028 25286 18080
rect 34885 18071 34943 18077
rect 34885 18037 34897 18071
rect 34931 18068 34943 18071
rect 36354 18068 36360 18080
rect 34931 18040 36360 18068
rect 34931 18037 34943 18040
rect 34885 18031 34943 18037
rect 36354 18028 36360 18040
rect 36412 18028 36418 18080
rect 50614 18028 50620 18080
rect 50672 18068 50678 18080
rect 52089 18071 52147 18077
rect 52089 18068 52101 18071
rect 50672 18040 52101 18068
rect 50672 18028 50678 18040
rect 52089 18037 52101 18040
rect 52135 18037 52147 18071
rect 52089 18031 52147 18037
rect 54294 18028 54300 18080
rect 54352 18068 54358 18080
rect 55309 18071 55367 18077
rect 55309 18068 55321 18071
rect 54352 18040 55321 18068
rect 54352 18028 54358 18040
rect 55309 18037 55321 18040
rect 55355 18037 55367 18071
rect 55309 18031 55367 18037
rect 55858 18028 55864 18080
rect 55916 18068 55922 18080
rect 57333 18071 57391 18077
rect 57333 18068 57345 18071
rect 55916 18040 57345 18068
rect 55916 18028 55922 18040
rect 57333 18037 57345 18040
rect 57379 18037 57391 18071
rect 57333 18031 57391 18037
rect 1104 17978 59340 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 59340 17978
rect 1104 17904 59340 17926
rect 22278 17864 22284 17876
rect 22239 17836 22284 17864
rect 22278 17824 22284 17836
rect 22336 17824 22342 17876
rect 37090 17824 37096 17876
rect 37148 17864 37154 17876
rect 37461 17867 37519 17873
rect 37461 17864 37473 17867
rect 37148 17836 37473 17864
rect 37148 17824 37154 17836
rect 37461 17833 37473 17836
rect 37507 17833 37519 17867
rect 38286 17864 38292 17876
rect 37461 17827 37519 17833
rect 37936 17836 38292 17864
rect 1578 17688 1584 17740
rect 1636 17728 1642 17740
rect 2498 17728 2504 17740
rect 1636 17700 2504 17728
rect 1636 17688 1642 17700
rect 2498 17688 2504 17700
rect 2556 17728 2562 17740
rect 3789 17731 3847 17737
rect 3789 17728 3801 17731
rect 2556 17700 3801 17728
rect 2556 17688 2562 17700
rect 3789 17697 3801 17700
rect 3835 17697 3847 17731
rect 14090 17728 14096 17740
rect 14051 17700 14096 17728
rect 3789 17691 3847 17697
rect 14090 17688 14096 17700
rect 14148 17688 14154 17740
rect 29914 17688 29920 17740
rect 29972 17728 29978 17740
rect 30929 17731 30987 17737
rect 30929 17728 30941 17731
rect 29972 17700 30941 17728
rect 29972 17688 29978 17700
rect 30929 17697 30941 17700
rect 30975 17697 30987 17731
rect 32766 17728 32772 17740
rect 32727 17700 32772 17728
rect 30929 17691 30987 17697
rect 32766 17688 32772 17700
rect 32824 17688 32830 17740
rect 37366 17688 37372 17740
rect 37424 17728 37430 17740
rect 37936 17737 37964 17836
rect 38286 17824 38292 17836
rect 38344 17824 38350 17876
rect 39114 17824 39120 17876
rect 39172 17864 39178 17876
rect 39301 17867 39359 17873
rect 39301 17864 39313 17867
rect 39172 17836 39313 17864
rect 39172 17824 39178 17836
rect 39301 17833 39313 17836
rect 39347 17833 39359 17867
rect 42426 17864 42432 17876
rect 39301 17827 39359 17833
rect 42168 17836 42432 17864
rect 42168 17737 42196 17836
rect 42426 17824 42432 17836
rect 42484 17824 42490 17876
rect 43530 17864 43536 17876
rect 43491 17836 43536 17864
rect 43530 17824 43536 17836
rect 43588 17824 43594 17876
rect 46382 17864 46388 17876
rect 46343 17836 46388 17864
rect 46382 17824 46388 17836
rect 46440 17824 46446 17876
rect 52638 17864 52644 17876
rect 52599 17836 52644 17864
rect 52638 17824 52644 17836
rect 52696 17824 52702 17876
rect 53834 17864 53840 17876
rect 53116 17836 53840 17864
rect 37921 17731 37979 17737
rect 37921 17728 37933 17731
rect 37424 17700 37933 17728
rect 37424 17688 37430 17700
rect 37921 17697 37933 17700
rect 37967 17697 37979 17731
rect 37921 17691 37979 17697
rect 42153 17731 42211 17737
rect 42153 17697 42165 17731
rect 42199 17697 42211 17731
rect 45002 17728 45008 17740
rect 44963 17700 45008 17728
rect 42153 17691 42211 17697
rect 45002 17688 45008 17700
rect 45060 17688 45066 17740
rect 47210 17688 47216 17740
rect 47268 17728 47274 17740
rect 47673 17731 47731 17737
rect 47673 17728 47685 17731
rect 47268 17700 47685 17728
rect 47268 17688 47274 17700
rect 47673 17697 47685 17700
rect 47719 17697 47731 17731
rect 51258 17728 51264 17740
rect 51219 17700 51264 17728
rect 47673 17691 47731 17697
rect 51258 17688 51264 17700
rect 51316 17688 51322 17740
rect 4522 17620 4528 17672
rect 4580 17660 4586 17672
rect 5442 17660 5448 17672
rect 4580 17632 5448 17660
rect 4580 17620 4586 17632
rect 5442 17620 5448 17632
rect 5500 17660 5506 17672
rect 6273 17663 6331 17669
rect 6273 17660 6285 17663
rect 5500 17632 6285 17660
rect 5500 17620 5506 17632
rect 6273 17629 6285 17632
rect 6319 17629 6331 17663
rect 8938 17660 8944 17672
rect 8851 17632 8944 17660
rect 6273 17623 6331 17629
rect 8938 17620 8944 17632
rect 8996 17660 9002 17672
rect 10781 17663 10839 17669
rect 10781 17660 10793 17663
rect 8996 17632 10793 17660
rect 8996 17620 9002 17632
rect 10781 17629 10793 17632
rect 10827 17660 10839 17663
rect 11606 17660 11612 17672
rect 10827 17632 11612 17660
rect 10827 17629 10839 17632
rect 10781 17623 10839 17629
rect 11606 17620 11612 17632
rect 11664 17620 11670 17672
rect 14360 17663 14418 17669
rect 14360 17629 14372 17663
rect 14406 17660 14418 17663
rect 15562 17660 15568 17672
rect 14406 17632 15568 17660
rect 14406 17629 14418 17632
rect 14360 17623 14418 17629
rect 15562 17620 15568 17632
rect 15620 17620 15626 17672
rect 15933 17663 15991 17669
rect 15933 17629 15945 17663
rect 15979 17660 15991 17663
rect 17310 17660 17316 17672
rect 15979 17632 17316 17660
rect 15979 17629 15991 17632
rect 15933 17623 15991 17629
rect 17310 17620 17316 17632
rect 17368 17620 17374 17672
rect 20898 17660 20904 17672
rect 20811 17632 20904 17660
rect 20898 17620 20904 17632
rect 20956 17660 20962 17672
rect 21726 17660 21732 17672
rect 20956 17632 21732 17660
rect 20956 17620 20962 17632
rect 21726 17620 21732 17632
rect 21784 17620 21790 17672
rect 24394 17620 24400 17672
rect 24452 17660 24458 17672
rect 25133 17663 25191 17669
rect 25133 17660 25145 17663
rect 24452 17632 25145 17660
rect 24452 17620 24458 17632
rect 25133 17629 25145 17632
rect 25179 17629 25191 17663
rect 25133 17623 25191 17629
rect 3878 17552 3884 17604
rect 3936 17592 3942 17604
rect 4034 17595 4092 17601
rect 4034 17592 4046 17595
rect 3936 17564 4046 17592
rect 3936 17552 3942 17564
rect 4034 17561 4046 17564
rect 4080 17561 4092 17595
rect 4034 17555 4092 17561
rect 6540 17595 6598 17601
rect 6540 17561 6552 17595
rect 6586 17592 6598 17595
rect 7742 17592 7748 17604
rect 6586 17564 7748 17592
rect 6586 17561 6598 17564
rect 6540 17555 6598 17561
rect 7742 17552 7748 17564
rect 7800 17552 7806 17604
rect 9208 17595 9266 17601
rect 9208 17561 9220 17595
rect 9254 17592 9266 17595
rect 10226 17592 10232 17604
rect 9254 17564 10232 17592
rect 9254 17561 9266 17564
rect 9208 17555 9266 17561
rect 10226 17552 10232 17564
rect 10284 17552 10290 17604
rect 11026 17595 11084 17601
rect 11026 17592 11038 17595
rect 10336 17564 11038 17592
rect 4614 17484 4620 17536
rect 4672 17524 4678 17536
rect 5169 17527 5227 17533
rect 5169 17524 5181 17527
rect 4672 17496 5181 17524
rect 4672 17484 4678 17496
rect 5169 17493 5181 17496
rect 5215 17493 5227 17527
rect 5169 17487 5227 17493
rect 7653 17527 7711 17533
rect 7653 17493 7665 17527
rect 7699 17524 7711 17527
rect 8386 17524 8392 17536
rect 7699 17496 8392 17524
rect 7699 17493 7711 17496
rect 7653 17487 7711 17493
rect 8386 17484 8392 17496
rect 8444 17484 8450 17536
rect 10336 17533 10364 17564
rect 11026 17561 11038 17564
rect 11072 17561 11084 17595
rect 11026 17555 11084 17561
rect 15838 17552 15844 17604
rect 15896 17592 15902 17604
rect 16178 17595 16236 17601
rect 16178 17592 16190 17595
rect 15896 17564 16190 17592
rect 15896 17552 15902 17564
rect 16178 17561 16190 17564
rect 16224 17561 16236 17595
rect 16178 17555 16236 17561
rect 21168 17595 21226 17601
rect 21168 17561 21180 17595
rect 21214 17592 21226 17595
rect 23198 17592 23204 17604
rect 21214 17564 23204 17592
rect 21214 17561 21226 17564
rect 21168 17555 21226 17561
rect 23198 17552 23204 17564
rect 23256 17552 23262 17604
rect 25148 17592 25176 17623
rect 25222 17620 25228 17672
rect 25280 17660 25286 17672
rect 25389 17663 25447 17669
rect 25389 17660 25401 17663
rect 25280 17632 25401 17660
rect 25280 17620 25286 17632
rect 25389 17629 25401 17632
rect 25435 17629 25447 17663
rect 27614 17660 27620 17672
rect 25389 17623 25447 17629
rect 26206 17632 27620 17660
rect 26206 17592 26234 17632
rect 27614 17620 27620 17632
rect 27672 17620 27678 17672
rect 36081 17663 36139 17669
rect 36081 17629 36093 17663
rect 36127 17660 36139 17663
rect 37384 17660 37412 17688
rect 36127 17632 37412 17660
rect 38188 17663 38246 17669
rect 36127 17629 36139 17632
rect 36081 17623 36139 17629
rect 38188 17629 38200 17663
rect 38234 17660 38246 17663
rect 39298 17660 39304 17672
rect 38234 17632 39304 17660
rect 38234 17629 38246 17632
rect 38188 17623 38246 17629
rect 39298 17620 39304 17632
rect 39356 17620 39362 17672
rect 51276 17660 51304 17688
rect 53116 17669 53144 17836
rect 53834 17824 53840 17836
rect 53892 17824 53898 17876
rect 53101 17663 53159 17669
rect 53101 17660 53113 17663
rect 51276 17632 53113 17660
rect 53101 17629 53113 17632
rect 53147 17629 53159 17663
rect 53101 17623 53159 17629
rect 53368 17663 53426 17669
rect 53368 17629 53380 17663
rect 53414 17660 53426 17663
rect 54294 17660 54300 17672
rect 53414 17632 54300 17660
rect 53414 17629 53426 17632
rect 53368 17623 53426 17629
rect 54294 17620 54300 17632
rect 54352 17620 54358 17672
rect 55950 17620 55956 17672
rect 56008 17660 56014 17672
rect 56781 17663 56839 17669
rect 56781 17660 56793 17663
rect 56008 17632 56793 17660
rect 56008 17620 56014 17632
rect 56781 17629 56793 17632
rect 56827 17629 56839 17663
rect 56781 17623 56839 17629
rect 25148 17564 26234 17592
rect 27884 17595 27942 17601
rect 27884 17561 27896 17595
rect 27930 17592 27942 17595
rect 29730 17592 29736 17604
rect 27930 17564 29736 17592
rect 27930 17561 27942 17564
rect 27884 17555 27942 17561
rect 29730 17552 29736 17564
rect 29788 17552 29794 17604
rect 31196 17595 31254 17601
rect 31196 17561 31208 17595
rect 31242 17592 31254 17595
rect 31570 17592 31576 17604
rect 31242 17564 31576 17592
rect 31242 17561 31254 17564
rect 31196 17555 31254 17561
rect 31570 17552 31576 17564
rect 31628 17552 31634 17604
rect 33036 17595 33094 17601
rect 33036 17561 33048 17595
rect 33082 17592 33094 17595
rect 35342 17592 35348 17604
rect 33082 17564 35348 17592
rect 33082 17561 33094 17564
rect 33036 17555 33094 17561
rect 35342 17552 35348 17564
rect 35400 17552 35406 17604
rect 36348 17595 36406 17601
rect 36348 17561 36360 17595
rect 36394 17592 36406 17595
rect 38838 17592 38844 17604
rect 36394 17564 38844 17592
rect 36394 17561 36406 17564
rect 36348 17555 36406 17561
rect 38838 17552 38844 17564
rect 38896 17552 38902 17604
rect 42420 17595 42478 17601
rect 42420 17561 42432 17595
rect 42466 17592 42478 17595
rect 43806 17592 43812 17604
rect 42466 17564 43812 17592
rect 42466 17561 42478 17564
rect 42420 17555 42478 17561
rect 43806 17552 43812 17564
rect 43864 17552 43870 17604
rect 45272 17595 45330 17601
rect 45272 17561 45284 17595
rect 45318 17592 45330 17595
rect 46290 17592 46296 17604
rect 45318 17564 46296 17592
rect 45318 17561 45330 17564
rect 45272 17555 45330 17561
rect 46290 17552 46296 17564
rect 46348 17552 46354 17604
rect 47940 17595 47998 17601
rect 47940 17561 47952 17595
rect 47986 17592 47998 17595
rect 48774 17592 48780 17604
rect 47986 17564 48780 17592
rect 47986 17561 47998 17564
rect 47940 17555 47998 17561
rect 48774 17552 48780 17564
rect 48832 17552 48838 17604
rect 51528 17595 51586 17601
rect 51528 17561 51540 17595
rect 51574 17592 51586 17595
rect 57048 17595 57106 17601
rect 51574 17564 54524 17592
rect 51574 17561 51586 17564
rect 51528 17555 51586 17561
rect 10321 17527 10379 17533
rect 10321 17493 10333 17527
rect 10367 17493 10379 17527
rect 10321 17487 10379 17493
rect 11330 17484 11336 17536
rect 11388 17524 11394 17536
rect 12161 17527 12219 17533
rect 12161 17524 12173 17527
rect 11388 17496 12173 17524
rect 11388 17484 11394 17496
rect 12161 17493 12173 17496
rect 12207 17493 12219 17527
rect 15470 17524 15476 17536
rect 15431 17496 15476 17524
rect 12161 17487 12219 17493
rect 15470 17484 15476 17496
rect 15528 17484 15534 17536
rect 15746 17484 15752 17536
rect 15804 17524 15810 17536
rect 17313 17527 17371 17533
rect 17313 17524 17325 17527
rect 15804 17496 17325 17524
rect 15804 17484 15810 17496
rect 17313 17493 17325 17496
rect 17359 17493 17371 17527
rect 26510 17524 26516 17536
rect 26471 17496 26516 17524
rect 17313 17487 17371 17493
rect 26510 17484 26516 17496
rect 26568 17484 26574 17536
rect 28994 17524 29000 17536
rect 28955 17496 29000 17524
rect 28994 17484 29000 17496
rect 29052 17484 29058 17536
rect 30466 17484 30472 17536
rect 30524 17524 30530 17536
rect 32309 17527 32367 17533
rect 32309 17524 32321 17527
rect 30524 17496 32321 17524
rect 30524 17484 30530 17496
rect 32309 17493 32321 17496
rect 32355 17493 32367 17527
rect 32309 17487 32367 17493
rect 34149 17527 34207 17533
rect 34149 17493 34161 17527
rect 34195 17524 34207 17527
rect 34790 17524 34796 17536
rect 34195 17496 34796 17524
rect 34195 17493 34207 17496
rect 34149 17487 34207 17493
rect 34790 17484 34796 17496
rect 34848 17484 34854 17536
rect 49050 17524 49056 17536
rect 49011 17496 49056 17524
rect 49050 17484 49056 17496
rect 49108 17484 49114 17536
rect 54496 17533 54524 17564
rect 57048 17561 57060 17595
rect 57094 17592 57106 17595
rect 57330 17592 57336 17604
rect 57094 17564 57336 17592
rect 57094 17561 57106 17564
rect 57048 17555 57106 17561
rect 57330 17552 57336 17564
rect 57388 17552 57394 17604
rect 54481 17527 54539 17533
rect 54481 17493 54493 17527
rect 54527 17493 54539 17527
rect 58158 17524 58164 17536
rect 58119 17496 58164 17524
rect 54481 17487 54539 17493
rect 58158 17484 58164 17496
rect 58216 17484 58222 17536
rect 1104 17434 59340 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 59340 17434
rect 1104 17360 59340 17382
rect 3878 17320 3884 17332
rect 3839 17292 3884 17320
rect 3878 17280 3884 17292
rect 3936 17280 3942 17332
rect 7742 17320 7748 17332
rect 7703 17292 7748 17320
rect 7742 17280 7748 17292
rect 7800 17280 7806 17332
rect 9398 17280 9404 17332
rect 9456 17320 9462 17332
rect 9585 17323 9643 17329
rect 9585 17320 9597 17323
rect 9456 17292 9597 17320
rect 9456 17280 9462 17292
rect 9585 17289 9597 17292
rect 9631 17289 9643 17323
rect 12894 17320 12900 17332
rect 12855 17292 12900 17320
rect 9585 17283 9643 17289
rect 12894 17280 12900 17292
rect 12952 17280 12958 17332
rect 21266 17320 21272 17332
rect 21227 17292 21272 17320
rect 21266 17280 21272 17292
rect 21324 17280 21330 17332
rect 23198 17320 23204 17332
rect 23159 17292 23204 17320
rect 23198 17280 23204 17292
rect 23256 17280 23262 17332
rect 28994 17280 29000 17332
rect 29052 17320 29058 17332
rect 35342 17320 35348 17332
rect 29052 17292 32413 17320
rect 35303 17292 35348 17320
rect 29052 17280 29058 17292
rect 2768 17255 2826 17261
rect 2768 17221 2780 17255
rect 2814 17252 2826 17255
rect 4982 17252 4988 17264
rect 2814 17224 4988 17252
rect 2814 17221 2826 17224
rect 2768 17215 2826 17221
rect 4982 17212 4988 17224
rect 5040 17212 5046 17264
rect 8938 17252 8944 17264
rect 8220 17224 8944 17252
rect 2498 17184 2504 17196
rect 2459 17156 2504 17184
rect 2498 17144 2504 17156
rect 2556 17144 2562 17196
rect 4341 17187 4399 17193
rect 4341 17153 4353 17187
rect 4387 17184 4399 17187
rect 4430 17184 4436 17196
rect 4387 17156 4436 17184
rect 4387 17153 4399 17156
rect 4341 17147 4399 17153
rect 4430 17144 4436 17156
rect 4488 17144 4494 17196
rect 4608 17187 4666 17193
rect 4608 17153 4620 17187
rect 4654 17184 4666 17187
rect 5166 17184 5172 17196
rect 4654 17156 5172 17184
rect 4654 17153 4666 17156
rect 4608 17147 4666 17153
rect 5166 17144 5172 17156
rect 5224 17144 5230 17196
rect 5442 17144 5448 17196
rect 5500 17184 5506 17196
rect 6365 17187 6423 17193
rect 6365 17184 6377 17187
rect 5500 17156 6377 17184
rect 5500 17144 5506 17156
rect 6365 17153 6377 17156
rect 6411 17153 6423 17187
rect 6365 17147 6423 17153
rect 6632 17187 6690 17193
rect 6632 17153 6644 17187
rect 6678 17184 6690 17187
rect 7006 17184 7012 17196
rect 6678 17156 7012 17184
rect 6678 17153 6690 17156
rect 6632 17147 6690 17153
rect 7006 17144 7012 17156
rect 7064 17144 7070 17196
rect 8220 17193 8248 17224
rect 8938 17212 8944 17224
rect 8996 17212 9002 17264
rect 14360 17255 14418 17261
rect 14360 17221 14372 17255
rect 14406 17252 14418 17255
rect 15470 17252 15476 17264
rect 14406 17224 15476 17252
rect 14406 17221 14418 17224
rect 14360 17215 14418 17221
rect 15470 17212 15476 17224
rect 15528 17212 15534 17264
rect 20156 17255 20214 17261
rect 20156 17221 20168 17255
rect 20202 17252 20214 17255
rect 20714 17252 20720 17264
rect 20202 17224 20720 17252
rect 20202 17221 20214 17224
rect 20156 17215 20214 17221
rect 20714 17212 20720 17224
rect 20772 17212 20778 17264
rect 24664 17255 24722 17261
rect 24664 17221 24676 17255
rect 24710 17252 24722 17255
rect 26510 17252 26516 17264
rect 24710 17224 26516 17252
rect 24710 17221 24722 17224
rect 24664 17215 24722 17221
rect 26510 17212 26516 17224
rect 26568 17212 26574 17264
rect 30466 17261 30472 17264
rect 30460 17252 30472 17261
rect 30427 17224 30472 17252
rect 30460 17215 30472 17224
rect 30466 17212 30472 17215
rect 30524 17212 30530 17264
rect 32385 17261 32413 17292
rect 35342 17280 35348 17292
rect 35400 17280 35406 17332
rect 36998 17280 37004 17332
rect 37056 17320 37062 17332
rect 38746 17320 38752 17332
rect 37056 17292 37780 17320
rect 38707 17292 38752 17320
rect 37056 17280 37062 17292
rect 32370 17255 32428 17261
rect 32370 17221 32382 17255
rect 32416 17221 32428 17255
rect 32370 17215 32428 17221
rect 32766 17212 32772 17264
rect 32824 17252 32830 17264
rect 32824 17224 34008 17252
rect 32824 17212 32830 17224
rect 8205 17187 8263 17193
rect 8205 17153 8217 17187
rect 8251 17153 8263 17187
rect 8205 17147 8263 17153
rect 8472 17187 8530 17193
rect 8472 17153 8484 17187
rect 8518 17184 8530 17187
rect 9398 17184 9404 17196
rect 8518 17156 9404 17184
rect 8518 17153 8530 17156
rect 8472 17147 8530 17153
rect 9398 17144 9404 17156
rect 9456 17144 9462 17196
rect 11517 17187 11575 17193
rect 11517 17153 11529 17187
rect 11563 17184 11575 17187
rect 11606 17184 11612 17196
rect 11563 17156 11612 17184
rect 11563 17153 11575 17156
rect 11517 17147 11575 17153
rect 11606 17144 11612 17156
rect 11664 17144 11670 17196
rect 11784 17187 11842 17193
rect 11784 17153 11796 17187
rect 11830 17184 11842 17187
rect 12158 17184 12164 17196
rect 11830 17156 12164 17184
rect 11830 17153 11842 17156
rect 11784 17147 11842 17153
rect 12158 17144 12164 17156
rect 12216 17144 12222 17196
rect 14090 17184 14096 17196
rect 14051 17156 14096 17184
rect 14090 17144 14096 17156
rect 14148 17144 14154 17196
rect 17221 17187 17279 17193
rect 17221 17153 17233 17187
rect 17267 17184 17279 17187
rect 17310 17184 17316 17196
rect 17267 17156 17316 17184
rect 17267 17153 17279 17156
rect 17221 17147 17279 17153
rect 17310 17144 17316 17156
rect 17368 17144 17374 17196
rect 17488 17187 17546 17193
rect 17488 17153 17500 17187
rect 17534 17184 17546 17187
rect 18506 17184 18512 17196
rect 17534 17156 18512 17184
rect 17534 17153 17546 17156
rect 17488 17147 17546 17153
rect 18506 17144 18512 17156
rect 18564 17144 18570 17196
rect 19889 17187 19947 17193
rect 19889 17153 19901 17187
rect 19935 17184 19947 17187
rect 20898 17184 20904 17196
rect 19935 17156 20904 17184
rect 19935 17153 19947 17156
rect 19889 17147 19947 17153
rect 20898 17144 20904 17156
rect 20956 17144 20962 17196
rect 21818 17184 21824 17196
rect 21779 17156 21824 17184
rect 21818 17144 21824 17156
rect 21876 17144 21882 17196
rect 22088 17187 22146 17193
rect 22088 17153 22100 17187
rect 22134 17184 22146 17187
rect 23198 17184 23204 17196
rect 22134 17156 23204 17184
rect 22134 17153 22146 17156
rect 22088 17147 22146 17153
rect 23198 17144 23204 17156
rect 23256 17144 23262 17196
rect 23658 17144 23664 17196
rect 23716 17184 23722 17196
rect 24394 17184 24400 17196
rect 23716 17156 24400 17184
rect 23716 17144 23722 17156
rect 24394 17144 24400 17156
rect 24452 17144 24458 17196
rect 28620 17187 28678 17193
rect 28620 17153 28632 17187
rect 28666 17184 28678 17187
rect 33502 17184 33508 17196
rect 28666 17156 33508 17184
rect 28666 17153 28678 17156
rect 28620 17147 28678 17153
rect 33502 17144 33508 17156
rect 33560 17144 33566 17196
rect 33980 17193 34008 17224
rect 37458 17212 37464 17264
rect 37516 17252 37522 17264
rect 37614 17255 37672 17261
rect 37614 17252 37626 17255
rect 37516 17224 37626 17252
rect 37516 17212 37522 17224
rect 37614 17221 37626 17224
rect 37660 17221 37672 17255
rect 37752 17252 37780 17292
rect 38746 17280 38752 17292
rect 38804 17280 38810 17332
rect 40589 17323 40647 17329
rect 40589 17289 40601 17323
rect 40635 17320 40647 17323
rect 40678 17320 40684 17332
rect 40635 17292 40684 17320
rect 40635 17289 40647 17292
rect 40589 17283 40647 17289
rect 40678 17280 40684 17292
rect 40736 17280 40742 17332
rect 43806 17320 43812 17332
rect 43767 17292 43812 17320
rect 43806 17280 43812 17292
rect 43864 17280 43870 17332
rect 46290 17280 46296 17332
rect 46348 17320 46354 17332
rect 46385 17323 46443 17329
rect 46385 17320 46397 17323
rect 46348 17292 46397 17320
rect 46348 17280 46354 17292
rect 46385 17289 46397 17292
rect 46431 17289 46443 17323
rect 52178 17320 52184 17332
rect 52139 17292 52184 17320
rect 46385 17283 46443 17289
rect 52178 17280 52184 17292
rect 52236 17280 52242 17332
rect 57238 17280 57244 17332
rect 57296 17320 57302 17332
rect 57333 17323 57391 17329
rect 57333 17320 57345 17323
rect 57296 17292 57345 17320
rect 57296 17280 57302 17292
rect 57333 17289 57345 17292
rect 57379 17289 57391 17323
rect 57333 17283 57391 17289
rect 39454 17255 39512 17261
rect 39454 17252 39466 17255
rect 37752 17224 39466 17252
rect 37614 17215 37672 17221
rect 39454 17221 39466 17224
rect 39500 17221 39512 17255
rect 50798 17252 50804 17264
rect 39454 17215 39512 17221
rect 48976 17224 50804 17252
rect 33965 17187 34023 17193
rect 33965 17153 33977 17187
rect 34011 17153 34023 17187
rect 33965 17147 34023 17153
rect 34232 17187 34290 17193
rect 34232 17153 34244 17187
rect 34278 17184 34290 17187
rect 37274 17184 37280 17196
rect 34278 17156 37280 17184
rect 34278 17153 34290 17156
rect 34232 17147 34290 17153
rect 37274 17144 37280 17156
rect 37332 17144 37338 17196
rect 37366 17144 37372 17196
rect 37424 17184 37430 17196
rect 37424 17156 37469 17184
rect 37424 17144 37430 17156
rect 37918 17144 37924 17196
rect 37976 17184 37982 17196
rect 39209 17187 39267 17193
rect 39209 17184 39221 17187
rect 37976 17156 39221 17184
rect 37976 17144 37982 17156
rect 39209 17153 39221 17156
rect 39255 17153 39267 17187
rect 39209 17147 39267 17153
rect 42696 17187 42754 17193
rect 42696 17153 42708 17187
rect 42742 17184 42754 17187
rect 43898 17184 43904 17196
rect 42742 17156 43904 17184
rect 42742 17153 42754 17156
rect 42696 17147 42754 17153
rect 43898 17144 43904 17156
rect 43956 17144 43962 17196
rect 45002 17184 45008 17196
rect 44963 17156 45008 17184
rect 45002 17144 45008 17156
rect 45060 17144 45066 17196
rect 45272 17187 45330 17193
rect 45272 17153 45284 17187
rect 45318 17184 45330 17187
rect 46382 17184 46388 17196
rect 45318 17156 46388 17184
rect 45318 17153 45330 17156
rect 45272 17147 45330 17153
rect 46382 17144 46388 17156
rect 46440 17144 46446 17196
rect 47210 17144 47216 17196
rect 47268 17184 47274 17196
rect 48976 17193 49004 17224
rect 50798 17212 50804 17224
rect 50856 17212 50862 17264
rect 54380 17255 54438 17261
rect 54380 17221 54392 17255
rect 54426 17252 54438 17255
rect 55858 17252 55864 17264
rect 54426 17224 55864 17252
rect 54426 17221 54438 17224
rect 54380 17215 54438 17221
rect 55858 17212 55864 17224
rect 55916 17212 55922 17264
rect 56220 17255 56278 17261
rect 56220 17221 56232 17255
rect 56266 17252 56278 17255
rect 58158 17252 58164 17264
rect 56266 17224 58164 17252
rect 56266 17221 56278 17224
rect 56220 17215 56278 17221
rect 58158 17212 58164 17224
rect 58216 17212 58222 17264
rect 48961 17187 49019 17193
rect 48961 17184 48973 17187
rect 47268 17156 48973 17184
rect 47268 17144 47274 17156
rect 48961 17153 48973 17156
rect 49007 17153 49019 17187
rect 48961 17147 49019 17153
rect 49228 17187 49286 17193
rect 49228 17153 49240 17187
rect 49274 17184 49286 17187
rect 50890 17184 50896 17196
rect 49274 17156 50896 17184
rect 49274 17153 49286 17156
rect 49228 17147 49286 17153
rect 50890 17144 50896 17156
rect 50948 17144 50954 17196
rect 51068 17187 51126 17193
rect 51068 17153 51080 17187
rect 51114 17184 51126 17187
rect 52914 17184 52920 17196
rect 51114 17156 52920 17184
rect 51114 17153 51126 17156
rect 51068 17147 51126 17153
rect 52914 17144 52920 17156
rect 52972 17144 52978 17196
rect 53834 17144 53840 17196
rect 53892 17184 53898 17196
rect 54113 17187 54171 17193
rect 54113 17184 54125 17187
rect 53892 17156 54125 17184
rect 53892 17144 53898 17156
rect 54113 17153 54125 17156
rect 54159 17184 54171 17187
rect 55950 17184 55956 17196
rect 54159 17156 55956 17184
rect 54159 17153 54171 17156
rect 54113 17147 54171 17153
rect 55950 17144 55956 17156
rect 56008 17144 56014 17196
rect 27614 17076 27620 17128
rect 27672 17116 27678 17128
rect 28353 17119 28411 17125
rect 28353 17116 28365 17119
rect 27672 17088 28365 17116
rect 27672 17076 27678 17088
rect 28353 17085 28365 17088
rect 28399 17085 28411 17119
rect 28353 17079 28411 17085
rect 4706 16940 4712 16992
rect 4764 16980 4770 16992
rect 5721 16983 5779 16989
rect 5721 16980 5733 16983
rect 4764 16952 5733 16980
rect 4764 16940 4770 16952
rect 5721 16949 5733 16952
rect 5767 16949 5779 16983
rect 15470 16980 15476 16992
rect 15431 16952 15476 16980
rect 5721 16943 5779 16949
rect 15470 16940 15476 16952
rect 15528 16940 15534 16992
rect 18601 16983 18659 16989
rect 18601 16949 18613 16983
rect 18647 16980 18659 16983
rect 19334 16980 19340 16992
rect 18647 16952 19340 16980
rect 18647 16949 18659 16952
rect 18601 16943 18659 16949
rect 19334 16940 19340 16952
rect 19392 16940 19398 16992
rect 25774 16980 25780 16992
rect 25735 16952 25780 16980
rect 25774 16940 25780 16952
rect 25832 16940 25838 16992
rect 28368 16980 28396 17079
rect 29914 17076 29920 17128
rect 29972 17116 29978 17128
rect 30193 17119 30251 17125
rect 30193 17116 30205 17119
rect 29972 17088 30205 17116
rect 29972 17076 29978 17088
rect 30193 17085 30205 17088
rect 30239 17085 30251 17119
rect 30193 17079 30251 17085
rect 32125 17119 32183 17125
rect 32125 17085 32137 17119
rect 32171 17085 32183 17119
rect 42426 17116 42432 17128
rect 42387 17088 42432 17116
rect 32125 17079 32183 17085
rect 29730 17048 29736 17060
rect 29691 17020 29736 17048
rect 29730 17008 29736 17020
rect 29788 17008 29794 17060
rect 32140 17048 32168 17079
rect 42426 17076 42432 17088
rect 42484 17076 42490 17128
rect 50798 17116 50804 17128
rect 50759 17088 50804 17116
rect 50798 17076 50804 17088
rect 50856 17076 50862 17128
rect 31128 17020 32168 17048
rect 31128 16980 31156 17020
rect 28368 16952 31156 16980
rect 31573 16983 31631 16989
rect 31573 16949 31585 16983
rect 31619 16980 31631 16983
rect 32306 16980 32312 16992
rect 31619 16952 32312 16980
rect 31619 16949 31631 16952
rect 31573 16943 31631 16949
rect 32306 16940 32312 16952
rect 32364 16940 32370 16992
rect 33226 16940 33232 16992
rect 33284 16980 33290 16992
rect 33505 16983 33563 16989
rect 33505 16980 33517 16983
rect 33284 16952 33517 16980
rect 33284 16940 33290 16952
rect 33505 16949 33517 16952
rect 33551 16949 33563 16983
rect 33505 16943 33563 16949
rect 49326 16940 49332 16992
rect 49384 16980 49390 16992
rect 50341 16983 50399 16989
rect 50341 16980 50353 16983
rect 49384 16952 50353 16980
rect 49384 16940 49390 16952
rect 50341 16949 50353 16952
rect 50387 16949 50399 16983
rect 55490 16980 55496 16992
rect 55451 16952 55496 16980
rect 50341 16943 50399 16949
rect 55490 16940 55496 16952
rect 55548 16940 55554 16992
rect 1104 16890 59340 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 59340 16890
rect 1104 16816 59340 16838
rect 5166 16776 5172 16788
rect 5127 16748 5172 16776
rect 5166 16736 5172 16748
rect 5224 16736 5230 16788
rect 7006 16776 7012 16788
rect 6967 16748 7012 16776
rect 7006 16736 7012 16748
rect 7064 16736 7070 16788
rect 9306 16776 9312 16788
rect 8956 16748 9312 16776
rect 8956 16649 8984 16748
rect 9306 16736 9312 16748
rect 9364 16736 9370 16788
rect 10226 16736 10232 16788
rect 10284 16776 10290 16788
rect 10321 16779 10379 16785
rect 10321 16776 10333 16779
rect 10284 16748 10333 16776
rect 10284 16736 10290 16748
rect 10321 16745 10333 16748
rect 10367 16745 10379 16779
rect 12158 16776 12164 16788
rect 12119 16748 12164 16776
rect 10321 16739 10379 16745
rect 12158 16736 12164 16748
rect 12216 16736 12222 16788
rect 15473 16779 15531 16785
rect 15473 16745 15485 16779
rect 15519 16776 15531 16779
rect 15838 16776 15844 16788
rect 15519 16748 15844 16776
rect 15519 16745 15531 16748
rect 15473 16739 15531 16745
rect 15838 16736 15844 16748
rect 15896 16736 15902 16788
rect 18506 16776 18512 16788
rect 18467 16748 18512 16776
rect 18506 16736 18512 16748
rect 18564 16736 18570 16788
rect 37274 16736 37280 16788
rect 37332 16776 37338 16788
rect 37461 16779 37519 16785
rect 37461 16776 37473 16779
rect 37332 16748 37473 16776
rect 37332 16736 37338 16748
rect 37461 16745 37473 16748
rect 37507 16745 37519 16779
rect 43898 16776 43904 16788
rect 43859 16748 43904 16776
rect 37461 16739 37519 16745
rect 43898 16736 43904 16748
rect 43956 16736 43962 16788
rect 46382 16776 46388 16788
rect 46343 16748 46388 16776
rect 46382 16736 46388 16748
rect 46440 16736 46446 16788
rect 48774 16776 48780 16788
rect 48735 16748 48780 16776
rect 48774 16736 48780 16748
rect 48832 16736 48838 16788
rect 52914 16776 52920 16788
rect 52875 16748 52920 16776
rect 52914 16736 52920 16748
rect 52972 16736 52978 16788
rect 8941 16643 8999 16649
rect 8941 16609 8953 16643
rect 8987 16609 8999 16643
rect 8941 16603 8999 16609
rect 13998 16600 14004 16652
rect 14056 16640 14062 16652
rect 14093 16643 14151 16649
rect 14093 16640 14105 16643
rect 14056 16612 14105 16640
rect 14056 16600 14062 16612
rect 14093 16609 14105 16612
rect 14139 16609 14151 16643
rect 24394 16640 24400 16652
rect 24355 16612 24400 16640
rect 14093 16603 14151 16609
rect 24394 16600 24400 16612
rect 24452 16600 24458 16652
rect 36078 16640 36084 16652
rect 36039 16612 36084 16640
rect 36078 16600 36084 16612
rect 36136 16600 36142 16652
rect 37826 16600 37832 16652
rect 37884 16640 37890 16652
rect 37921 16643 37979 16649
rect 37921 16640 37933 16643
rect 37884 16612 37933 16640
rect 37884 16600 37890 16612
rect 37921 16609 37933 16612
rect 37967 16609 37979 16643
rect 37921 16603 37979 16609
rect 39758 16600 39764 16652
rect 39816 16640 39822 16652
rect 40681 16643 40739 16649
rect 40681 16640 40693 16643
rect 39816 16612 40693 16640
rect 39816 16600 39822 16612
rect 40681 16609 40693 16612
rect 40727 16609 40739 16643
rect 40681 16603 40739 16609
rect 42426 16600 42432 16652
rect 42484 16640 42490 16652
rect 42521 16643 42579 16649
rect 42521 16640 42533 16643
rect 42484 16612 42533 16640
rect 42484 16600 42490 16612
rect 42521 16609 42533 16612
rect 42567 16609 42579 16643
rect 47394 16640 47400 16652
rect 42521 16603 42579 16609
rect 46032 16612 47400 16640
rect 2682 16532 2688 16584
rect 2740 16572 2746 16584
rect 3789 16575 3847 16581
rect 3789 16572 3801 16575
rect 2740 16544 3801 16572
rect 2740 16532 2746 16544
rect 3789 16541 3801 16544
rect 3835 16541 3847 16575
rect 3789 16535 3847 16541
rect 4056 16575 4114 16581
rect 4056 16541 4068 16575
rect 4102 16572 4114 16575
rect 4614 16572 4620 16584
rect 4102 16544 4620 16572
rect 4102 16541 4114 16544
rect 4056 16535 4114 16541
rect 4614 16532 4620 16544
rect 4672 16532 4678 16584
rect 5534 16532 5540 16584
rect 5592 16572 5598 16584
rect 5629 16575 5687 16581
rect 5629 16572 5641 16575
rect 5592 16544 5641 16572
rect 5592 16532 5598 16544
rect 5629 16541 5641 16544
rect 5675 16541 5687 16575
rect 5629 16535 5687 16541
rect 9208 16575 9266 16581
rect 9208 16541 9220 16575
rect 9254 16572 9266 16575
rect 9582 16572 9588 16584
rect 9254 16544 9588 16572
rect 9254 16541 9266 16544
rect 9208 16535 9266 16541
rect 9582 16532 9588 16544
rect 9640 16532 9646 16584
rect 10410 16532 10416 16584
rect 10468 16572 10474 16584
rect 10781 16575 10839 16581
rect 10781 16572 10793 16575
rect 10468 16544 10793 16572
rect 10468 16532 10474 16544
rect 10781 16541 10793 16544
rect 10827 16541 10839 16575
rect 10781 16535 10839 16541
rect 11048 16575 11106 16581
rect 11048 16541 11060 16575
rect 11094 16572 11106 16575
rect 11330 16572 11336 16584
rect 11094 16544 11336 16572
rect 11094 16541 11106 16544
rect 11048 16535 11106 16541
rect 11330 16532 11336 16544
rect 11388 16532 11394 16584
rect 14360 16575 14418 16581
rect 14360 16541 14372 16575
rect 14406 16572 14418 16575
rect 15470 16572 15476 16584
rect 14406 16544 15476 16572
rect 14406 16541 14418 16544
rect 14360 16535 14418 16541
rect 15470 16532 15476 16544
rect 15528 16532 15534 16584
rect 16666 16532 16672 16584
rect 16724 16572 16730 16584
rect 17129 16575 17187 16581
rect 17129 16572 17141 16575
rect 16724 16544 17141 16572
rect 16724 16532 16730 16544
rect 17129 16541 17141 16544
rect 17175 16541 17187 16575
rect 17129 16535 17187 16541
rect 19150 16532 19156 16584
rect 19208 16572 19214 16584
rect 20898 16572 20904 16584
rect 19208 16544 20904 16572
rect 19208 16532 19214 16544
rect 20898 16532 20904 16544
rect 20956 16532 20962 16584
rect 24664 16575 24722 16581
rect 24664 16541 24676 16575
rect 24710 16572 24722 16575
rect 25774 16572 25780 16584
rect 24710 16544 25780 16572
rect 24710 16541 24722 16544
rect 24664 16535 24722 16541
rect 25774 16532 25780 16544
rect 25832 16532 25838 16584
rect 26234 16532 26240 16584
rect 26292 16572 26298 16584
rect 31021 16575 31079 16581
rect 26292 16544 26337 16572
rect 26292 16532 26298 16544
rect 31021 16541 31033 16575
rect 31067 16572 31079 16575
rect 31754 16572 31760 16584
rect 31067 16544 31760 16572
rect 31067 16541 31079 16544
rect 31021 16535 31079 16541
rect 31754 16532 31760 16544
rect 31812 16532 31818 16584
rect 36354 16581 36360 16584
rect 36348 16535 36360 16581
rect 36412 16572 36418 16584
rect 45002 16572 45008 16584
rect 36412 16544 36448 16572
rect 44963 16544 45008 16572
rect 36354 16532 36360 16535
rect 36412 16532 36418 16544
rect 45002 16532 45008 16544
rect 45060 16572 45066 16584
rect 46032 16572 46060 16612
rect 47394 16600 47400 16612
rect 47452 16600 47458 16652
rect 53377 16643 53435 16649
rect 53377 16640 53389 16643
rect 52564 16612 53389 16640
rect 45060 16544 46060 16572
rect 47664 16575 47722 16581
rect 45060 16532 45066 16544
rect 47664 16541 47676 16575
rect 47710 16572 47722 16575
rect 49326 16572 49332 16584
rect 47710 16544 49332 16572
rect 47710 16541 47722 16544
rect 47664 16535 47722 16541
rect 49326 16532 49332 16544
rect 49384 16532 49390 16584
rect 51534 16572 51540 16584
rect 51495 16544 51540 16572
rect 51534 16532 51540 16544
rect 51592 16532 51598 16584
rect 51810 16581 51816 16584
rect 51804 16535 51816 16581
rect 51868 16572 51874 16584
rect 52564 16572 52592 16612
rect 53377 16609 53389 16612
rect 53423 16609 53435 16643
rect 53377 16603 53435 16609
rect 51868 16544 51904 16572
rect 52380 16544 52592 16572
rect 51810 16532 51816 16535
rect 51868 16532 51874 16544
rect 5896 16507 5954 16513
rect 5896 16473 5908 16507
rect 5942 16504 5954 16507
rect 7742 16504 7748 16516
rect 5942 16476 7748 16504
rect 5942 16473 5954 16476
rect 5896 16467 5954 16473
rect 7742 16464 7748 16476
rect 7800 16464 7806 16516
rect 9306 16464 9312 16516
rect 9364 16504 9370 16516
rect 10428 16504 10456 16532
rect 9364 16476 10456 16504
rect 17396 16507 17454 16513
rect 9364 16464 9370 16476
rect 17396 16473 17408 16507
rect 17442 16504 17454 16507
rect 19242 16504 19248 16516
rect 17442 16476 19248 16504
rect 17442 16473 17454 16476
rect 17396 16467 17454 16473
rect 19242 16464 19248 16476
rect 19300 16464 19306 16516
rect 21168 16507 21226 16513
rect 21168 16473 21180 16507
rect 21214 16504 21226 16507
rect 23474 16504 23480 16516
rect 21214 16476 23480 16504
rect 21214 16473 21226 16476
rect 21168 16467 21226 16473
rect 23474 16464 23480 16476
rect 23532 16464 23538 16516
rect 25866 16464 25872 16516
rect 25924 16504 25930 16516
rect 26482 16507 26540 16513
rect 26482 16504 26494 16507
rect 25924 16476 26494 16504
rect 25924 16464 25930 16476
rect 26482 16473 26494 16476
rect 26528 16473 26540 16507
rect 26482 16467 26540 16473
rect 31288 16507 31346 16513
rect 31288 16473 31300 16507
rect 31334 16504 31346 16507
rect 31846 16504 31852 16516
rect 31334 16476 31852 16504
rect 31334 16473 31346 16476
rect 31288 16467 31346 16473
rect 31846 16464 31852 16476
rect 31904 16464 31910 16516
rect 38188 16507 38246 16513
rect 38188 16473 38200 16507
rect 38234 16504 38246 16507
rect 39850 16504 39856 16516
rect 38234 16476 39856 16504
rect 38234 16473 38246 16476
rect 38188 16467 38246 16473
rect 39850 16464 39856 16476
rect 39908 16464 39914 16516
rect 40948 16507 41006 16513
rect 40948 16473 40960 16507
rect 40994 16504 41006 16507
rect 42610 16504 42616 16516
rect 40994 16476 42616 16504
rect 40994 16473 41006 16476
rect 40948 16467 41006 16473
rect 42610 16464 42616 16476
rect 42668 16464 42674 16516
rect 42788 16507 42846 16513
rect 42788 16473 42800 16507
rect 42834 16504 42846 16507
rect 43806 16504 43812 16516
rect 42834 16476 43812 16504
rect 42834 16473 42846 16476
rect 42788 16467 42846 16473
rect 43806 16464 43812 16476
rect 43864 16464 43870 16516
rect 45272 16507 45330 16513
rect 45272 16473 45284 16507
rect 45318 16504 45330 16507
rect 46382 16504 46388 16516
rect 45318 16476 46388 16504
rect 45318 16473 45330 16476
rect 45272 16467 45330 16473
rect 46382 16464 46388 16476
rect 46440 16464 46446 16516
rect 51552 16504 51580 16532
rect 52380 16504 52408 16544
rect 55950 16532 55956 16584
rect 56008 16572 56014 16584
rect 56505 16575 56563 16581
rect 56505 16572 56517 16575
rect 56008 16544 56517 16572
rect 56008 16532 56014 16544
rect 56505 16541 56517 16544
rect 56551 16541 56563 16575
rect 56505 16535 56563 16541
rect 51552 16476 52408 16504
rect 53644 16507 53702 16513
rect 53644 16473 53656 16507
rect 53690 16504 53702 16507
rect 55398 16504 55404 16516
rect 53690 16476 55404 16504
rect 53690 16473 53702 16476
rect 53644 16467 53702 16473
rect 55398 16464 55404 16476
rect 55456 16464 55462 16516
rect 56772 16507 56830 16513
rect 56772 16473 56784 16507
rect 56818 16504 56830 16507
rect 57790 16504 57796 16516
rect 56818 16476 57796 16504
rect 56818 16473 56830 16476
rect 56772 16467 56830 16473
rect 57790 16464 57796 16476
rect 57848 16464 57854 16516
rect 22278 16436 22284 16448
rect 22239 16408 22284 16436
rect 22278 16396 22284 16408
rect 22336 16396 22342 16448
rect 25774 16436 25780 16448
rect 25735 16408 25780 16436
rect 25774 16396 25780 16408
rect 25832 16396 25838 16448
rect 27062 16396 27068 16448
rect 27120 16436 27126 16448
rect 27617 16439 27675 16445
rect 27617 16436 27629 16439
rect 27120 16408 27629 16436
rect 27120 16396 27126 16408
rect 27617 16405 27629 16408
rect 27663 16405 27675 16439
rect 27617 16399 27675 16405
rect 32214 16396 32220 16448
rect 32272 16436 32278 16448
rect 32401 16439 32459 16445
rect 32401 16436 32413 16439
rect 32272 16408 32413 16436
rect 32272 16396 32278 16408
rect 32401 16405 32413 16408
rect 32447 16405 32459 16439
rect 32401 16399 32459 16405
rect 39301 16439 39359 16445
rect 39301 16405 39313 16439
rect 39347 16436 39359 16439
rect 39942 16436 39948 16448
rect 39347 16408 39948 16436
rect 39347 16405 39359 16408
rect 39301 16399 39359 16405
rect 39942 16396 39948 16408
rect 40000 16396 40006 16448
rect 42058 16436 42064 16448
rect 42019 16408 42064 16436
rect 42058 16396 42064 16408
rect 42116 16396 42122 16448
rect 54754 16436 54760 16448
rect 54715 16408 54760 16436
rect 54754 16396 54760 16408
rect 54812 16396 54818 16448
rect 57882 16436 57888 16448
rect 57843 16408 57888 16436
rect 57882 16396 57888 16408
rect 57940 16396 57946 16448
rect 1104 16346 59340 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 59340 16346
rect 1104 16272 59340 16294
rect 7742 16232 7748 16244
rect 7703 16204 7748 16232
rect 7742 16192 7748 16204
rect 7800 16192 7806 16244
rect 8386 16192 8392 16244
rect 8444 16232 8450 16244
rect 8444 16204 8524 16232
rect 8444 16192 8450 16204
rect 3596 16167 3654 16173
rect 3596 16133 3608 16167
rect 3642 16164 3654 16167
rect 4706 16164 4712 16176
rect 3642 16136 4712 16164
rect 3642 16133 3654 16136
rect 3596 16127 3654 16133
rect 4706 16124 4712 16136
rect 4764 16124 4770 16176
rect 8496 16173 8524 16204
rect 9398 16192 9404 16244
rect 9456 16232 9462 16244
rect 9585 16235 9643 16241
rect 9585 16232 9597 16235
rect 9456 16204 9597 16232
rect 9456 16192 9462 16204
rect 9585 16201 9597 16204
rect 9631 16201 9643 16235
rect 9585 16195 9643 16201
rect 19334 16192 19340 16244
rect 19392 16232 19398 16244
rect 20530 16232 20536 16244
rect 19392 16204 19472 16232
rect 20491 16204 20536 16232
rect 19392 16192 19398 16204
rect 8472 16167 8530 16173
rect 6380 16136 8248 16164
rect 1756 16099 1814 16105
rect 1756 16065 1768 16099
rect 1802 16096 1814 16099
rect 1802 16068 4752 16096
rect 1802 16065 1814 16068
rect 1756 16059 1814 16065
rect 1489 16031 1547 16037
rect 1489 15997 1501 16031
rect 1535 15997 1547 16031
rect 2682 16028 2688 16040
rect 2595 16000 2688 16028
rect 1489 15991 1547 15997
rect 1504 15892 1532 15991
rect 2682 15988 2688 16000
rect 2740 16028 2746 16040
rect 3329 16031 3387 16037
rect 3329 16028 3341 16031
rect 2740 16000 3341 16028
rect 2740 15988 2746 16000
rect 3329 15997 3341 16000
rect 3375 15997 3387 16031
rect 3329 15991 3387 15997
rect 1762 15892 1768 15904
rect 1504 15864 1768 15892
rect 1762 15852 1768 15864
rect 1820 15892 1826 15904
rect 2700 15892 2728 15988
rect 4724 15969 4752 16068
rect 5534 15988 5540 16040
rect 5592 16028 5598 16040
rect 6380 16037 6408 16136
rect 6632 16099 6690 16105
rect 6632 16065 6644 16099
rect 6678 16096 6690 16099
rect 6914 16096 6920 16108
rect 6678 16068 6920 16096
rect 6678 16065 6690 16068
rect 6632 16059 6690 16065
rect 6914 16056 6920 16068
rect 6972 16056 6978 16108
rect 8220 16105 8248 16136
rect 8472 16133 8484 16167
rect 8518 16133 8530 16167
rect 8472 16127 8530 16133
rect 14636 16167 14694 16173
rect 14636 16133 14648 16167
rect 14682 16164 14694 16167
rect 15746 16164 15752 16176
rect 14682 16136 15752 16164
rect 14682 16133 14694 16136
rect 14636 16127 14694 16133
rect 15746 16124 15752 16136
rect 15804 16124 15810 16176
rect 19444 16173 19472 16204
rect 20530 16192 20536 16204
rect 20588 16192 20594 16244
rect 23198 16232 23204 16244
rect 23159 16204 23204 16232
rect 23198 16192 23204 16204
rect 23256 16192 23262 16244
rect 26234 16232 26240 16244
rect 24412 16204 26240 16232
rect 19420 16167 19478 16173
rect 17328 16136 19196 16164
rect 17328 16108 17356 16136
rect 19168 16108 19196 16136
rect 19420 16133 19432 16167
rect 19466 16133 19478 16167
rect 19420 16127 19478 16133
rect 22088 16167 22146 16173
rect 22088 16133 22100 16167
rect 22134 16164 22146 16167
rect 22278 16164 22284 16176
rect 22134 16136 22284 16164
rect 22134 16133 22146 16136
rect 22088 16127 22146 16133
rect 22278 16124 22284 16136
rect 22336 16124 22342 16176
rect 24412 16108 24440 16204
rect 26234 16192 26240 16204
rect 26292 16232 26298 16244
rect 26786 16232 26792 16244
rect 26292 16204 26792 16232
rect 26292 16192 26298 16204
rect 26786 16192 26792 16204
rect 26844 16192 26850 16244
rect 31570 16232 31576 16244
rect 31531 16204 31576 16232
rect 31570 16192 31576 16204
rect 31628 16192 31634 16244
rect 32306 16192 32312 16244
rect 32364 16232 32370 16244
rect 33502 16232 33508 16244
rect 32364 16204 32444 16232
rect 33463 16204 33508 16232
rect 32364 16192 32370 16204
rect 24664 16167 24722 16173
rect 24664 16133 24676 16167
rect 24710 16164 24722 16167
rect 25774 16164 25780 16176
rect 24710 16136 25780 16164
rect 24710 16133 24722 16136
rect 24664 16127 24722 16133
rect 25774 16124 25780 16136
rect 25832 16124 25838 16176
rect 30460 16167 30518 16173
rect 30460 16133 30472 16167
rect 30506 16164 30518 16167
rect 32214 16164 32220 16176
rect 30506 16136 32220 16164
rect 30506 16133 30518 16136
rect 30460 16127 30518 16133
rect 32214 16124 32220 16136
rect 32272 16124 32278 16176
rect 32416 16173 32444 16204
rect 33502 16192 33508 16204
rect 33560 16192 33566 16244
rect 43806 16232 43812 16244
rect 43767 16204 43812 16232
rect 43806 16192 43812 16204
rect 43864 16192 43870 16244
rect 46382 16232 46388 16244
rect 46343 16204 46388 16232
rect 46382 16192 46388 16204
rect 46440 16192 46446 16244
rect 50890 16192 50896 16244
rect 50948 16232 50954 16244
rect 51721 16235 51779 16241
rect 51721 16232 51733 16235
rect 50948 16204 51733 16232
rect 50948 16192 50954 16204
rect 51721 16201 51733 16204
rect 51767 16201 51779 16235
rect 57330 16232 57336 16244
rect 57291 16204 57336 16232
rect 51721 16195 51779 16201
rect 57330 16192 57336 16204
rect 57388 16192 57394 16244
rect 32392 16167 32450 16173
rect 32392 16133 32404 16167
rect 32438 16133 32450 16167
rect 32392 16127 32450 16133
rect 34790 16124 34796 16176
rect 34848 16164 34854 16176
rect 34946 16167 35004 16173
rect 34946 16164 34958 16167
rect 34848 16136 34958 16164
rect 34848 16124 34854 16136
rect 34946 16133 34958 16136
rect 34992 16133 35004 16167
rect 39758 16164 39764 16176
rect 34946 16127 35004 16133
rect 37936 16136 39764 16164
rect 8205 16099 8263 16105
rect 8205 16065 8217 16099
rect 8251 16065 8263 16099
rect 8205 16059 8263 16065
rect 14274 16056 14280 16108
rect 14332 16096 14338 16108
rect 14369 16099 14427 16105
rect 14369 16096 14381 16099
rect 14332 16068 14381 16096
rect 14332 16056 14338 16068
rect 14369 16065 14381 16068
rect 14415 16096 14427 16099
rect 16666 16096 16672 16108
rect 14415 16068 16672 16096
rect 14415 16065 14427 16068
rect 14369 16059 14427 16065
rect 16666 16056 16672 16068
rect 16724 16056 16730 16108
rect 17310 16096 17316 16108
rect 17271 16068 17316 16096
rect 17310 16056 17316 16068
rect 17368 16056 17374 16108
rect 17580 16099 17638 16105
rect 17580 16065 17592 16099
rect 17626 16096 17638 16099
rect 18690 16096 18696 16108
rect 17626 16068 18696 16096
rect 17626 16065 17638 16068
rect 17580 16059 17638 16065
rect 18690 16056 18696 16068
rect 18748 16056 18754 16108
rect 19150 16096 19156 16108
rect 19063 16068 19156 16096
rect 19150 16056 19156 16068
rect 19208 16056 19214 16108
rect 24394 16096 24400 16108
rect 24307 16068 24400 16096
rect 24394 16056 24400 16068
rect 24452 16056 24458 16108
rect 26326 16056 26332 16108
rect 26384 16096 26390 16108
rect 27229 16099 27287 16105
rect 27229 16096 27241 16099
rect 26384 16068 27241 16096
rect 26384 16056 26390 16068
rect 27229 16065 27241 16068
rect 27275 16065 27287 16099
rect 27229 16059 27287 16065
rect 30193 16099 30251 16105
rect 30193 16065 30205 16099
rect 30239 16096 30251 16099
rect 31754 16096 31760 16108
rect 30239 16068 31760 16096
rect 30239 16065 30251 16068
rect 30193 16059 30251 16065
rect 31754 16056 31760 16068
rect 31812 16096 31818 16108
rect 32125 16099 32183 16105
rect 32125 16096 32137 16099
rect 31812 16068 32137 16096
rect 31812 16056 31818 16068
rect 32125 16065 32137 16068
rect 32171 16096 32183 16099
rect 32858 16096 32864 16108
rect 32171 16068 32864 16096
rect 32171 16065 32183 16068
rect 32125 16059 32183 16065
rect 32858 16056 32864 16068
rect 32916 16056 32922 16108
rect 6365 16031 6423 16037
rect 6365 16028 6377 16031
rect 5592 16000 6377 16028
rect 5592 15988 5598 16000
rect 6365 15997 6377 16000
rect 6411 15997 6423 16031
rect 6365 15991 6423 15997
rect 20898 15988 20904 16040
rect 20956 16028 20962 16040
rect 21821 16031 21879 16037
rect 21821 16028 21833 16031
rect 20956 16000 21833 16028
rect 20956 15988 20962 16000
rect 21821 15997 21833 16000
rect 21867 15997 21879 16031
rect 21821 15991 21879 15997
rect 26786 15988 26792 16040
rect 26844 16028 26850 16040
rect 26973 16031 27031 16037
rect 26973 16028 26985 16031
rect 26844 16000 26985 16028
rect 26844 15988 26850 16000
rect 26973 15997 26985 16000
rect 27019 15997 27031 16031
rect 34698 16028 34704 16040
rect 34659 16000 34704 16028
rect 26973 15991 27031 15997
rect 34698 15988 34704 16000
rect 34756 15988 34762 16040
rect 37826 16028 37832 16040
rect 37739 16000 37832 16028
rect 37826 15988 37832 16000
rect 37884 16028 37890 16040
rect 37936 16028 37964 16136
rect 39758 16124 39764 16136
rect 39816 16124 39822 16176
rect 40144 16136 41368 16164
rect 38096 16099 38154 16105
rect 38096 16065 38108 16099
rect 38142 16096 38154 16099
rect 39022 16096 39028 16108
rect 38142 16068 39028 16096
rect 38142 16065 38154 16068
rect 38096 16059 38154 16065
rect 39022 16056 39028 16068
rect 39080 16056 39086 16108
rect 37884 16000 37964 16028
rect 37884 15988 37890 16000
rect 40034 15988 40040 16040
rect 40092 16028 40098 16040
rect 40144 16037 40172 16136
rect 40396 16099 40454 16105
rect 40396 16065 40408 16099
rect 40442 16096 40454 16099
rect 41230 16096 41236 16108
rect 40442 16068 41236 16096
rect 40442 16065 40454 16068
rect 40396 16059 40454 16065
rect 41230 16056 41236 16068
rect 41288 16056 41294 16108
rect 41340 16096 41368 16136
rect 42058 16124 42064 16176
rect 42116 16164 42122 16176
rect 42674 16167 42732 16173
rect 42674 16164 42686 16167
rect 42116 16136 42686 16164
rect 42116 16124 42122 16136
rect 42674 16133 42686 16136
rect 42720 16133 42732 16167
rect 42674 16127 42732 16133
rect 47940 16167 47998 16173
rect 47940 16133 47952 16167
rect 47986 16164 47998 16167
rect 49050 16164 49056 16176
rect 47986 16136 49056 16164
rect 47986 16133 47998 16136
rect 47940 16127 47998 16133
rect 49050 16124 49056 16136
rect 49108 16124 49114 16176
rect 50614 16173 50620 16176
rect 50608 16164 50620 16173
rect 50575 16136 50620 16164
rect 50608 16127 50620 16136
rect 50614 16124 50620 16127
rect 50672 16124 50678 16176
rect 54380 16167 54438 16173
rect 54380 16133 54392 16167
rect 54426 16164 54438 16167
rect 55490 16164 55496 16176
rect 54426 16136 55496 16164
rect 54426 16133 54438 16136
rect 54380 16127 54438 16133
rect 55490 16124 55496 16136
rect 55548 16124 55554 16176
rect 56220 16167 56278 16173
rect 56220 16133 56232 16167
rect 56266 16164 56278 16167
rect 57882 16164 57888 16176
rect 56266 16136 57888 16164
rect 56266 16133 56278 16136
rect 56220 16127 56278 16133
rect 57882 16124 57888 16136
rect 57940 16124 57946 16176
rect 42426 16096 42432 16108
rect 41340 16068 42432 16096
rect 42426 16056 42432 16068
rect 42484 16056 42490 16108
rect 45002 16096 45008 16108
rect 44963 16068 45008 16096
rect 45002 16056 45008 16068
rect 45060 16056 45066 16108
rect 45272 16099 45330 16105
rect 45272 16065 45284 16099
rect 45318 16096 45330 16099
rect 46382 16096 46388 16108
rect 45318 16068 46388 16096
rect 45318 16065 45330 16068
rect 45272 16059 45330 16065
rect 46382 16056 46388 16068
rect 46440 16056 46446 16108
rect 50341 16099 50399 16105
rect 50341 16065 50353 16099
rect 50387 16096 50399 16099
rect 51534 16096 51540 16108
rect 50387 16068 51540 16096
rect 50387 16065 50399 16068
rect 50341 16059 50399 16065
rect 51534 16056 51540 16068
rect 51592 16096 51598 16108
rect 51994 16096 52000 16108
rect 51592 16068 52000 16096
rect 51592 16056 51598 16068
rect 51994 16056 52000 16068
rect 52052 16056 52058 16108
rect 40129 16031 40187 16037
rect 40129 16028 40141 16031
rect 40092 16000 40141 16028
rect 40092 15988 40098 16000
rect 40129 15997 40141 16000
rect 40175 15997 40187 16031
rect 40129 15991 40187 15997
rect 47578 15988 47584 16040
rect 47636 16028 47642 16040
rect 47673 16031 47731 16037
rect 47673 16028 47685 16031
rect 47636 16000 47685 16028
rect 47636 15988 47642 16000
rect 47673 15997 47685 16000
rect 47719 15997 47731 16031
rect 47673 15991 47731 15997
rect 54113 16031 54171 16037
rect 54113 15997 54125 16031
rect 54159 15997 54171 16031
rect 55950 16028 55956 16040
rect 54113 15991 54171 15997
rect 55186 16000 55956 16028
rect 4709 15963 4767 15969
rect 4709 15929 4721 15963
rect 4755 15929 4767 15963
rect 4709 15923 4767 15929
rect 2866 15892 2872 15904
rect 1820 15864 2728 15892
rect 2827 15864 2872 15892
rect 1820 15852 1826 15864
rect 2866 15852 2872 15864
rect 2924 15852 2930 15904
rect 15746 15892 15752 15904
rect 15707 15864 15752 15892
rect 15746 15852 15752 15864
rect 15804 15852 15810 15904
rect 18693 15895 18751 15901
rect 18693 15861 18705 15895
rect 18739 15892 18751 15895
rect 19334 15892 19340 15904
rect 18739 15864 19340 15892
rect 18739 15861 18751 15864
rect 18693 15855 18751 15861
rect 19334 15852 19340 15864
rect 19392 15852 19398 15904
rect 25774 15892 25780 15904
rect 25735 15864 25780 15892
rect 25774 15852 25780 15864
rect 25832 15852 25838 15904
rect 28350 15892 28356 15904
rect 28311 15864 28356 15892
rect 28350 15852 28356 15864
rect 28408 15852 28414 15904
rect 36078 15892 36084 15904
rect 36039 15864 36084 15892
rect 36078 15852 36084 15864
rect 36136 15852 36142 15904
rect 39206 15892 39212 15904
rect 39167 15864 39212 15892
rect 39206 15852 39212 15864
rect 39264 15852 39270 15904
rect 41506 15892 41512 15904
rect 41467 15864 41512 15892
rect 41506 15852 41512 15864
rect 41564 15852 41570 15904
rect 49050 15892 49056 15904
rect 49011 15864 49056 15892
rect 49050 15852 49056 15864
rect 49108 15852 49114 15904
rect 54128 15892 54156 15991
rect 55186 15892 55214 16000
rect 55950 15988 55956 16000
rect 56008 15988 56014 16040
rect 55398 15920 55404 15972
rect 55456 15960 55462 15972
rect 55493 15963 55551 15969
rect 55493 15960 55505 15963
rect 55456 15932 55505 15960
rect 55456 15920 55462 15932
rect 55493 15929 55505 15932
rect 55539 15929 55551 15963
rect 55493 15923 55551 15929
rect 54128 15864 55214 15892
rect 1104 15802 59340 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 59340 15802
rect 1104 15728 59340 15750
rect 6914 15648 6920 15700
rect 6972 15688 6978 15700
rect 18690 15688 18696 15700
rect 6972 15660 7017 15688
rect 18651 15660 18696 15688
rect 6972 15648 6978 15660
rect 18690 15648 18696 15660
rect 18748 15648 18754 15700
rect 20898 15648 20904 15700
rect 20956 15688 20962 15700
rect 21177 15691 21235 15697
rect 21177 15688 21189 15691
rect 20956 15660 21189 15688
rect 20956 15648 20962 15660
rect 21177 15657 21189 15660
rect 21223 15657 21235 15691
rect 23474 15688 23480 15700
rect 23435 15660 23480 15688
rect 21177 15651 21235 15657
rect 13998 15512 14004 15564
rect 14056 15552 14062 15564
rect 14369 15555 14427 15561
rect 14369 15552 14381 15555
rect 14056 15524 14381 15552
rect 14056 15512 14062 15524
rect 14369 15521 14381 15524
rect 14415 15521 14427 15555
rect 21192 15552 21220 15651
rect 23474 15648 23480 15660
rect 23532 15648 23538 15700
rect 25777 15691 25835 15697
rect 25777 15657 25789 15691
rect 25823 15688 25835 15691
rect 25866 15688 25872 15700
rect 25823 15660 25872 15688
rect 25823 15657 25835 15660
rect 25777 15651 25835 15657
rect 25866 15648 25872 15660
rect 25924 15648 25930 15700
rect 39022 15688 39028 15700
rect 38983 15660 39028 15688
rect 39022 15648 39028 15660
rect 39080 15648 39086 15700
rect 41230 15688 41236 15700
rect 41191 15660 41236 15688
rect 41230 15648 41236 15660
rect 41288 15648 41294 15700
rect 42610 15648 42616 15700
rect 42668 15688 42674 15700
rect 43073 15691 43131 15697
rect 43073 15688 43085 15691
rect 42668 15660 43085 15688
rect 42668 15648 42674 15660
rect 43073 15657 43085 15660
rect 43119 15657 43131 15691
rect 46382 15688 46388 15700
rect 46343 15660 46388 15688
rect 43073 15651 43131 15657
rect 46382 15648 46388 15660
rect 46440 15648 46446 15700
rect 57790 15688 57796 15700
rect 57751 15660 57796 15688
rect 57790 15648 57796 15660
rect 57848 15648 57854 15700
rect 22097 15555 22155 15561
rect 22097 15552 22109 15555
rect 21192 15524 22109 15552
rect 14369 15515 14427 15521
rect 22097 15521 22109 15524
rect 22143 15521 22155 15555
rect 24394 15552 24400 15564
rect 24355 15524 24400 15552
rect 22097 15515 22155 15521
rect 24394 15512 24400 15524
rect 24452 15512 24458 15564
rect 39758 15512 39764 15564
rect 39816 15552 39822 15564
rect 39853 15555 39911 15561
rect 39853 15552 39865 15555
rect 39816 15524 39865 15552
rect 39816 15512 39822 15524
rect 39853 15521 39865 15524
rect 39899 15521 39911 15555
rect 48130 15552 48136 15564
rect 39853 15515 39911 15521
rect 47872 15524 48136 15552
rect 1762 15444 1768 15496
rect 1820 15484 1826 15496
rect 1857 15487 1915 15493
rect 1857 15484 1869 15487
rect 1820 15456 1869 15484
rect 1820 15444 1826 15456
rect 1857 15453 1869 15456
rect 1903 15453 1915 15487
rect 1857 15447 1915 15453
rect 2124 15487 2182 15493
rect 2124 15453 2136 15487
rect 2170 15484 2182 15487
rect 2866 15484 2872 15496
rect 2170 15456 2872 15484
rect 2170 15453 2182 15456
rect 2124 15447 2182 15453
rect 2866 15444 2872 15456
rect 2924 15444 2930 15496
rect 5534 15484 5540 15496
rect 5495 15456 5540 15484
rect 5534 15444 5540 15456
rect 5592 15444 5598 15496
rect 9766 15444 9772 15496
rect 9824 15484 9830 15496
rect 10410 15484 10416 15496
rect 9824 15456 10416 15484
rect 9824 15444 9830 15456
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 14636 15487 14694 15493
rect 14636 15453 14648 15487
rect 14682 15484 14694 15487
rect 15746 15484 15752 15496
rect 14682 15456 15752 15484
rect 14682 15453 14694 15456
rect 14636 15447 14694 15453
rect 15746 15444 15752 15456
rect 15804 15444 15810 15496
rect 17310 15484 17316 15496
rect 17271 15456 17316 15484
rect 17310 15444 17316 15456
rect 17368 15444 17374 15496
rect 24664 15487 24722 15493
rect 24664 15453 24676 15487
rect 24710 15484 24722 15487
rect 25774 15484 25780 15496
rect 24710 15456 25780 15484
rect 24710 15453 24722 15456
rect 24664 15447 24722 15453
rect 25774 15444 25780 15456
rect 25832 15444 25838 15496
rect 26786 15484 26792 15496
rect 26747 15456 26792 15484
rect 26786 15444 26792 15456
rect 26844 15444 26850 15496
rect 27056 15487 27114 15493
rect 27056 15453 27068 15487
rect 27102 15484 27114 15487
rect 28350 15484 28356 15496
rect 27102 15456 28356 15484
rect 27102 15453 27114 15456
rect 27056 15447 27114 15453
rect 28350 15444 28356 15456
rect 28408 15444 28414 15496
rect 30745 15487 30803 15493
rect 30745 15453 30757 15487
rect 30791 15484 30803 15487
rect 32769 15487 32827 15493
rect 32769 15484 32781 15487
rect 30791 15456 32781 15484
rect 30791 15453 30803 15456
rect 30745 15447 30803 15453
rect 32769 15453 32781 15456
rect 32815 15484 32827 15487
rect 32858 15484 32864 15496
rect 32815 15456 32864 15484
rect 32815 15453 32827 15456
rect 32769 15447 32827 15453
rect 32858 15444 32864 15456
rect 32916 15444 32922 15496
rect 34606 15444 34612 15496
rect 34664 15484 34670 15496
rect 34701 15487 34759 15493
rect 34701 15484 34713 15487
rect 34664 15456 34713 15484
rect 34664 15444 34670 15456
rect 34701 15453 34713 15456
rect 34747 15453 34759 15487
rect 34701 15447 34759 15453
rect 34968 15487 35026 15493
rect 34968 15453 34980 15487
rect 35014 15484 35026 15487
rect 36078 15484 36084 15496
rect 35014 15456 36084 15484
rect 35014 15453 35026 15456
rect 34968 15447 35026 15453
rect 36078 15444 36084 15456
rect 36136 15444 36142 15496
rect 37645 15487 37703 15493
rect 37645 15453 37657 15487
rect 37691 15484 37703 15487
rect 37734 15484 37740 15496
rect 37691 15456 37740 15484
rect 37691 15453 37703 15456
rect 37645 15447 37703 15453
rect 37734 15444 37740 15456
rect 37792 15444 37798 15496
rect 39942 15444 39948 15496
rect 40000 15484 40006 15496
rect 40109 15487 40167 15493
rect 40109 15484 40121 15487
rect 40000 15456 40121 15484
rect 40000 15444 40006 15456
rect 40109 15453 40121 15456
rect 40155 15453 40167 15487
rect 40109 15447 40167 15453
rect 41693 15487 41751 15493
rect 41693 15453 41705 15487
rect 41739 15484 41751 15487
rect 45002 15484 45008 15496
rect 41739 15456 45008 15484
rect 41739 15453 41751 15456
rect 41693 15447 41751 15453
rect 45002 15444 45008 15456
rect 45060 15444 45066 15496
rect 47872 15493 47900 15524
rect 48130 15512 48136 15524
rect 48188 15552 48194 15564
rect 48188 15524 50292 15552
rect 48188 15512 48194 15524
rect 47857 15487 47915 15493
rect 47857 15453 47869 15487
rect 47903 15453 47915 15487
rect 50157 15487 50215 15493
rect 50157 15484 50169 15487
rect 47857 15447 47915 15453
rect 49528 15456 50169 15484
rect 5804 15419 5862 15425
rect 5804 15385 5816 15419
rect 5850 15416 5862 15419
rect 7926 15416 7932 15428
rect 5850 15388 7932 15416
rect 5850 15385 5862 15388
rect 5804 15379 5862 15385
rect 7926 15376 7932 15388
rect 7984 15376 7990 15428
rect 10680 15419 10738 15425
rect 10680 15385 10692 15419
rect 10726 15416 10738 15419
rect 12158 15416 12164 15428
rect 10726 15388 12164 15416
rect 10726 15385 10738 15388
rect 10680 15379 10738 15385
rect 12158 15376 12164 15388
rect 12216 15376 12222 15428
rect 17580 15419 17638 15425
rect 17580 15385 17592 15419
rect 17626 15416 17638 15419
rect 18782 15416 18788 15428
rect 17626 15388 18788 15416
rect 17626 15385 17638 15388
rect 17580 15379 17638 15385
rect 18782 15376 18788 15388
rect 18840 15376 18846 15428
rect 19426 15376 19432 15428
rect 19484 15416 19490 15428
rect 19889 15419 19947 15425
rect 19889 15416 19901 15419
rect 19484 15388 19901 15416
rect 19484 15376 19490 15388
rect 19889 15385 19901 15388
rect 19935 15385 19947 15419
rect 19889 15379 19947 15385
rect 22364 15419 22422 15425
rect 22364 15385 22376 15419
rect 22410 15416 22422 15419
rect 23658 15416 23664 15428
rect 22410 15388 23664 15416
rect 22410 15385 22422 15388
rect 22364 15379 22422 15385
rect 23658 15376 23664 15388
rect 23716 15376 23722 15428
rect 31012 15419 31070 15425
rect 31012 15385 31024 15419
rect 31058 15416 31070 15419
rect 33036 15419 33094 15425
rect 31058 15388 32996 15416
rect 31058 15385 31070 15388
rect 31012 15379 31070 15385
rect 3234 15348 3240 15360
rect 3195 15320 3240 15348
rect 3234 15308 3240 15320
rect 3292 15308 3298 15360
rect 11790 15348 11796 15360
rect 11751 15320 11796 15348
rect 11790 15308 11796 15320
rect 11848 15308 11854 15360
rect 15746 15348 15752 15360
rect 15707 15320 15752 15348
rect 15746 15308 15752 15320
rect 15804 15308 15810 15360
rect 28166 15348 28172 15360
rect 28127 15320 28172 15348
rect 28166 15308 28172 15320
rect 28224 15308 28230 15360
rect 32122 15348 32128 15360
rect 32083 15320 32128 15348
rect 32122 15308 32128 15320
rect 32180 15308 32186 15360
rect 32968 15348 32996 15388
rect 33036 15385 33048 15419
rect 33082 15416 33094 15419
rect 33962 15416 33968 15428
rect 33082 15388 33968 15416
rect 33082 15385 33094 15388
rect 33036 15379 33094 15385
rect 33962 15376 33968 15388
rect 34020 15376 34026 15428
rect 37912 15419 37970 15425
rect 37912 15385 37924 15419
rect 37958 15416 37970 15419
rect 38930 15416 38936 15428
rect 37958 15388 38936 15416
rect 37958 15385 37970 15388
rect 37912 15379 37970 15385
rect 38930 15376 38936 15388
rect 38988 15376 38994 15428
rect 41598 15376 41604 15428
rect 41656 15416 41662 15428
rect 41938 15419 41996 15425
rect 41938 15416 41950 15419
rect 41656 15388 41950 15416
rect 41656 15376 41662 15388
rect 41938 15385 41950 15388
rect 41984 15385 41996 15419
rect 41938 15379 41996 15385
rect 45272 15419 45330 15425
rect 45272 15385 45284 15419
rect 45318 15416 45330 15419
rect 46382 15416 46388 15428
rect 45318 15388 46388 15416
rect 45318 15385 45330 15388
rect 45272 15379 45330 15385
rect 46382 15376 46388 15388
rect 46440 15376 46446 15428
rect 49528 15360 49556 15456
rect 50157 15453 50169 15456
rect 50203 15453 50215 15487
rect 50264 15484 50292 15524
rect 51994 15484 52000 15496
rect 50264 15456 51580 15484
rect 51955 15456 52000 15484
rect 50157 15447 50215 15453
rect 50424 15419 50482 15425
rect 50424 15385 50436 15419
rect 50470 15416 50482 15419
rect 51442 15416 51448 15428
rect 50470 15388 51448 15416
rect 50470 15385 50482 15388
rect 50424 15379 50482 15385
rect 51442 15376 51448 15388
rect 51500 15376 51506 15428
rect 51552 15416 51580 15456
rect 51994 15444 52000 15456
rect 52052 15444 52058 15496
rect 55950 15444 55956 15496
rect 56008 15484 56014 15496
rect 56410 15484 56416 15496
rect 56008 15456 56416 15484
rect 56008 15444 56014 15456
rect 56410 15444 56416 15456
rect 56468 15444 56474 15496
rect 52264 15419 52322 15425
rect 51552 15388 52224 15416
rect 33686 15348 33692 15360
rect 32968 15320 33692 15348
rect 33686 15308 33692 15320
rect 33744 15308 33750 15360
rect 34146 15348 34152 15360
rect 34107 15320 34152 15348
rect 34146 15308 34152 15320
rect 34204 15308 34210 15360
rect 36078 15348 36084 15360
rect 36039 15320 36084 15348
rect 36078 15308 36084 15320
rect 36136 15308 36142 15360
rect 47578 15308 47584 15360
rect 47636 15348 47642 15360
rect 49145 15351 49203 15357
rect 49145 15348 49157 15351
rect 47636 15320 49157 15348
rect 47636 15308 47642 15320
rect 49145 15317 49157 15320
rect 49191 15348 49203 15351
rect 49510 15348 49516 15360
rect 49191 15320 49516 15348
rect 49191 15317 49203 15320
rect 49145 15311 49203 15317
rect 49510 15308 49516 15320
rect 49568 15308 49574 15360
rect 51537 15351 51595 15357
rect 51537 15317 51549 15351
rect 51583 15348 51595 15351
rect 52086 15348 52092 15360
rect 51583 15320 52092 15348
rect 51583 15317 51595 15320
rect 51537 15311 51595 15317
rect 52086 15308 52092 15320
rect 52144 15308 52150 15360
rect 52196 15348 52224 15388
rect 52264 15385 52276 15419
rect 52310 15416 52322 15419
rect 53282 15416 53288 15428
rect 52310 15388 53288 15416
rect 52310 15385 52322 15388
rect 52264 15379 52322 15385
rect 53282 15376 53288 15388
rect 53340 15376 53346 15428
rect 56680 15419 56738 15425
rect 56680 15385 56692 15419
rect 56726 15416 56738 15419
rect 57330 15416 57336 15428
rect 56726 15388 57336 15416
rect 56726 15385 56738 15388
rect 56680 15379 56738 15385
rect 57330 15376 57336 15388
rect 57388 15376 57394 15428
rect 53098 15348 53104 15360
rect 52196 15320 53104 15348
rect 53098 15308 53104 15320
rect 53156 15308 53162 15360
rect 53377 15351 53435 15357
rect 53377 15317 53389 15351
rect 53423 15348 53435 15351
rect 53742 15348 53748 15360
rect 53423 15320 53748 15348
rect 53423 15317 53435 15320
rect 53377 15311 53435 15317
rect 53742 15308 53748 15320
rect 53800 15308 53806 15360
rect 1104 15258 59340 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 59340 15258
rect 1104 15184 59340 15206
rect 7926 15144 7932 15156
rect 7887 15116 7932 15144
rect 7926 15104 7932 15116
rect 7984 15104 7990 15156
rect 18782 15144 18788 15156
rect 18743 15116 18788 15144
rect 18782 15104 18788 15116
rect 18840 15104 18846 15156
rect 19242 15104 19248 15156
rect 19300 15144 19306 15156
rect 20625 15147 20683 15153
rect 20625 15144 20637 15147
rect 19300 15116 20637 15144
rect 19300 15104 19306 15116
rect 20625 15113 20637 15116
rect 20671 15113 20683 15147
rect 26326 15144 26332 15156
rect 26287 15116 26332 15144
rect 20625 15107 20683 15113
rect 26326 15104 26332 15116
rect 26384 15104 26390 15156
rect 38930 15144 38936 15156
rect 38891 15116 38936 15144
rect 38930 15104 38936 15116
rect 38988 15104 38994 15156
rect 39850 15104 39856 15156
rect 39908 15144 39914 15156
rect 40865 15147 40923 15153
rect 40865 15144 40877 15147
rect 39908 15116 40877 15144
rect 39908 15104 39914 15116
rect 40865 15113 40877 15116
rect 40911 15113 40923 15147
rect 46382 15144 46388 15156
rect 46343 15116 46388 15144
rect 40865 15107 40923 15113
rect 46382 15104 46388 15116
rect 46440 15104 46446 15156
rect 57330 15144 57336 15156
rect 57291 15116 57336 15144
rect 57330 15104 57336 15116
rect 57388 15104 57394 15156
rect 1940 15079 1998 15085
rect 1940 15045 1952 15079
rect 1986 15076 1998 15079
rect 3234 15076 3240 15088
rect 1986 15048 3240 15076
rect 1986 15045 1998 15048
rect 1940 15039 1998 15045
rect 3234 15036 3240 15048
rect 3292 15036 3298 15088
rect 9766 15076 9772 15088
rect 8496 15048 9772 15076
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 1762 15008 1768 15020
rect 1719 14980 1768 15008
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 6816 15011 6874 15017
rect 6816 14977 6828 15011
rect 6862 15008 6874 15011
rect 8110 15008 8116 15020
rect 6862 14980 8116 15008
rect 6862 14977 6874 14980
rect 6816 14971 6874 14977
rect 8110 14968 8116 14980
rect 8168 14968 8174 15020
rect 8496 15017 8524 15048
rect 9766 15036 9772 15048
rect 9824 15036 9830 15088
rect 12520 15079 12578 15085
rect 12520 15045 12532 15079
rect 12566 15076 12578 15079
rect 14544 15079 14602 15085
rect 12566 15048 14504 15076
rect 12566 15045 12578 15048
rect 12520 15039 12578 15045
rect 8481 15011 8539 15017
rect 8481 14977 8493 15011
rect 8527 14977 8539 15011
rect 8481 14971 8539 14977
rect 8748 15011 8806 15017
rect 8748 14977 8760 15011
rect 8794 15008 8806 15011
rect 10962 15008 10968 15020
rect 8794 14980 10968 15008
rect 8794 14977 8806 14980
rect 8748 14971 8806 14977
rect 10962 14968 10968 14980
rect 11020 14968 11026 15020
rect 14274 15008 14280 15020
rect 14235 14980 14280 15008
rect 14274 14968 14280 14980
rect 14332 14968 14338 15020
rect 14476 15008 14504 15048
rect 14544 15045 14556 15079
rect 14590 15076 14602 15079
rect 15746 15076 15752 15088
rect 14590 15048 15752 15076
rect 14590 15045 14602 15048
rect 14544 15039 14602 15045
rect 15746 15036 15752 15048
rect 15804 15036 15810 15088
rect 23376 15079 23434 15085
rect 23376 15045 23388 15079
rect 23422 15076 23434 15079
rect 25216 15079 25274 15085
rect 23422 15048 25084 15076
rect 23422 15045 23434 15048
rect 23376 15039 23434 15045
rect 15378 15008 15384 15020
rect 14476 14980 15384 15008
rect 15378 14968 15384 14980
rect 15436 14968 15442 15020
rect 17672 15011 17730 15017
rect 17672 14977 17684 15011
rect 17718 15008 17730 15011
rect 18506 15008 18512 15020
rect 17718 14980 18512 15008
rect 17718 14977 17730 14980
rect 17672 14971 17730 14977
rect 18506 14968 18512 14980
rect 18564 14968 18570 15020
rect 19150 14968 19156 15020
rect 19208 15008 19214 15020
rect 19245 15011 19303 15017
rect 19245 15008 19257 15011
rect 19208 14980 19257 15008
rect 19208 14968 19214 14980
rect 19245 14977 19257 14980
rect 19291 14977 19303 15011
rect 19245 14971 19303 14977
rect 19334 14968 19340 15020
rect 19392 15008 19398 15020
rect 19501 15011 19559 15017
rect 19501 15008 19513 15011
rect 19392 14980 19513 15008
rect 19392 14968 19398 14980
rect 19501 14977 19513 14980
rect 19547 14977 19559 15011
rect 19501 14971 19559 14977
rect 23109 15011 23167 15017
rect 23109 14977 23121 15011
rect 23155 15008 23167 15011
rect 24394 15008 24400 15020
rect 23155 14980 24400 15008
rect 23155 14977 23167 14980
rect 23109 14971 23167 14977
rect 24394 14968 24400 14980
rect 24452 15008 24458 15020
rect 24949 15011 25007 15017
rect 24949 15008 24961 15011
rect 24452 14980 24961 15008
rect 24452 14968 24458 14980
rect 24949 14977 24961 14980
rect 24995 14977 25007 15011
rect 24949 14971 25007 14977
rect 6270 14900 6276 14952
rect 6328 14940 6334 14952
rect 6549 14943 6607 14949
rect 6549 14940 6561 14943
rect 6328 14912 6561 14940
rect 6328 14900 6334 14912
rect 6549 14909 6561 14912
rect 6595 14909 6607 14943
rect 12250 14940 12256 14952
rect 12211 14912 12256 14940
rect 6549 14903 6607 14909
rect 12250 14900 12256 14912
rect 12308 14900 12314 14952
rect 16666 14900 16672 14952
rect 16724 14940 16730 14952
rect 17310 14940 17316 14952
rect 16724 14912 17316 14940
rect 16724 14900 16730 14912
rect 17310 14900 17316 14912
rect 17368 14940 17374 14952
rect 17405 14943 17463 14949
rect 17405 14940 17417 14943
rect 17368 14912 17417 14940
rect 17368 14900 17374 14912
rect 17405 14909 17417 14912
rect 17451 14909 17463 14943
rect 25056 14940 25084 15048
rect 25216 15045 25228 15079
rect 25262 15076 25274 15079
rect 27062 15076 27068 15088
rect 25262 15048 27068 15076
rect 25262 15045 25274 15048
rect 25216 15039 25274 15045
rect 27062 15036 27068 15048
rect 27120 15036 27126 15088
rect 27240 15079 27298 15085
rect 27240 15045 27252 15079
rect 27286 15076 27298 15079
rect 28166 15076 28172 15088
rect 27286 15048 28172 15076
rect 27286 15045 27298 15048
rect 27240 15039 27298 15045
rect 28166 15036 28172 15048
rect 28224 15036 28230 15088
rect 29080 15079 29138 15085
rect 29080 15045 29092 15079
rect 29126 15076 29138 15079
rect 33226 15076 33232 15088
rect 29126 15048 33232 15076
rect 29126 15045 29138 15048
rect 29080 15039 29138 15045
rect 33226 15036 33232 15048
rect 33284 15036 33290 15088
rect 34968 15079 35026 15085
rect 34968 15045 34980 15079
rect 35014 15076 35026 15079
rect 36078 15076 36084 15088
rect 35014 15048 36084 15076
rect 35014 15045 35026 15048
rect 34968 15039 35026 15045
rect 36078 15036 36084 15048
rect 36136 15036 36142 15088
rect 37734 15036 37740 15088
rect 37792 15036 37798 15088
rect 39206 15036 39212 15088
rect 39264 15076 39270 15088
rect 39730 15079 39788 15085
rect 39730 15076 39742 15079
rect 39264 15048 39742 15076
rect 39264 15036 39270 15048
rect 39730 15045 39742 15048
rect 39776 15045 39788 15079
rect 45554 15076 45560 15088
rect 39730 15039 39788 15045
rect 45020 15048 45560 15076
rect 26786 14968 26792 15020
rect 26844 15008 26850 15020
rect 26973 15011 27031 15017
rect 26973 15008 26985 15011
rect 26844 14980 26985 15008
rect 26844 14968 26850 14980
rect 26973 14977 26985 14980
rect 27019 14977 27031 15011
rect 26973 14971 27031 14977
rect 33128 15011 33186 15017
rect 33128 14977 33140 15011
rect 33174 15008 33186 15011
rect 34514 15008 34520 15020
rect 33174 14980 34520 15008
rect 33174 14977 33186 14980
rect 33128 14971 33186 14977
rect 34514 14968 34520 14980
rect 34572 14968 34578 15020
rect 34606 14968 34612 15020
rect 34664 15008 34670 15020
rect 34701 15011 34759 15017
rect 34701 15008 34713 15011
rect 34664 14980 34713 15008
rect 34664 14968 34670 14980
rect 34701 14977 34713 14980
rect 34747 14977 34759 15011
rect 37550 15008 37556 15020
rect 37463 14980 37556 15008
rect 34701 14971 34759 14977
rect 37550 14968 37556 14980
rect 37608 15008 37614 15020
rect 37752 15008 37780 15036
rect 37608 14980 37780 15008
rect 37820 15011 37878 15017
rect 37608 14968 37614 14980
rect 37820 14977 37832 15011
rect 37866 15008 37878 15011
rect 38930 15008 38936 15020
rect 37866 14980 38936 15008
rect 37866 14977 37878 14980
rect 37820 14971 37878 14977
rect 38930 14968 38936 14980
rect 38988 14968 38994 15020
rect 39485 15011 39543 15017
rect 39485 14977 39497 15011
rect 39531 15008 39543 15011
rect 40034 15008 40040 15020
rect 39531 14980 40040 15008
rect 39531 14977 39543 14980
rect 39485 14971 39543 14977
rect 40034 14968 40040 14980
rect 40092 14968 40098 15020
rect 45020 15017 45048 15048
rect 45554 15036 45560 15048
rect 45612 15036 45618 15088
rect 47940 15079 47998 15085
rect 47940 15045 47952 15079
rect 47986 15076 47998 15079
rect 49050 15076 49056 15088
rect 47986 15048 49056 15076
rect 47986 15045 47998 15048
rect 47940 15039 47998 15045
rect 49050 15036 49056 15048
rect 49108 15036 49114 15088
rect 52748 15048 54984 15076
rect 45005 15011 45063 15017
rect 45005 14977 45017 15011
rect 45051 14977 45063 15011
rect 45005 14971 45063 14977
rect 45272 15011 45330 15017
rect 45272 14977 45284 15011
rect 45318 15008 45330 15011
rect 46658 15008 46664 15020
rect 45318 14980 46664 15008
rect 45318 14977 45330 14980
rect 45272 14971 45330 14977
rect 46658 14968 46664 14980
rect 46716 14968 46722 15020
rect 49142 14968 49148 15020
rect 49200 15008 49206 15020
rect 49769 15011 49827 15017
rect 49769 15008 49781 15011
rect 49200 14980 49781 15008
rect 49200 14968 49206 14980
rect 49769 14977 49781 14980
rect 49815 14977 49827 15011
rect 49769 14971 49827 14977
rect 51994 14968 52000 15020
rect 52052 15008 52058 15020
rect 52748 15017 52776 15048
rect 52733 15011 52791 15017
rect 52733 15008 52745 15011
rect 52052 14980 52745 15008
rect 52052 14968 52058 14980
rect 52733 14977 52745 14980
rect 52779 14977 52791 15011
rect 52733 14971 52791 14977
rect 53000 15011 53058 15017
rect 53000 14977 53012 15011
rect 53046 15008 53058 15011
rect 54846 15008 54852 15020
rect 53046 14980 54852 15008
rect 53046 14977 53058 14980
rect 53000 14971 53058 14977
rect 54846 14968 54852 14980
rect 54904 14968 54910 15020
rect 54956 14952 54984 15048
rect 56220 15011 56278 15017
rect 56220 14977 56232 15011
rect 56266 15008 56278 15011
rect 57330 15008 57336 15020
rect 56266 14980 57336 15008
rect 56266 14977 56278 14980
rect 56220 14971 56278 14977
rect 57330 14968 57336 14980
rect 57388 14968 57394 15020
rect 28810 14940 28816 14952
rect 17405 14903 17463 14909
rect 24964 14912 25084 14940
rect 28771 14912 28816 14940
rect 3050 14804 3056 14816
rect 3011 14776 3056 14804
rect 3050 14764 3056 14776
rect 3108 14764 3114 14816
rect 9674 14764 9680 14816
rect 9732 14804 9738 14816
rect 9861 14807 9919 14813
rect 9861 14804 9873 14807
rect 9732 14776 9873 14804
rect 9732 14764 9738 14776
rect 9861 14773 9873 14776
rect 9907 14773 9919 14807
rect 13630 14804 13636 14816
rect 13591 14776 13636 14804
rect 9861 14767 9919 14773
rect 13630 14764 13636 14776
rect 13688 14764 13694 14816
rect 15654 14804 15660 14816
rect 15615 14776 15660 14804
rect 15654 14764 15660 14776
rect 15712 14764 15718 14816
rect 24486 14804 24492 14816
rect 24447 14776 24492 14804
rect 24486 14764 24492 14776
rect 24544 14764 24550 14816
rect 24964 14804 24992 14912
rect 28810 14900 28816 14912
rect 28868 14900 28874 14952
rect 32858 14940 32864 14952
rect 32819 14912 32864 14940
rect 32858 14900 32864 14912
rect 32916 14900 32922 14952
rect 47578 14900 47584 14952
rect 47636 14940 47642 14952
rect 47673 14943 47731 14949
rect 47673 14940 47685 14943
rect 47636 14912 47685 14940
rect 47636 14900 47642 14912
rect 47673 14909 47685 14912
rect 47719 14909 47731 14943
rect 49510 14940 49516 14952
rect 49471 14912 49516 14940
rect 47673 14903 47731 14909
rect 49510 14900 49516 14912
rect 49568 14900 49574 14952
rect 54938 14900 54944 14952
rect 54996 14940 55002 14952
rect 55953 14943 56011 14949
rect 55953 14940 55965 14943
rect 54996 14912 55965 14940
rect 54996 14900 55002 14912
rect 55953 14909 55965 14912
rect 55999 14909 56011 14943
rect 55953 14903 56011 14909
rect 26694 14804 26700 14816
rect 24964 14776 26700 14804
rect 26694 14764 26700 14776
rect 26752 14764 26758 14816
rect 28350 14804 28356 14816
rect 28311 14776 28356 14804
rect 28350 14764 28356 14776
rect 28408 14764 28414 14816
rect 30190 14804 30196 14816
rect 30151 14776 30196 14804
rect 30190 14764 30196 14776
rect 30248 14764 30254 14816
rect 34241 14807 34299 14813
rect 34241 14773 34253 14807
rect 34287 14804 34299 14807
rect 34698 14804 34704 14816
rect 34287 14776 34704 14804
rect 34287 14773 34299 14776
rect 34241 14767 34299 14773
rect 34698 14764 34704 14776
rect 34756 14764 34762 14816
rect 36078 14804 36084 14816
rect 36039 14776 36084 14804
rect 36078 14764 36084 14776
rect 36136 14764 36142 14816
rect 49050 14804 49056 14816
rect 49011 14776 49056 14804
rect 49050 14764 49056 14776
rect 49108 14764 49114 14816
rect 49786 14764 49792 14816
rect 49844 14804 49850 14816
rect 50893 14807 50951 14813
rect 50893 14804 50905 14807
rect 49844 14776 50905 14804
rect 49844 14764 49850 14776
rect 50893 14773 50905 14776
rect 50939 14773 50951 14807
rect 50893 14767 50951 14773
rect 53650 14764 53656 14816
rect 53708 14804 53714 14816
rect 54113 14807 54171 14813
rect 54113 14804 54125 14807
rect 53708 14776 54125 14804
rect 53708 14764 53714 14776
rect 54113 14773 54125 14776
rect 54159 14773 54171 14807
rect 54113 14767 54171 14773
rect 1104 14714 59340 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 59340 14714
rect 1104 14640 59340 14662
rect 8110 14600 8116 14612
rect 8071 14572 8116 14600
rect 8110 14560 8116 14572
rect 8168 14560 8174 14612
rect 18506 14600 18512 14612
rect 18467 14572 18512 14600
rect 18506 14560 18512 14572
rect 18564 14560 18570 14612
rect 23658 14600 23664 14612
rect 23619 14572 23664 14600
rect 23658 14560 23664 14572
rect 23716 14560 23722 14612
rect 31846 14600 31852 14612
rect 31807 14572 31852 14600
rect 31846 14560 31852 14572
rect 31904 14560 31910 14612
rect 41233 14603 41291 14609
rect 41233 14569 41245 14603
rect 41279 14600 41291 14603
rect 41598 14600 41604 14612
rect 41279 14572 41604 14600
rect 41279 14569 41291 14572
rect 41233 14563 41291 14569
rect 41598 14560 41604 14572
rect 41656 14560 41662 14612
rect 46658 14600 46664 14612
rect 46619 14572 46664 14600
rect 46658 14560 46664 14572
rect 46716 14560 46722 14612
rect 19150 14424 19156 14476
rect 19208 14464 19214 14476
rect 20441 14467 20499 14473
rect 20441 14464 20453 14467
rect 19208 14436 20453 14464
rect 19208 14424 19214 14436
rect 20441 14433 20453 14436
rect 20487 14433 20499 14467
rect 20441 14427 20499 14433
rect 32858 14424 32864 14476
rect 32916 14464 32922 14476
rect 34057 14467 34115 14473
rect 34057 14464 34069 14467
rect 32916 14436 34069 14464
rect 32916 14424 32922 14436
rect 34057 14433 34069 14436
rect 34103 14464 34115 14467
rect 34606 14464 34612 14476
rect 34103 14436 34612 14464
rect 34103 14433 34115 14436
rect 34057 14427 34115 14433
rect 34606 14424 34612 14436
rect 34664 14424 34670 14476
rect 34790 14424 34796 14476
rect 34848 14464 34854 14476
rect 34885 14467 34943 14473
rect 34885 14464 34897 14467
rect 34848 14436 34897 14464
rect 34848 14424 34854 14436
rect 34885 14433 34897 14436
rect 34931 14433 34943 14467
rect 34885 14427 34943 14433
rect 39301 14467 39359 14473
rect 39301 14433 39313 14467
rect 39347 14464 39359 14467
rect 39758 14464 39764 14476
rect 39347 14436 39764 14464
rect 39347 14433 39359 14436
rect 39301 14427 39359 14433
rect 39758 14424 39764 14436
rect 39816 14464 39822 14476
rect 39853 14467 39911 14473
rect 39853 14464 39865 14467
rect 39816 14436 39865 14464
rect 39816 14424 39822 14436
rect 39853 14433 39865 14436
rect 39899 14433 39911 14467
rect 39853 14427 39911 14433
rect 45002 14424 45008 14476
rect 45060 14464 45066 14476
rect 45281 14467 45339 14473
rect 45281 14464 45293 14467
rect 45060 14436 45293 14464
rect 45060 14424 45066 14436
rect 45281 14433 45293 14436
rect 45327 14433 45339 14467
rect 51994 14464 52000 14476
rect 51955 14436 52000 14464
rect 45281 14427 45339 14433
rect 51994 14424 52000 14436
rect 52052 14424 52058 14476
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 1762 14396 1768 14408
rect 1719 14368 1768 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 1762 14356 1768 14368
rect 1820 14356 1826 14408
rect 1940 14399 1998 14405
rect 1940 14365 1952 14399
rect 1986 14396 1998 14399
rect 3050 14396 3056 14408
rect 1986 14368 3056 14396
rect 1986 14365 1998 14368
rect 1940 14359 1998 14365
rect 3050 14356 3056 14368
rect 3108 14356 3114 14408
rect 6270 14356 6276 14408
rect 6328 14396 6334 14408
rect 6733 14399 6791 14405
rect 6733 14396 6745 14399
rect 6328 14368 6745 14396
rect 6328 14356 6334 14368
rect 6733 14365 6745 14368
rect 6779 14365 6791 14399
rect 9861 14399 9919 14405
rect 9861 14396 9873 14399
rect 6733 14359 6791 14365
rect 6886 14368 9873 14396
rect 4525 14331 4583 14337
rect 4525 14297 4537 14331
rect 4571 14328 4583 14331
rect 6886 14328 6914 14368
rect 9861 14365 9873 14368
rect 9907 14396 9919 14399
rect 11054 14396 11060 14408
rect 9907 14368 11060 14396
rect 9907 14365 9919 14368
rect 9861 14359 9919 14365
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 12161 14399 12219 14405
rect 12161 14396 12173 14399
rect 11164 14368 12173 14396
rect 4571 14300 6914 14328
rect 7000 14331 7058 14337
rect 4571 14297 4583 14300
rect 4525 14291 4583 14297
rect 7000 14297 7012 14331
rect 7046 14328 7058 14331
rect 7926 14328 7932 14340
rect 7046 14300 7932 14328
rect 7046 14297 7058 14300
rect 7000 14291 7058 14297
rect 7926 14288 7932 14300
rect 7984 14288 7990 14340
rect 3050 14260 3056 14272
rect 3011 14232 3056 14260
rect 3050 14220 3056 14232
rect 3108 14220 3114 14272
rect 5534 14220 5540 14272
rect 5592 14260 5598 14272
rect 5813 14263 5871 14269
rect 5813 14260 5825 14263
rect 5592 14232 5825 14260
rect 5592 14220 5598 14232
rect 5813 14229 5825 14232
rect 5859 14229 5871 14263
rect 5813 14223 5871 14229
rect 10778 14220 10784 14272
rect 10836 14260 10842 14272
rect 11164 14269 11192 14368
rect 12161 14365 12173 14368
rect 12207 14396 12219 14399
rect 12250 14396 12256 14408
rect 12207 14368 12256 14396
rect 12207 14365 12219 14368
rect 12161 14359 12219 14365
rect 12250 14356 12256 14368
rect 12308 14356 12314 14408
rect 14093 14399 14151 14405
rect 14093 14365 14105 14399
rect 14139 14396 14151 14399
rect 14182 14396 14188 14408
rect 14139 14368 14188 14396
rect 14139 14365 14151 14368
rect 14093 14359 14151 14365
rect 14182 14356 14188 14368
rect 14240 14356 14246 14408
rect 14360 14399 14418 14405
rect 14360 14365 14372 14399
rect 14406 14396 14418 14399
rect 15654 14396 15660 14408
rect 14406 14368 15660 14396
rect 14406 14365 14418 14368
rect 14360 14359 14418 14365
rect 15654 14356 15660 14368
rect 15712 14356 15718 14408
rect 16758 14356 16764 14408
rect 16816 14396 16822 14408
rect 17129 14399 17187 14405
rect 17129 14396 17141 14399
rect 16816 14368 17141 14396
rect 16816 14356 16822 14368
rect 17129 14365 17141 14368
rect 17175 14365 17187 14399
rect 22281 14399 22339 14405
rect 17129 14359 17187 14365
rect 20640 14368 22232 14396
rect 12428 14331 12486 14337
rect 12428 14297 12440 14331
rect 12474 14328 12486 14331
rect 14550 14328 14556 14340
rect 12474 14300 14556 14328
rect 12474 14297 12486 14300
rect 12428 14291 12486 14297
rect 14550 14288 14556 14300
rect 14608 14288 14614 14340
rect 17396 14331 17454 14337
rect 17396 14297 17408 14331
rect 17442 14328 17454 14331
rect 20640 14328 20668 14368
rect 17442 14300 20668 14328
rect 20708 14331 20766 14337
rect 17442 14297 17454 14300
rect 17396 14291 17454 14297
rect 20708 14297 20720 14331
rect 20754 14328 20766 14331
rect 21266 14328 21272 14340
rect 20754 14300 21272 14328
rect 20754 14297 20766 14300
rect 20708 14291 20766 14297
rect 21266 14288 21272 14300
rect 21324 14288 21330 14340
rect 22204 14328 22232 14368
rect 22281 14365 22293 14399
rect 22327 14396 22339 14399
rect 24394 14396 24400 14408
rect 22327 14368 24400 14396
rect 22327 14365 22339 14368
rect 22281 14359 22339 14365
rect 24394 14356 24400 14368
rect 24452 14356 24458 14408
rect 28810 14356 28816 14408
rect 28868 14396 28874 14408
rect 30469 14399 30527 14405
rect 30469 14396 30481 14399
rect 28868 14368 30481 14396
rect 28868 14356 28874 14368
rect 30469 14365 30481 14368
rect 30515 14365 30527 14399
rect 30469 14359 30527 14365
rect 30736 14399 30794 14405
rect 30736 14365 30748 14399
rect 30782 14396 30794 14399
rect 32122 14396 32128 14408
rect 30782 14368 32128 14396
rect 30782 14365 30794 14368
rect 30736 14359 30794 14365
rect 22370 14328 22376 14340
rect 22204 14300 22376 14328
rect 22370 14288 22376 14300
rect 22428 14288 22434 14340
rect 22548 14331 22606 14337
rect 22548 14297 22560 14331
rect 22594 14328 22606 14331
rect 23198 14328 23204 14340
rect 22594 14300 23204 14328
rect 22594 14297 22606 14300
rect 22548 14291 22606 14297
rect 23198 14288 23204 14300
rect 23256 14288 23262 14340
rect 25961 14331 26019 14337
rect 25961 14297 25973 14331
rect 26007 14328 26019 14331
rect 26234 14328 26240 14340
rect 26007 14300 26240 14328
rect 26007 14297 26019 14300
rect 25961 14291 26019 14297
rect 26234 14288 26240 14300
rect 26292 14288 26298 14340
rect 27522 14328 27528 14340
rect 27483 14300 27528 14328
rect 27522 14288 27528 14300
rect 27580 14288 27586 14340
rect 11149 14263 11207 14269
rect 11149 14260 11161 14263
rect 10836 14232 11161 14260
rect 10836 14220 10842 14232
rect 11149 14229 11161 14232
rect 11195 14229 11207 14263
rect 11149 14223 11207 14229
rect 13541 14263 13599 14269
rect 13541 14229 13553 14263
rect 13587 14260 13599 14263
rect 14182 14260 14188 14272
rect 13587 14232 14188 14260
rect 13587 14229 13599 14232
rect 13541 14223 13599 14229
rect 14182 14220 14188 14232
rect 14240 14220 14246 14272
rect 15470 14260 15476 14272
rect 15431 14232 15476 14260
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 21818 14260 21824 14272
rect 21779 14232 21824 14260
rect 21818 14220 21824 14232
rect 21876 14220 21882 14272
rect 30484 14260 30512 14359
rect 32122 14356 32128 14368
rect 32180 14356 32186 14408
rect 35152 14399 35210 14405
rect 35152 14365 35164 14399
rect 35198 14396 35210 14399
rect 36078 14396 36084 14408
rect 35198 14368 36084 14396
rect 35198 14365 35210 14368
rect 35152 14359 35210 14365
rect 36078 14356 36084 14368
rect 36136 14356 36142 14408
rect 40120 14399 40178 14405
rect 40120 14365 40132 14399
rect 40166 14396 40178 14399
rect 41506 14396 41512 14408
rect 40166 14368 41512 14396
rect 40166 14365 40178 14368
rect 40120 14359 40178 14365
rect 41506 14356 41512 14368
rect 41564 14356 41570 14408
rect 47578 14396 47584 14408
rect 47539 14368 47584 14396
rect 47578 14356 47584 14368
rect 47636 14356 47642 14408
rect 47848 14399 47906 14405
rect 47848 14365 47860 14399
rect 47894 14396 47906 14399
rect 49050 14396 49056 14408
rect 47894 14368 49056 14396
rect 47894 14365 47906 14368
rect 47848 14359 47906 14365
rect 49050 14356 49056 14368
rect 49108 14356 49114 14408
rect 50157 14399 50215 14405
rect 50157 14365 50169 14399
rect 50203 14396 50215 14399
rect 52012 14396 52040 14424
rect 50203 14368 52040 14396
rect 50203 14365 50215 14368
rect 50157 14359 50215 14365
rect 52086 14356 52092 14408
rect 52144 14396 52150 14408
rect 52253 14399 52311 14405
rect 52253 14396 52265 14399
rect 52144 14368 52265 14396
rect 52144 14356 52150 14368
rect 52253 14365 52265 14368
rect 52299 14365 52311 14399
rect 52253 14359 52311 14365
rect 55950 14356 55956 14408
rect 56008 14396 56014 14408
rect 56410 14396 56416 14408
rect 56008 14368 56416 14396
rect 56008 14356 56014 14368
rect 56410 14356 56416 14368
rect 56468 14396 56474 14408
rect 56689 14399 56747 14405
rect 56689 14396 56701 14399
rect 56468 14368 56701 14396
rect 56468 14356 56474 14368
rect 56689 14365 56701 14368
rect 56735 14365 56747 14399
rect 56689 14359 56747 14365
rect 32306 14328 32312 14340
rect 32267 14300 32312 14328
rect 32306 14288 32312 14300
rect 32364 14328 32370 14340
rect 37553 14331 37611 14337
rect 37553 14328 37565 14331
rect 32364 14300 37565 14328
rect 32364 14288 32370 14300
rect 37553 14297 37565 14300
rect 37599 14328 37611 14331
rect 39850 14328 39856 14340
rect 37599 14300 39856 14328
rect 37599 14297 37611 14300
rect 37553 14291 37611 14297
rect 39850 14288 39856 14300
rect 39908 14288 39914 14340
rect 45548 14331 45606 14337
rect 45548 14297 45560 14331
rect 45594 14328 45606 14331
rect 46382 14328 46388 14340
rect 45594 14300 46388 14328
rect 45594 14297 45606 14300
rect 45548 14291 45606 14297
rect 46382 14288 46388 14300
rect 46440 14288 46446 14340
rect 49694 14288 49700 14340
rect 49752 14328 49758 14340
rect 50402 14331 50460 14337
rect 50402 14328 50414 14331
rect 49752 14300 50414 14328
rect 49752 14288 49758 14300
rect 50402 14297 50414 14300
rect 50448 14297 50460 14331
rect 50402 14291 50460 14297
rect 55582 14288 55588 14340
rect 55640 14328 55646 14340
rect 56934 14331 56992 14337
rect 56934 14328 56946 14331
rect 55640 14300 56946 14328
rect 55640 14288 55646 14300
rect 56934 14297 56946 14300
rect 56980 14297 56992 14331
rect 56934 14291 56992 14297
rect 32858 14260 32864 14272
rect 30484 14232 32864 14260
rect 32858 14220 32864 14232
rect 32916 14220 32922 14272
rect 36262 14260 36268 14272
rect 36223 14232 36268 14260
rect 36262 14220 36268 14232
rect 36320 14220 36326 14272
rect 48958 14260 48964 14272
rect 48919 14232 48964 14260
rect 48958 14220 48964 14232
rect 49016 14220 49022 14272
rect 51534 14260 51540 14272
rect 51495 14232 51540 14260
rect 51534 14220 51540 14232
rect 51592 14220 51598 14272
rect 53374 14260 53380 14272
rect 53335 14232 53380 14260
rect 53374 14220 53380 14232
rect 53432 14220 53438 14272
rect 58066 14260 58072 14272
rect 58027 14232 58072 14260
rect 58066 14220 58072 14232
rect 58124 14220 58130 14272
rect 1104 14170 59340 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 59340 14170
rect 1104 14096 59340 14118
rect 7926 14056 7932 14068
rect 7887 14028 7932 14056
rect 7926 14016 7932 14028
rect 7984 14016 7990 14068
rect 12897 14059 12955 14065
rect 12897 14025 12909 14059
rect 12943 14025 12955 14059
rect 12897 14019 12955 14025
rect 18049 14059 18107 14065
rect 18049 14025 18061 14059
rect 18095 14025 18107 14059
rect 18049 14019 18107 14025
rect 21269 14059 21327 14065
rect 21269 14025 21281 14059
rect 21315 14056 21327 14059
rect 23198 14056 23204 14068
rect 21315 14028 21956 14056
rect 23159 14028 23204 14056
rect 21315 14025 21327 14028
rect 21269 14019 21327 14025
rect 1940 13991 1998 13997
rect 1940 13957 1952 13991
rect 1986 13988 1998 13991
rect 3050 13988 3056 14000
rect 1986 13960 3056 13988
rect 1986 13957 1998 13960
rect 1940 13951 1998 13957
rect 3050 13948 3056 13960
rect 3108 13948 3114 14000
rect 9852 13991 9910 13997
rect 9852 13957 9864 13991
rect 9898 13988 9910 13991
rect 12912 13988 12940 14019
rect 9898 13960 12940 13988
rect 14360 13991 14418 13997
rect 9898 13957 9910 13960
rect 9852 13951 9910 13957
rect 14360 13957 14372 13991
rect 14406 13988 14418 13991
rect 15470 13988 15476 14000
rect 14406 13960 15476 13988
rect 14406 13957 14418 13960
rect 14360 13951 14418 13957
rect 15470 13948 15476 13960
rect 15528 13948 15534 14000
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13920 1731 13923
rect 1762 13920 1768 13932
rect 1719 13892 1768 13920
rect 1719 13889 1731 13892
rect 1673 13883 1731 13889
rect 1762 13880 1768 13892
rect 1820 13880 1826 13932
rect 6816 13923 6874 13929
rect 6816 13889 6828 13923
rect 6862 13920 6874 13923
rect 8202 13920 8208 13932
rect 6862 13892 8208 13920
rect 6862 13889 6874 13892
rect 6816 13883 6874 13889
rect 8202 13880 8208 13892
rect 8260 13880 8266 13932
rect 11784 13923 11842 13929
rect 11784 13889 11796 13923
rect 11830 13920 11842 13923
rect 13630 13920 13636 13932
rect 11830 13892 13636 13920
rect 11830 13889 11842 13892
rect 11784 13883 11842 13889
rect 13630 13880 13636 13892
rect 13688 13880 13694 13932
rect 14090 13920 14096 13932
rect 14051 13892 14096 13920
rect 14090 13880 14096 13892
rect 14148 13880 14154 13932
rect 16669 13923 16727 13929
rect 16669 13889 16681 13923
rect 16715 13920 16727 13923
rect 16758 13920 16764 13932
rect 16715 13892 16764 13920
rect 16715 13889 16727 13892
rect 16669 13883 16727 13889
rect 16758 13880 16764 13892
rect 16816 13880 16822 13932
rect 16936 13923 16994 13929
rect 16936 13889 16948 13923
rect 16982 13920 16994 13923
rect 18064 13920 18092 14019
rect 20156 13991 20214 13997
rect 20156 13957 20168 13991
rect 20202 13988 20214 13991
rect 21818 13988 21824 14000
rect 20202 13960 21824 13988
rect 20202 13957 20214 13960
rect 20156 13951 20214 13957
rect 21818 13948 21824 13960
rect 21876 13948 21882 14000
rect 21928 13988 21956 14028
rect 23198 14016 23204 14028
rect 23256 14016 23262 14068
rect 30190 14056 30196 14068
rect 26206 14028 30196 14056
rect 22066 13991 22124 13997
rect 22066 13988 22078 13991
rect 21928 13960 22078 13988
rect 22066 13957 22078 13960
rect 22112 13957 22124 13991
rect 22066 13951 22124 13957
rect 22186 13948 22192 14000
rect 22244 13948 22250 14000
rect 25308 13991 25366 13997
rect 25308 13957 25320 13991
rect 25354 13988 25366 13991
rect 26206 13988 26234 14028
rect 30190 14016 30196 14028
rect 30248 14016 30254 14068
rect 33962 14016 33968 14068
rect 34020 14056 34026 14068
rect 34149 14059 34207 14065
rect 34149 14056 34161 14059
rect 34020 14028 34161 14056
rect 34020 14016 34026 14028
rect 34149 14025 34161 14028
rect 34195 14025 34207 14059
rect 38930 14056 38936 14068
rect 38891 14028 38936 14056
rect 34149 14019 34207 14025
rect 38930 14016 38936 14028
rect 38988 14016 38994 14068
rect 44542 14016 44548 14068
rect 44600 14056 44606 14068
rect 46109 14059 46167 14065
rect 46109 14056 46121 14059
rect 44600 14028 46121 14056
rect 44600 14016 44606 14028
rect 46109 14025 46121 14028
rect 46155 14025 46167 14059
rect 46109 14019 46167 14025
rect 49053 14059 49111 14065
rect 49053 14025 49065 14059
rect 49099 14056 49111 14059
rect 49142 14056 49148 14068
rect 49099 14028 49148 14056
rect 49099 14025 49111 14028
rect 49053 14019 49111 14025
rect 49142 14016 49148 14028
rect 49200 14016 49206 14068
rect 56686 14056 56692 14068
rect 55186 14028 56692 14056
rect 25354 13960 26234 13988
rect 27240 13991 27298 13997
rect 25354 13957 25366 13960
rect 25308 13951 25366 13957
rect 27240 13957 27252 13991
rect 27286 13988 27298 13991
rect 28350 13988 28356 14000
rect 27286 13960 28356 13988
rect 27286 13957 27298 13960
rect 27240 13951 27298 13957
rect 28350 13948 28356 13960
rect 28408 13948 28414 14000
rect 33036 13991 33094 13997
rect 33036 13957 33048 13991
rect 33082 13988 33094 13991
rect 35244 13991 35302 13997
rect 33082 13960 35204 13988
rect 33082 13957 33094 13960
rect 33036 13951 33094 13957
rect 22204 13920 22232 13948
rect 16982 13892 18000 13920
rect 18064 13892 22232 13920
rect 16982 13889 16994 13892
rect 16936 13883 16994 13889
rect 6270 13812 6276 13864
rect 6328 13852 6334 13864
rect 6549 13855 6607 13861
rect 6549 13852 6561 13855
rect 6328 13824 6561 13852
rect 6328 13812 6334 13824
rect 6549 13821 6561 13824
rect 6595 13821 6607 13855
rect 6549 13815 6607 13821
rect 9585 13855 9643 13861
rect 9585 13821 9597 13855
rect 9631 13821 9643 13855
rect 9585 13815 9643 13821
rect 3050 13716 3056 13728
rect 3011 13688 3056 13716
rect 3050 13676 3056 13688
rect 3108 13676 3114 13728
rect 9600 13716 9628 13815
rect 10778 13812 10784 13864
rect 10836 13852 10842 13864
rect 11517 13855 11575 13861
rect 11517 13852 11529 13855
rect 10836 13824 11529 13852
rect 10836 13812 10842 13824
rect 11517 13821 11529 13824
rect 11563 13821 11575 13855
rect 17972 13852 18000 13892
rect 24394 13880 24400 13932
rect 24452 13920 24458 13932
rect 25041 13923 25099 13929
rect 25041 13920 25053 13923
rect 24452 13892 25053 13920
rect 24452 13880 24458 13892
rect 25041 13889 25053 13892
rect 25087 13920 25099 13923
rect 26973 13923 27031 13929
rect 26973 13920 26985 13923
rect 25087 13892 26985 13920
rect 25087 13889 25099 13892
rect 25041 13883 25099 13889
rect 26973 13889 26985 13892
rect 27019 13920 27031 13923
rect 27062 13920 27068 13932
rect 27019 13892 27068 13920
rect 27019 13889 27031 13892
rect 26973 13883 27031 13889
rect 27062 13880 27068 13892
rect 27120 13920 27126 13932
rect 27522 13920 27528 13932
rect 27120 13892 27528 13920
rect 27120 13880 27126 13892
rect 27522 13880 27528 13892
rect 27580 13920 27586 13932
rect 29086 13929 29092 13932
rect 28813 13923 28871 13929
rect 28813 13920 28825 13923
rect 27580 13892 28825 13920
rect 27580 13880 27586 13892
rect 28813 13889 28825 13892
rect 28859 13889 28871 13923
rect 28813 13883 28871 13889
rect 29080 13883 29092 13929
rect 29144 13920 29150 13932
rect 32769 13923 32827 13929
rect 29144 13892 29180 13920
rect 29086 13880 29092 13883
rect 29144 13880 29150 13892
rect 32769 13889 32781 13923
rect 32815 13920 32827 13923
rect 32858 13920 32864 13932
rect 32815 13892 32864 13920
rect 32815 13889 32827 13892
rect 32769 13883 32827 13889
rect 32858 13880 32864 13892
rect 32916 13880 32922 13932
rect 34790 13880 34796 13932
rect 34848 13920 34854 13932
rect 34977 13923 35035 13929
rect 34977 13920 34989 13923
rect 34848 13892 34989 13920
rect 34848 13880 34854 13892
rect 34977 13889 34989 13892
rect 35023 13889 35035 13923
rect 35176 13920 35204 13960
rect 35244 13957 35256 13991
rect 35290 13988 35302 13991
rect 36262 13988 36268 14000
rect 35290 13960 36268 13988
rect 35290 13957 35302 13960
rect 35244 13951 35302 13957
rect 36262 13948 36268 13960
rect 36320 13948 36326 14000
rect 44910 13988 44916 14000
rect 42904 13960 44916 13988
rect 36078 13920 36084 13932
rect 35176 13892 36084 13920
rect 34977 13883 35035 13889
rect 36078 13880 36084 13892
rect 36136 13880 36142 13932
rect 37550 13920 37556 13932
rect 37511 13892 37556 13920
rect 37550 13880 37556 13892
rect 37608 13880 37614 13932
rect 37820 13923 37878 13929
rect 37820 13889 37832 13923
rect 37866 13920 37878 13923
rect 38930 13920 38936 13932
rect 37866 13892 38936 13920
rect 37866 13889 37878 13892
rect 37820 13883 37878 13889
rect 38930 13880 38936 13892
rect 38988 13880 38994 13932
rect 18230 13852 18236 13864
rect 17972 13824 18236 13852
rect 11517 13815 11575 13821
rect 18230 13812 18236 13824
rect 18288 13812 18294 13864
rect 19150 13812 19156 13864
rect 19208 13852 19214 13864
rect 42904 13861 42932 13960
rect 42978 13880 42984 13932
rect 43036 13920 43042 13932
rect 44744 13929 44772 13960
rect 44910 13948 44916 13960
rect 44968 13948 44974 14000
rect 47940 13991 47998 13997
rect 47940 13957 47952 13991
rect 47986 13988 47998 13991
rect 48958 13988 48964 14000
rect 47986 13960 48964 13988
rect 47986 13957 47998 13960
rect 47940 13951 47998 13957
rect 48958 13948 48964 13960
rect 49016 13948 49022 14000
rect 50056 13991 50114 13997
rect 50056 13957 50068 13991
rect 50102 13988 50114 13991
rect 51534 13988 51540 14000
rect 50102 13960 51540 13988
rect 50102 13957 50114 13960
rect 50056 13951 50114 13957
rect 51534 13948 51540 13960
rect 51592 13948 51598 14000
rect 54849 13991 54907 13997
rect 54849 13957 54861 13991
rect 54895 13988 54907 13991
rect 54938 13988 54944 14000
rect 54895 13960 54944 13988
rect 54895 13957 54907 13960
rect 54849 13951 54907 13957
rect 54938 13948 54944 13960
rect 54996 13948 55002 14000
rect 43145 13923 43203 13929
rect 43145 13920 43157 13923
rect 43036 13892 43157 13920
rect 43036 13880 43042 13892
rect 43145 13889 43157 13892
rect 43191 13889 43203 13923
rect 43145 13883 43203 13889
rect 44729 13923 44787 13929
rect 44729 13889 44741 13923
rect 44775 13889 44787 13923
rect 44729 13883 44787 13889
rect 44996 13923 45054 13929
rect 44996 13889 45008 13923
rect 45042 13920 45054 13923
rect 46750 13920 46756 13932
rect 45042 13892 46756 13920
rect 45042 13889 45054 13892
rect 44996 13883 45054 13889
rect 46750 13880 46756 13892
rect 46808 13880 46814 13932
rect 49510 13880 49516 13932
rect 49568 13920 49574 13932
rect 49789 13923 49847 13929
rect 49789 13920 49801 13923
rect 49568 13892 49801 13920
rect 49568 13880 49574 13892
rect 49789 13889 49801 13892
rect 49835 13889 49847 13923
rect 53098 13920 53104 13932
rect 53011 13892 53104 13920
rect 49789 13883 49847 13889
rect 53098 13880 53104 13892
rect 53156 13920 53162 13932
rect 55186 13920 55214 14028
rect 56686 14016 56692 14028
rect 56744 14016 56750 14068
rect 57330 14056 57336 14068
rect 57291 14028 57336 14056
rect 57330 14016 57336 14028
rect 57388 14016 57394 14068
rect 56220 13991 56278 13997
rect 56220 13957 56232 13991
rect 56266 13988 56278 13991
rect 58066 13988 58072 14000
rect 56266 13960 58072 13988
rect 56266 13957 56278 13960
rect 56220 13951 56278 13957
rect 58066 13948 58072 13960
rect 58124 13948 58130 14000
rect 53156 13892 55214 13920
rect 53156 13880 53162 13892
rect 19889 13855 19947 13861
rect 19889 13852 19901 13855
rect 19208 13824 19901 13852
rect 19208 13812 19214 13824
rect 19889 13821 19901 13824
rect 19935 13821 19947 13855
rect 19889 13815 19947 13821
rect 21821 13855 21879 13861
rect 21821 13821 21833 13855
rect 21867 13821 21879 13855
rect 21821 13815 21879 13821
rect 42889 13855 42947 13861
rect 42889 13821 42901 13855
rect 42935 13821 42947 13855
rect 42889 13815 42947 13821
rect 9766 13716 9772 13728
rect 9600 13688 9772 13716
rect 9766 13676 9772 13688
rect 9824 13676 9830 13728
rect 10965 13719 11023 13725
rect 10965 13685 10977 13719
rect 11011 13716 11023 13719
rect 11054 13716 11060 13728
rect 11011 13688 11060 13716
rect 11011 13685 11023 13688
rect 10965 13679 11023 13685
rect 11054 13676 11060 13688
rect 11112 13676 11118 13728
rect 15470 13716 15476 13728
rect 15431 13688 15476 13716
rect 15470 13676 15476 13688
rect 15528 13676 15534 13728
rect 19904 13716 19932 13815
rect 21836 13784 21864 13815
rect 47578 13812 47584 13864
rect 47636 13852 47642 13864
rect 47673 13855 47731 13861
rect 47673 13852 47685 13855
rect 47636 13824 47685 13852
rect 47636 13812 47642 13824
rect 47673 13821 47685 13824
rect 47719 13821 47731 13855
rect 55950 13852 55956 13864
rect 55911 13824 55956 13852
rect 47673 13815 47731 13821
rect 20824 13756 21864 13784
rect 20824 13728 20852 13756
rect 20806 13716 20812 13728
rect 19904 13688 20812 13716
rect 20806 13676 20812 13688
rect 20864 13676 20870 13728
rect 26418 13716 26424 13728
rect 26379 13688 26424 13716
rect 26418 13676 26424 13688
rect 26476 13676 26482 13728
rect 28350 13716 28356 13728
rect 28311 13688 28356 13716
rect 28350 13676 28356 13688
rect 28408 13676 28414 13728
rect 30190 13716 30196 13728
rect 30151 13688 30196 13716
rect 30190 13676 30196 13688
rect 30248 13676 30254 13728
rect 36354 13716 36360 13728
rect 36315 13688 36360 13716
rect 36354 13676 36360 13688
rect 36412 13676 36418 13728
rect 44266 13716 44272 13728
rect 44227 13688 44272 13716
rect 44266 13676 44272 13688
rect 44324 13676 44330 13728
rect 47688 13716 47716 13815
rect 55950 13812 55956 13824
rect 56008 13812 56014 13864
rect 47946 13716 47952 13728
rect 47688 13688 47952 13716
rect 47946 13676 47952 13688
rect 48004 13676 48010 13728
rect 51166 13716 51172 13728
rect 51127 13688 51172 13716
rect 51166 13676 51172 13688
rect 51224 13676 51230 13728
rect 1104 13626 59340 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 59340 13626
rect 1104 13552 59340 13574
rect 8202 13512 8208 13524
rect 8163 13484 8208 13512
rect 8202 13472 8208 13484
rect 8260 13472 8266 13524
rect 12158 13512 12164 13524
rect 12119 13484 12164 13512
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 26694 13512 26700 13524
rect 26655 13484 26700 13512
rect 26694 13472 26700 13484
rect 26752 13472 26758 13524
rect 34514 13472 34520 13524
rect 34572 13512 34578 13524
rect 36357 13515 36415 13521
rect 36357 13512 36369 13515
rect 34572 13484 36369 13512
rect 34572 13472 34578 13484
rect 36357 13481 36369 13484
rect 36403 13481 36415 13515
rect 38930 13512 38936 13524
rect 38891 13484 38936 13512
rect 36357 13475 36415 13481
rect 38930 13472 38936 13484
rect 38988 13472 38994 13524
rect 42797 13515 42855 13521
rect 42797 13481 42809 13515
rect 42843 13512 42855 13515
rect 42978 13512 42984 13524
rect 42843 13484 42984 13512
rect 42843 13481 42855 13484
rect 42797 13475 42855 13481
rect 42978 13472 42984 13484
rect 43036 13472 43042 13524
rect 46382 13512 46388 13524
rect 46343 13484 46388 13512
rect 46382 13472 46388 13484
rect 46440 13472 46446 13524
rect 49329 13515 49387 13521
rect 49329 13481 49341 13515
rect 49375 13512 49387 13515
rect 49694 13512 49700 13524
rect 49375 13484 49700 13512
rect 49375 13481 49387 13484
rect 49329 13475 49387 13481
rect 49694 13472 49700 13484
rect 49752 13472 49758 13524
rect 51442 13472 51448 13524
rect 51500 13512 51506 13524
rect 51537 13515 51595 13521
rect 51537 13512 51549 13515
rect 51500 13484 51549 13512
rect 51500 13472 51506 13484
rect 51537 13481 51549 13484
rect 51583 13481 51595 13515
rect 51537 13475 51595 13481
rect 53282 13472 53288 13524
rect 53340 13512 53346 13524
rect 53377 13515 53435 13521
rect 53377 13512 53389 13515
rect 53340 13484 53389 13512
rect 53340 13472 53346 13484
rect 53377 13481 53389 13484
rect 53423 13481 53435 13515
rect 53377 13475 53435 13481
rect 24394 13336 24400 13388
rect 24452 13376 24458 13388
rect 25317 13379 25375 13385
rect 25317 13376 25329 13379
rect 24452 13348 25329 13376
rect 24452 13336 24458 13348
rect 25317 13345 25329 13348
rect 25363 13345 25375 13379
rect 25317 13339 25375 13345
rect 27062 13336 27068 13388
rect 27120 13376 27126 13388
rect 27157 13379 27215 13385
rect 27157 13376 27169 13379
rect 27120 13348 27169 13376
rect 27120 13336 27126 13348
rect 27157 13345 27169 13348
rect 27203 13345 27215 13379
rect 27157 13339 27215 13345
rect 34790 13336 34796 13388
rect 34848 13376 34854 13388
rect 34977 13379 35035 13385
rect 34977 13376 34989 13379
rect 34848 13348 34989 13376
rect 34848 13336 34854 13348
rect 34977 13345 34989 13348
rect 35023 13345 35035 13379
rect 37550 13376 37556 13388
rect 37511 13348 37556 13376
rect 34977 13339 35035 13345
rect 1854 13308 1860 13320
rect 1815 13280 1860 13308
rect 1854 13268 1860 13280
rect 1912 13268 1918 13320
rect 2124 13311 2182 13317
rect 2124 13277 2136 13311
rect 2170 13308 2182 13311
rect 3050 13308 3056 13320
rect 2170 13280 3056 13308
rect 2170 13277 2182 13280
rect 2124 13271 2182 13277
rect 3050 13268 3056 13280
rect 3108 13268 3114 13320
rect 4985 13311 5043 13317
rect 4985 13277 4997 13311
rect 5031 13308 5043 13311
rect 5534 13308 5540 13320
rect 5031 13280 5540 13308
rect 5031 13277 5043 13280
rect 4985 13271 5043 13277
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 6270 13268 6276 13320
rect 6328 13308 6334 13320
rect 6825 13311 6883 13317
rect 6825 13308 6837 13311
rect 6328 13280 6837 13308
rect 6328 13268 6334 13280
rect 6825 13277 6837 13280
rect 6871 13308 6883 13311
rect 8941 13311 8999 13317
rect 8941 13308 8953 13311
rect 6871 13280 8953 13308
rect 6871 13277 6883 13280
rect 6825 13271 6883 13277
rect 8941 13277 8953 13280
rect 8987 13308 8999 13311
rect 9766 13308 9772 13320
rect 8987 13280 9772 13308
rect 8987 13277 8999 13280
rect 8941 13271 8999 13277
rect 9766 13268 9772 13280
rect 9824 13308 9830 13320
rect 10778 13308 10784 13320
rect 9824 13280 10784 13308
rect 9824 13268 9830 13280
rect 10778 13268 10784 13280
rect 10836 13268 10842 13320
rect 11054 13317 11060 13320
rect 11048 13308 11060 13317
rect 11015 13280 11060 13308
rect 11048 13271 11060 13280
rect 11054 13268 11060 13271
rect 11112 13268 11118 13320
rect 20717 13311 20775 13317
rect 20717 13277 20729 13311
rect 20763 13308 20775 13311
rect 20806 13308 20812 13320
rect 20763 13280 20812 13308
rect 20763 13277 20775 13280
rect 20717 13271 20775 13277
rect 20806 13268 20812 13280
rect 20864 13268 20870 13320
rect 25584 13311 25642 13317
rect 25584 13277 25596 13311
rect 25630 13308 25642 13311
rect 26418 13308 26424 13320
rect 25630 13280 26424 13308
rect 25630 13277 25642 13280
rect 25584 13271 25642 13277
rect 26418 13268 26424 13280
rect 26476 13268 26482 13320
rect 27424 13311 27482 13317
rect 27424 13277 27436 13311
rect 27470 13308 27482 13311
rect 28350 13308 28356 13320
rect 27470 13280 28356 13308
rect 27470 13277 27482 13280
rect 27424 13271 27482 13277
rect 28350 13268 28356 13280
rect 28408 13268 28414 13320
rect 30929 13311 30987 13317
rect 30929 13277 30941 13311
rect 30975 13308 30987 13311
rect 32769 13311 32827 13317
rect 32769 13308 32781 13311
rect 30975 13280 32781 13308
rect 30975 13277 30987 13280
rect 30929 13271 30987 13277
rect 32769 13277 32781 13280
rect 32815 13308 32827 13311
rect 32858 13308 32864 13320
rect 32815 13280 32864 13308
rect 32815 13277 32827 13280
rect 32769 13271 32827 13277
rect 32858 13268 32864 13280
rect 32916 13268 32922 13320
rect 5252 13243 5310 13249
rect 5252 13209 5264 13243
rect 5298 13240 5310 13243
rect 5810 13240 5816 13252
rect 5298 13212 5816 13240
rect 5298 13209 5310 13212
rect 5252 13203 5310 13209
rect 5810 13200 5816 13212
rect 5868 13200 5874 13252
rect 7092 13243 7150 13249
rect 7092 13209 7104 13243
rect 7138 13240 7150 13243
rect 7742 13240 7748 13252
rect 7138 13212 7748 13240
rect 7138 13209 7150 13212
rect 7092 13203 7150 13209
rect 7742 13200 7748 13212
rect 7800 13200 7806 13252
rect 9208 13243 9266 13249
rect 9208 13209 9220 13243
rect 9254 13240 9266 13243
rect 11790 13240 11796 13252
rect 9254 13212 11796 13240
rect 9254 13209 9266 13212
rect 9208 13203 9266 13209
rect 11790 13200 11796 13212
rect 11848 13200 11854 13252
rect 15286 13200 15292 13252
rect 15344 13240 15350 13252
rect 15565 13243 15623 13249
rect 15565 13240 15577 13243
rect 15344 13212 15577 13240
rect 15344 13200 15350 13212
rect 15565 13209 15577 13212
rect 15611 13209 15623 13243
rect 15565 13203 15623 13209
rect 20984 13243 21042 13249
rect 20984 13209 20996 13243
rect 21030 13240 21042 13243
rect 22278 13240 22284 13252
rect 21030 13212 22284 13240
rect 21030 13209 21042 13212
rect 20984 13203 21042 13209
rect 22278 13200 22284 13212
rect 22336 13200 22342 13252
rect 31196 13243 31254 13249
rect 31196 13209 31208 13243
rect 31242 13240 31254 13243
rect 31938 13240 31944 13252
rect 31242 13212 31944 13240
rect 31242 13209 31254 13212
rect 31196 13203 31254 13209
rect 31938 13200 31944 13212
rect 31996 13200 32002 13252
rect 33036 13243 33094 13249
rect 33036 13209 33048 13243
rect 33082 13240 33094 13243
rect 33778 13240 33784 13252
rect 33082 13212 33784 13240
rect 33082 13209 33094 13212
rect 33036 13203 33094 13209
rect 33778 13200 33784 13212
rect 33836 13200 33842 13252
rect 34992 13240 35020 13339
rect 37550 13336 37556 13348
rect 37608 13336 37614 13388
rect 51994 13376 52000 13388
rect 51955 13348 52000 13376
rect 51994 13336 52000 13348
rect 52052 13336 52058 13388
rect 35244 13311 35302 13317
rect 35244 13277 35256 13311
rect 35290 13308 35302 13311
rect 36354 13308 36360 13320
rect 35290 13280 36360 13308
rect 35290 13277 35302 13280
rect 35244 13271 35302 13277
rect 36354 13268 36360 13280
rect 36412 13268 36418 13320
rect 41417 13311 41475 13317
rect 41417 13277 41429 13311
rect 41463 13308 41475 13311
rect 42518 13308 42524 13320
rect 41463 13280 42524 13308
rect 41463 13277 41475 13280
rect 41417 13271 41475 13277
rect 42518 13268 42524 13280
rect 42576 13268 42582 13320
rect 45005 13311 45063 13317
rect 45005 13277 45017 13311
rect 45051 13308 45063 13311
rect 45554 13308 45560 13320
rect 45051 13280 45560 13308
rect 45051 13277 45063 13280
rect 45005 13271 45063 13277
rect 45554 13268 45560 13280
rect 45612 13268 45618 13320
rect 47946 13308 47952 13320
rect 47907 13280 47952 13308
rect 47946 13268 47952 13280
rect 48004 13268 48010 13320
rect 48216 13311 48274 13317
rect 48216 13277 48228 13311
rect 48262 13308 48274 13311
rect 49786 13308 49792 13320
rect 48262 13280 49792 13308
rect 48262 13277 48274 13280
rect 48216 13271 48274 13277
rect 49786 13268 49792 13280
rect 49844 13268 49850 13320
rect 50157 13311 50215 13317
rect 50157 13277 50169 13311
rect 50203 13277 50215 13311
rect 50157 13271 50215 13277
rect 50424 13311 50482 13317
rect 50424 13277 50436 13311
rect 50470 13308 50482 13311
rect 51166 13308 51172 13320
rect 50470 13280 51172 13308
rect 50470 13277 50482 13280
rect 50424 13271 50482 13277
rect 37550 13240 37556 13252
rect 34992 13212 37556 13240
rect 37550 13200 37556 13212
rect 37608 13200 37614 13252
rect 37820 13243 37878 13249
rect 37820 13209 37832 13243
rect 37866 13240 37878 13243
rect 38838 13240 38844 13252
rect 37866 13212 38844 13240
rect 37866 13209 37878 13212
rect 37820 13203 37878 13209
rect 38838 13200 38844 13212
rect 38896 13200 38902 13252
rect 41684 13243 41742 13249
rect 41684 13209 41696 13243
rect 41730 13240 41742 13243
rect 43898 13240 43904 13252
rect 41730 13212 43904 13240
rect 41730 13209 41742 13212
rect 41684 13203 41742 13209
rect 43898 13200 43904 13212
rect 43956 13200 43962 13252
rect 45272 13243 45330 13249
rect 45272 13209 45284 13243
rect 45318 13240 45330 13243
rect 45738 13240 45744 13252
rect 45318 13212 45744 13240
rect 45318 13209 45330 13212
rect 45272 13203 45330 13209
rect 45738 13200 45744 13212
rect 45796 13200 45802 13252
rect 50172 13240 50200 13271
rect 51166 13268 51172 13280
rect 51224 13268 51230 13320
rect 52264 13311 52322 13317
rect 52264 13277 52276 13311
rect 52310 13308 52322 13311
rect 53374 13308 53380 13320
rect 52310 13280 53380 13308
rect 52310 13277 52322 13280
rect 52264 13271 52322 13277
rect 53374 13268 53380 13280
rect 53432 13268 53438 13320
rect 56686 13308 56692 13320
rect 56647 13280 56692 13308
rect 56686 13268 56692 13280
rect 56744 13268 56750 13320
rect 50172 13212 51212 13240
rect 51184 13184 51212 13212
rect 3234 13172 3240 13184
rect 3195 13144 3240 13172
rect 3234 13132 3240 13144
rect 3292 13132 3298 13184
rect 6362 13172 6368 13184
rect 6323 13144 6368 13172
rect 6362 13132 6368 13144
rect 6420 13132 6426 13184
rect 10318 13172 10324 13184
rect 10279 13144 10324 13172
rect 10318 13132 10324 13144
rect 10376 13132 10382 13184
rect 16666 13132 16672 13184
rect 16724 13172 16730 13184
rect 16853 13175 16911 13181
rect 16853 13172 16865 13175
rect 16724 13144 16865 13172
rect 16724 13132 16730 13144
rect 16853 13141 16865 13144
rect 16899 13141 16911 13175
rect 22094 13172 22100 13184
rect 22055 13144 22100 13172
rect 16853 13135 16911 13141
rect 22094 13132 22100 13144
rect 22152 13132 22158 13184
rect 28534 13172 28540 13184
rect 28495 13144 28540 13172
rect 28534 13132 28540 13144
rect 28592 13132 28598 13184
rect 32309 13175 32367 13181
rect 32309 13141 32321 13175
rect 32355 13172 32367 13175
rect 32398 13172 32404 13184
rect 32355 13144 32404 13172
rect 32355 13141 32367 13144
rect 32309 13135 32367 13141
rect 32398 13132 32404 13144
rect 32456 13132 32462 13184
rect 34149 13175 34207 13181
rect 34149 13141 34161 13175
rect 34195 13172 34207 13175
rect 34238 13172 34244 13184
rect 34195 13144 34244 13172
rect 34195 13141 34207 13144
rect 34149 13135 34207 13141
rect 34238 13132 34244 13144
rect 34296 13132 34302 13184
rect 51166 13132 51172 13184
rect 51224 13132 51230 13184
rect 57238 13132 57244 13184
rect 57296 13172 57302 13184
rect 57977 13175 58035 13181
rect 57977 13172 57989 13175
rect 57296 13144 57989 13172
rect 57296 13132 57302 13144
rect 57977 13141 57989 13144
rect 58023 13141 58035 13175
rect 57977 13135 58035 13141
rect 1104 13082 59340 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 59340 13082
rect 1104 13008 59340 13030
rect 3513 12971 3571 12977
rect 3513 12937 3525 12971
rect 3559 12937 3571 12971
rect 7742 12968 7748 12980
rect 7703 12940 7748 12968
rect 3513 12931 3571 12937
rect 2400 12903 2458 12909
rect 2400 12869 2412 12903
rect 2446 12900 2458 12903
rect 3234 12900 3240 12912
rect 2446 12872 3240 12900
rect 2446 12869 2458 12872
rect 2400 12863 2458 12869
rect 3234 12860 3240 12872
rect 3292 12860 3298 12912
rect 3528 12900 3556 12931
rect 7742 12928 7748 12940
rect 7800 12928 7806 12980
rect 9766 12928 9772 12980
rect 9824 12928 9830 12980
rect 10962 12968 10968 12980
rect 10923 12940 10968 12968
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 14550 12928 14556 12980
rect 14608 12968 14614 12980
rect 15197 12971 15255 12977
rect 15197 12968 15209 12971
rect 14608 12940 15209 12968
rect 14608 12928 14614 12940
rect 15197 12937 15209 12940
rect 15243 12937 15255 12971
rect 21266 12968 21272 12980
rect 21227 12940 21272 12968
rect 15197 12931 15255 12937
rect 21266 12928 21272 12940
rect 21324 12928 21330 12980
rect 36078 12968 36084 12980
rect 36039 12940 36084 12968
rect 36078 12928 36084 12940
rect 36136 12928 36142 12980
rect 38838 12928 38844 12980
rect 38896 12968 38902 12980
rect 38933 12971 38991 12977
rect 38933 12968 38945 12971
rect 38896 12940 38945 12968
rect 38896 12928 38902 12940
rect 38933 12937 38945 12940
rect 38979 12937 38991 12971
rect 46750 12968 46756 12980
rect 46711 12940 46756 12968
rect 38933 12931 38991 12937
rect 46750 12928 46756 12940
rect 46808 12928 46814 12980
rect 51905 12971 51963 12977
rect 51905 12937 51917 12971
rect 51951 12937 51963 12971
rect 54846 12968 54852 12980
rect 54807 12940 54852 12968
rect 51905 12931 51963 12937
rect 4218 12903 4276 12909
rect 4218 12900 4230 12903
rect 3528 12872 4230 12900
rect 4218 12869 4230 12872
rect 4264 12869 4276 12903
rect 4218 12863 4276 12869
rect 1854 12792 1860 12844
rect 1912 12832 1918 12844
rect 2133 12835 2191 12841
rect 2133 12832 2145 12835
rect 1912 12804 2145 12832
rect 1912 12792 1918 12804
rect 2133 12801 2145 12804
rect 2179 12832 2191 12835
rect 6632 12835 6690 12841
rect 2179 12804 3924 12832
rect 2179 12801 2191 12804
rect 2133 12795 2191 12801
rect 3896 12776 3924 12804
rect 6632 12801 6644 12835
rect 6678 12832 6690 12835
rect 7742 12832 7748 12844
rect 6678 12804 7748 12832
rect 6678 12801 6690 12804
rect 6632 12795 6690 12801
rect 7742 12792 7748 12804
rect 7800 12792 7806 12844
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 9784 12832 9812 12928
rect 9852 12903 9910 12909
rect 9852 12869 9864 12903
rect 9898 12900 9910 12903
rect 10318 12900 10324 12912
rect 9898 12872 10324 12900
rect 9898 12869 9910 12872
rect 9852 12863 9910 12869
rect 10318 12860 10324 12872
rect 10376 12860 10382 12912
rect 14084 12903 14142 12909
rect 14084 12869 14096 12903
rect 14130 12900 14142 12903
rect 15470 12900 15476 12912
rect 14130 12872 15476 12900
rect 14130 12869 14142 12872
rect 14084 12863 14142 12869
rect 15470 12860 15476 12872
rect 15528 12860 15534 12912
rect 20156 12903 20214 12909
rect 20156 12869 20168 12903
rect 20202 12900 20214 12903
rect 22094 12900 22100 12912
rect 20202 12872 22100 12900
rect 20202 12869 20214 12872
rect 20156 12863 20214 12869
rect 22094 12860 22100 12872
rect 22152 12860 22158 12912
rect 24020 12903 24078 12909
rect 24020 12869 24032 12903
rect 24066 12900 24078 12903
rect 24486 12900 24492 12912
rect 24066 12872 24492 12900
rect 24066 12869 24078 12872
rect 24020 12863 24078 12869
rect 24486 12860 24492 12872
rect 24544 12860 24550 12912
rect 27516 12903 27574 12909
rect 27516 12869 27528 12903
rect 27562 12900 27574 12903
rect 28534 12900 28540 12912
rect 27562 12872 28540 12900
rect 27562 12869 27574 12872
rect 27516 12863 27574 12869
rect 28534 12860 28540 12872
rect 28592 12860 28598 12912
rect 32858 12900 32864 12912
rect 32140 12872 32864 12900
rect 32140 12844 32168 12872
rect 32858 12860 32864 12872
rect 32916 12860 32922 12912
rect 34698 12860 34704 12912
rect 34756 12900 34762 12912
rect 34946 12903 35004 12909
rect 34946 12900 34958 12903
rect 34756 12872 34958 12900
rect 34756 12860 34762 12872
rect 34946 12869 34958 12872
rect 34992 12869 35004 12903
rect 44910 12900 44916 12912
rect 44871 12872 44916 12900
rect 34946 12863 35004 12869
rect 44910 12860 44916 12872
rect 44968 12900 44974 12912
rect 48952 12903 49010 12909
rect 44968 12872 45416 12900
rect 44968 12860 44974 12872
rect 9631 12804 9812 12832
rect 16669 12835 16727 12841
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 16669 12801 16681 12835
rect 16715 12832 16727 12835
rect 16758 12832 16764 12844
rect 16715 12804 16764 12832
rect 16715 12801 16727 12804
rect 16669 12795 16727 12801
rect 16758 12792 16764 12804
rect 16816 12792 16822 12844
rect 16936 12835 16994 12841
rect 16936 12801 16948 12835
rect 16982 12832 16994 12835
rect 17954 12832 17960 12844
rect 16982 12804 17960 12832
rect 16982 12801 16994 12804
rect 16936 12795 16994 12801
rect 17954 12792 17960 12804
rect 18012 12792 18018 12844
rect 19889 12835 19947 12841
rect 19889 12801 19901 12835
rect 19935 12832 19947 12835
rect 20714 12832 20720 12844
rect 19935 12804 20720 12832
rect 19935 12801 19947 12804
rect 19889 12795 19947 12801
rect 20714 12792 20720 12804
rect 20772 12792 20778 12844
rect 23753 12835 23811 12841
rect 23753 12801 23765 12835
rect 23799 12832 23811 12835
rect 24394 12832 24400 12844
rect 23799 12804 24400 12832
rect 23799 12801 23811 12804
rect 23753 12795 23811 12801
rect 24394 12792 24400 12804
rect 24452 12792 24458 12844
rect 27249 12835 27307 12841
rect 27249 12801 27261 12835
rect 27295 12832 27307 12835
rect 27338 12832 27344 12844
rect 27295 12804 27344 12832
rect 27295 12801 27307 12804
rect 27249 12795 27307 12801
rect 27338 12792 27344 12804
rect 27396 12792 27402 12844
rect 28994 12792 29000 12844
rect 29052 12832 29058 12844
rect 29345 12835 29403 12841
rect 29345 12832 29357 12835
rect 29052 12804 29357 12832
rect 29052 12792 29058 12804
rect 29345 12801 29357 12804
rect 29391 12801 29403 12835
rect 32122 12832 32128 12844
rect 32035 12804 32128 12832
rect 29345 12795 29403 12801
rect 32122 12792 32128 12804
rect 32180 12792 32186 12844
rect 32392 12835 32450 12841
rect 32392 12801 32404 12835
rect 32438 12832 32450 12835
rect 33410 12832 33416 12844
rect 32438 12804 33416 12832
rect 32438 12801 32450 12804
rect 32392 12795 32450 12801
rect 33410 12792 33416 12804
rect 33468 12792 33474 12844
rect 34790 12832 34796 12844
rect 34716 12804 34796 12832
rect 3878 12724 3884 12776
rect 3936 12764 3942 12776
rect 3973 12767 4031 12773
rect 3973 12764 3985 12767
rect 3936 12736 3985 12764
rect 3936 12724 3942 12736
rect 3973 12733 3985 12736
rect 4019 12733 4031 12767
rect 3973 12727 4031 12733
rect 5626 12724 5632 12776
rect 5684 12764 5690 12776
rect 6270 12764 6276 12776
rect 5684 12736 6276 12764
rect 5684 12724 5690 12736
rect 6270 12724 6276 12736
rect 6328 12764 6334 12776
rect 6365 12767 6423 12773
rect 6365 12764 6377 12767
rect 6328 12736 6377 12764
rect 6328 12724 6334 12736
rect 6365 12733 6377 12736
rect 6411 12733 6423 12767
rect 13814 12764 13820 12776
rect 13775 12736 13820 12764
rect 6365 12727 6423 12733
rect 13814 12724 13820 12736
rect 13872 12724 13878 12776
rect 34716 12773 34744 12804
rect 34790 12792 34796 12804
rect 34848 12792 34854 12844
rect 37550 12832 37556 12844
rect 37511 12804 37556 12832
rect 37550 12792 37556 12804
rect 37608 12792 37614 12844
rect 37820 12835 37878 12841
rect 37820 12801 37832 12835
rect 37866 12832 37878 12835
rect 38930 12832 38936 12844
rect 37866 12804 38936 12832
rect 37866 12801 37878 12804
rect 37820 12795 37878 12801
rect 38930 12792 38936 12804
rect 38988 12792 38994 12844
rect 43162 12832 43168 12844
rect 43123 12804 43168 12832
rect 43162 12792 43168 12804
rect 43220 12792 43226 12844
rect 45388 12841 45416 12872
rect 48952 12869 48964 12903
rect 48998 12900 49010 12903
rect 51920 12900 51948 12931
rect 54846 12928 54852 12940
rect 54904 12928 54910 12980
rect 53742 12909 53748 12912
rect 53736 12900 53748 12909
rect 48998 12872 51948 12900
rect 53703 12872 53748 12900
rect 48998 12869 49010 12872
rect 48952 12863 49010 12869
rect 53736 12863 53748 12872
rect 53742 12860 53748 12863
rect 53800 12860 53806 12912
rect 45646 12841 45652 12844
rect 45373 12835 45431 12841
rect 45373 12801 45385 12835
rect 45419 12801 45431 12835
rect 45373 12795 45431 12801
rect 45640 12795 45652 12841
rect 45704 12832 45710 12844
rect 45704 12804 45740 12832
rect 45646 12792 45652 12795
rect 45704 12792 45710 12804
rect 48222 12792 48228 12844
rect 48280 12832 48286 12844
rect 48685 12835 48743 12841
rect 48685 12832 48697 12835
rect 48280 12804 48697 12832
rect 48280 12792 48286 12804
rect 48685 12801 48697 12804
rect 48731 12832 48743 12835
rect 48731 12804 50568 12832
rect 48731 12801 48743 12804
rect 48685 12795 48743 12801
rect 50540 12773 50568 12804
rect 50614 12792 50620 12844
rect 50672 12832 50678 12844
rect 50781 12835 50839 12841
rect 50781 12832 50793 12835
rect 50672 12804 50793 12832
rect 50672 12792 50678 12804
rect 50781 12801 50793 12804
rect 50827 12801 50839 12835
rect 50781 12795 50839 12801
rect 51994 12792 52000 12844
rect 52052 12832 52058 12844
rect 52362 12832 52368 12844
rect 52052 12804 52368 12832
rect 52052 12792 52058 12804
rect 52362 12792 52368 12804
rect 52420 12832 52426 12844
rect 53469 12835 53527 12841
rect 53469 12832 53481 12835
rect 52420 12804 53481 12832
rect 52420 12792 52426 12804
rect 53469 12801 53481 12804
rect 53515 12801 53527 12835
rect 53469 12795 53527 12801
rect 55490 12792 55496 12844
rect 55548 12832 55554 12844
rect 56209 12835 56267 12841
rect 56209 12832 56221 12835
rect 55548 12804 56221 12832
rect 55548 12792 55554 12804
rect 56209 12801 56221 12804
rect 56255 12801 56267 12835
rect 56209 12795 56267 12801
rect 29089 12767 29147 12773
rect 29089 12733 29101 12767
rect 29135 12733 29147 12767
rect 29089 12727 29147 12733
rect 34701 12767 34759 12773
rect 34701 12733 34713 12767
rect 34747 12733 34759 12767
rect 34701 12727 34759 12733
rect 50525 12767 50583 12773
rect 50525 12733 50537 12767
rect 50571 12733 50583 12767
rect 50525 12727 50583 12733
rect 5350 12628 5356 12640
rect 5311 12600 5356 12628
rect 5350 12588 5356 12600
rect 5408 12588 5414 12640
rect 18049 12631 18107 12637
rect 18049 12597 18061 12631
rect 18095 12628 18107 12631
rect 18138 12628 18144 12640
rect 18095 12600 18144 12628
rect 18095 12597 18107 12600
rect 18049 12591 18107 12597
rect 18138 12588 18144 12600
rect 18196 12588 18202 12640
rect 25130 12628 25136 12640
rect 25091 12600 25136 12628
rect 25130 12588 25136 12600
rect 25188 12588 25194 12640
rect 28626 12628 28632 12640
rect 28587 12600 28632 12628
rect 28626 12588 28632 12600
rect 28684 12588 28690 12640
rect 29104 12628 29132 12727
rect 29270 12628 29276 12640
rect 29104 12600 29276 12628
rect 29270 12588 29276 12600
rect 29328 12588 29334 12640
rect 29362 12588 29368 12640
rect 29420 12628 29426 12640
rect 30469 12631 30527 12637
rect 30469 12628 30481 12631
rect 29420 12600 30481 12628
rect 29420 12588 29426 12600
rect 30469 12597 30481 12600
rect 30515 12597 30527 12631
rect 33502 12628 33508 12640
rect 33463 12600 33508 12628
rect 30469 12591 30527 12597
rect 33502 12588 33508 12600
rect 33560 12588 33566 12640
rect 50062 12628 50068 12640
rect 50023 12600 50068 12628
rect 50062 12588 50068 12600
rect 50120 12588 50126 12640
rect 50540 12628 50568 12727
rect 55398 12724 55404 12776
rect 55456 12764 55462 12776
rect 55950 12764 55956 12776
rect 55456 12736 55956 12764
rect 55456 12724 55462 12736
rect 55950 12724 55956 12736
rect 56008 12724 56014 12776
rect 51166 12628 51172 12640
rect 50540 12600 51172 12628
rect 51166 12588 51172 12600
rect 51224 12588 51230 12640
rect 56594 12588 56600 12640
rect 56652 12628 56658 12640
rect 57333 12631 57391 12637
rect 57333 12628 57345 12631
rect 56652 12600 57345 12628
rect 56652 12588 56658 12600
rect 57333 12597 57345 12600
rect 57379 12597 57391 12631
rect 57333 12591 57391 12597
rect 1104 12538 59340 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 59340 12538
rect 1104 12464 59340 12486
rect 9766 12424 9772 12436
rect 9416 12396 9772 12424
rect 5626 12288 5632 12300
rect 5587 12260 5632 12288
rect 5626 12248 5632 12260
rect 5684 12248 5690 12300
rect 9416 12297 9444 12396
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 11146 12384 11152 12436
rect 11204 12424 11210 12436
rect 15286 12424 15292 12436
rect 11204 12396 15292 12424
rect 11204 12384 11210 12396
rect 15286 12384 15292 12396
rect 15344 12384 15350 12436
rect 15378 12384 15384 12436
rect 15436 12424 15442 12436
rect 15473 12427 15531 12433
rect 15473 12424 15485 12427
rect 15436 12396 15485 12424
rect 15436 12384 15442 12396
rect 15473 12393 15485 12396
rect 15519 12393 15531 12427
rect 22278 12424 22284 12436
rect 22239 12396 22284 12424
rect 15473 12387 15531 12393
rect 22278 12384 22284 12396
rect 22336 12384 22342 12436
rect 28813 12427 28871 12433
rect 28813 12393 28825 12427
rect 28859 12424 28871 12427
rect 28994 12424 29000 12436
rect 28859 12396 29000 12424
rect 28859 12393 28871 12396
rect 28813 12387 28871 12393
rect 28994 12384 29000 12396
rect 29052 12384 29058 12436
rect 38930 12424 38936 12436
rect 38891 12396 38936 12424
rect 38930 12384 38936 12396
rect 38988 12384 38994 12436
rect 39850 12384 39856 12436
rect 39908 12424 39914 12436
rect 41690 12424 41696 12436
rect 39908 12396 41696 12424
rect 39908 12384 39914 12396
rect 41690 12384 41696 12396
rect 41748 12424 41754 12436
rect 43162 12424 43168 12436
rect 41748 12396 43168 12424
rect 41748 12384 41754 12396
rect 43162 12384 43168 12396
rect 43220 12384 43226 12436
rect 43898 12424 43904 12436
rect 43859 12396 43904 12424
rect 43898 12384 43904 12396
rect 43956 12384 43962 12436
rect 9401 12291 9459 12297
rect 9401 12257 9413 12291
rect 9447 12257 9459 12291
rect 9401 12251 9459 12257
rect 24118 12248 24124 12300
rect 24176 12288 24182 12300
rect 24394 12288 24400 12300
rect 24176 12260 24400 12288
rect 24176 12248 24182 12260
rect 24394 12248 24400 12260
rect 24452 12248 24458 12300
rect 37550 12288 37556 12300
rect 37511 12260 37556 12288
rect 37550 12248 37556 12260
rect 37608 12248 37614 12300
rect 45554 12248 45560 12300
rect 45612 12288 45618 12300
rect 45830 12288 45836 12300
rect 45612 12260 45836 12288
rect 45612 12248 45618 12260
rect 45830 12248 45836 12260
rect 45888 12288 45894 12300
rect 46385 12291 46443 12297
rect 46385 12288 46397 12291
rect 45888 12260 46397 12288
rect 45888 12248 45894 12260
rect 46385 12257 46397 12260
rect 46431 12257 46443 12291
rect 48222 12288 48228 12300
rect 48183 12260 48228 12288
rect 46385 12251 46443 12257
rect 48222 12248 48228 12260
rect 48280 12248 48286 12300
rect 52362 12248 52368 12300
rect 52420 12288 52426 12300
rect 53009 12291 53067 12297
rect 53009 12288 53021 12291
rect 52420 12260 53021 12288
rect 52420 12248 52426 12260
rect 53009 12257 53021 12260
rect 53055 12257 53067 12291
rect 53009 12251 53067 12257
rect 56870 12248 56876 12300
rect 56928 12288 56934 12300
rect 57238 12288 57244 12300
rect 56928 12260 57244 12288
rect 56928 12248 56934 12260
rect 57238 12248 57244 12260
rect 57296 12248 57302 12300
rect 3789 12223 3847 12229
rect 3789 12189 3801 12223
rect 3835 12220 3847 12223
rect 3878 12220 3884 12232
rect 3835 12192 3884 12220
rect 3835 12189 3847 12192
rect 3789 12183 3847 12189
rect 3878 12180 3884 12192
rect 3936 12220 3942 12232
rect 5534 12220 5540 12232
rect 3936 12192 5540 12220
rect 3936 12180 3942 12192
rect 5534 12180 5540 12192
rect 5592 12220 5598 12232
rect 9674 12229 9680 12232
rect 9668 12220 9680 12229
rect 5592 12192 6132 12220
rect 9635 12192 9680 12220
rect 5592 12180 5598 12192
rect 6104 12164 6132 12192
rect 9668 12183 9680 12192
rect 9674 12180 9680 12183
rect 9732 12180 9738 12232
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13872 12192 14105 12220
rect 13872 12180 13878 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 4056 12155 4114 12161
rect 4056 12121 4068 12155
rect 4102 12152 4114 12155
rect 4246 12152 4252 12164
rect 4102 12124 4252 12152
rect 4102 12121 4114 12124
rect 4056 12115 4114 12121
rect 4246 12112 4252 12124
rect 4304 12112 4310 12164
rect 5874 12155 5932 12161
rect 5874 12152 5886 12155
rect 5184 12124 5886 12152
rect 5184 12093 5212 12124
rect 5874 12121 5886 12124
rect 5920 12121 5932 12155
rect 5874 12115 5932 12121
rect 6086 12112 6092 12164
rect 6144 12112 6150 12164
rect 14108 12152 14136 12183
rect 14182 12180 14188 12232
rect 14240 12220 14246 12232
rect 14349 12223 14407 12229
rect 14349 12220 14361 12223
rect 14240 12192 14361 12220
rect 14240 12180 14246 12192
rect 14349 12189 14361 12192
rect 14395 12189 14407 12223
rect 14349 12183 14407 12189
rect 15933 12223 15991 12229
rect 15933 12189 15945 12223
rect 15979 12220 15991 12223
rect 16666 12220 16672 12232
rect 15979 12192 16672 12220
rect 15979 12189 15991 12192
rect 15933 12183 15991 12189
rect 15948 12152 15976 12183
rect 16666 12180 16672 12192
rect 16724 12180 16730 12232
rect 20901 12223 20959 12229
rect 20901 12189 20913 12223
rect 20947 12220 20959 12223
rect 24136 12220 24164 12248
rect 20947 12192 24164 12220
rect 24664 12223 24722 12229
rect 20947 12189 20959 12192
rect 20901 12183 20959 12189
rect 24664 12189 24676 12223
rect 24710 12220 24722 12223
rect 25130 12220 25136 12232
rect 24710 12192 25136 12220
rect 24710 12189 24722 12192
rect 24664 12183 24722 12189
rect 25130 12180 25136 12192
rect 25188 12180 25194 12232
rect 27430 12220 27436 12232
rect 27391 12192 27436 12220
rect 27430 12180 27436 12192
rect 27488 12180 27494 12232
rect 27700 12223 27758 12229
rect 27700 12189 27712 12223
rect 27746 12220 27758 12223
rect 28626 12220 28632 12232
rect 27746 12192 28632 12220
rect 27746 12189 27758 12192
rect 27700 12183 27758 12189
rect 28626 12180 28632 12192
rect 28684 12180 28690 12232
rect 29270 12180 29276 12232
rect 29328 12220 29334 12232
rect 29549 12223 29607 12229
rect 29549 12220 29561 12223
rect 29328 12192 29561 12220
rect 29328 12180 29334 12192
rect 29549 12189 29561 12192
rect 29595 12189 29607 12223
rect 29549 12183 29607 12189
rect 29816 12223 29874 12229
rect 29816 12189 29828 12223
rect 29862 12220 29874 12223
rect 30190 12220 30196 12232
rect 29862 12192 30196 12220
rect 29862 12189 29874 12192
rect 29816 12183 29874 12189
rect 14108 12124 15976 12152
rect 16200 12155 16258 12161
rect 16200 12121 16212 12155
rect 16246 12152 16258 12155
rect 17218 12152 17224 12164
rect 16246 12124 17224 12152
rect 16246 12121 16258 12124
rect 16200 12115 16258 12121
rect 17218 12112 17224 12124
rect 17276 12112 17282 12164
rect 21168 12155 21226 12161
rect 21168 12121 21180 12155
rect 21214 12152 21226 12155
rect 23474 12152 23480 12164
rect 21214 12124 23480 12152
rect 21214 12121 21226 12124
rect 21168 12115 21226 12121
rect 23474 12112 23480 12124
rect 23532 12112 23538 12164
rect 29564 12152 29592 12183
rect 30190 12180 30196 12192
rect 30248 12180 30254 12232
rect 31389 12223 31447 12229
rect 31389 12220 31401 12223
rect 30300 12192 31401 12220
rect 30300 12152 30328 12192
rect 31389 12189 31401 12192
rect 31435 12220 31447 12223
rect 32122 12220 32128 12232
rect 31435 12192 32128 12220
rect 31435 12189 31447 12192
rect 31389 12183 31447 12189
rect 32122 12180 32128 12192
rect 32180 12180 32186 12232
rect 34701 12223 34759 12229
rect 34701 12189 34713 12223
rect 34747 12220 34759 12223
rect 34790 12220 34796 12232
rect 34747 12192 34796 12220
rect 34747 12189 34759 12192
rect 34701 12183 34759 12189
rect 34790 12180 34796 12192
rect 34848 12180 34854 12232
rect 40494 12180 40500 12232
rect 40552 12220 40558 12232
rect 40681 12223 40739 12229
rect 40681 12220 40693 12223
rect 40552 12192 40693 12220
rect 40552 12180 40558 12192
rect 40681 12189 40693 12192
rect 40727 12220 40739 12223
rect 42518 12220 42524 12232
rect 40727 12192 42524 12220
rect 40727 12189 40739 12192
rect 40681 12183 40739 12189
rect 42518 12180 42524 12192
rect 42576 12180 42582 12232
rect 51166 12220 51172 12232
rect 51079 12192 51172 12220
rect 51166 12180 51172 12192
rect 51224 12220 51230 12232
rect 52380 12220 52408 12248
rect 51224 12192 52408 12220
rect 53276 12223 53334 12229
rect 51224 12180 51230 12192
rect 53276 12189 53288 12223
rect 53322 12220 53334 12223
rect 53650 12220 53656 12232
rect 53322 12192 53656 12220
rect 53322 12189 53334 12192
rect 53276 12183 53334 12189
rect 53650 12180 53656 12192
rect 53708 12180 53714 12232
rect 55398 12220 55404 12232
rect 55359 12192 55404 12220
rect 55398 12180 55404 12192
rect 55456 12180 55462 12232
rect 55668 12223 55726 12229
rect 55668 12189 55680 12223
rect 55714 12220 55726 12223
rect 56594 12220 56600 12232
rect 55714 12192 56600 12220
rect 55714 12189 55726 12192
rect 55668 12183 55726 12189
rect 56594 12180 56600 12192
rect 56652 12180 56658 12232
rect 57514 12229 57520 12232
rect 57508 12183 57520 12229
rect 57572 12220 57578 12232
rect 57572 12192 57608 12220
rect 57514 12180 57520 12183
rect 57572 12180 57578 12192
rect 29564 12124 30328 12152
rect 31110 12112 31116 12164
rect 31168 12152 31174 12164
rect 31634 12155 31692 12161
rect 31634 12152 31646 12155
rect 31168 12124 31646 12152
rect 31168 12112 31174 12124
rect 31634 12121 31646 12124
rect 31680 12121 31692 12155
rect 31634 12115 31692 12121
rect 34968 12155 35026 12161
rect 34968 12121 34980 12155
rect 35014 12152 35026 12155
rect 35986 12152 35992 12164
rect 35014 12124 35992 12152
rect 35014 12121 35026 12124
rect 34968 12115 35026 12121
rect 35986 12112 35992 12124
rect 36044 12112 36050 12164
rect 37820 12155 37878 12161
rect 37820 12121 37832 12155
rect 37866 12152 37878 12155
rect 38838 12152 38844 12164
rect 37866 12124 38844 12152
rect 37866 12121 37878 12124
rect 37820 12115 37878 12121
rect 38838 12112 38844 12124
rect 38896 12112 38902 12164
rect 40948 12155 41006 12161
rect 40948 12121 40960 12155
rect 40994 12152 41006 12155
rect 41874 12152 41880 12164
rect 40994 12124 41880 12152
rect 40994 12121 41006 12124
rect 40948 12115 41006 12121
rect 41874 12112 41880 12124
rect 41932 12112 41938 12164
rect 42766 12155 42824 12161
rect 42766 12152 42778 12155
rect 42076 12124 42778 12152
rect 5169 12087 5227 12093
rect 5169 12053 5181 12087
rect 5215 12053 5227 12087
rect 7006 12084 7012 12096
rect 6967 12056 7012 12084
rect 5169 12047 5227 12053
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 10778 12084 10784 12096
rect 10739 12056 10784 12084
rect 10778 12044 10784 12056
rect 10836 12044 10842 12096
rect 17310 12084 17316 12096
rect 17271 12056 17316 12084
rect 17310 12044 17316 12056
rect 17368 12044 17374 12096
rect 25774 12084 25780 12096
rect 25735 12056 25780 12084
rect 25774 12044 25780 12056
rect 25832 12044 25838 12096
rect 30926 12084 30932 12096
rect 30887 12056 30932 12084
rect 30926 12044 30932 12056
rect 30984 12044 30990 12096
rect 31202 12044 31208 12096
rect 31260 12084 31266 12096
rect 32769 12087 32827 12093
rect 32769 12084 32781 12087
rect 31260 12056 32781 12084
rect 31260 12044 31266 12056
rect 32769 12053 32781 12056
rect 32815 12053 32827 12087
rect 36078 12084 36084 12096
rect 36039 12056 36084 12084
rect 32769 12047 32827 12053
rect 36078 12044 36084 12056
rect 36136 12044 36142 12096
rect 42076 12093 42104 12124
rect 42766 12121 42778 12124
rect 42812 12121 42824 12155
rect 42766 12115 42824 12121
rect 46652 12155 46710 12161
rect 46652 12121 46664 12155
rect 46698 12152 46710 12155
rect 48492 12155 48550 12161
rect 46698 12124 48176 12152
rect 46698 12121 46710 12124
rect 46652 12115 46710 12121
rect 42061 12087 42119 12093
rect 42061 12053 42073 12087
rect 42107 12053 42119 12087
rect 47762 12084 47768 12096
rect 47723 12056 47768 12084
rect 42061 12047 42119 12053
rect 47762 12044 47768 12056
rect 47820 12044 47826 12096
rect 48148 12084 48176 12124
rect 48492 12121 48504 12155
rect 48538 12152 48550 12155
rect 50154 12152 50160 12164
rect 48538 12124 50160 12152
rect 48538 12121 48550 12124
rect 48492 12115 48550 12121
rect 50154 12112 50160 12124
rect 50212 12112 50218 12164
rect 51436 12155 51494 12161
rect 51436 12121 51448 12155
rect 51482 12152 51494 12155
rect 52914 12152 52920 12164
rect 51482 12124 52920 12152
rect 51482 12121 51494 12124
rect 51436 12115 51494 12121
rect 52914 12112 52920 12124
rect 52972 12112 52978 12164
rect 49605 12087 49663 12093
rect 49605 12084 49617 12087
rect 48148 12056 49617 12084
rect 49605 12053 49617 12056
rect 49651 12053 49663 12087
rect 49605 12047 49663 12053
rect 52549 12087 52607 12093
rect 52549 12053 52561 12087
rect 52595 12084 52607 12087
rect 53650 12084 53656 12096
rect 52595 12056 53656 12084
rect 52595 12053 52607 12056
rect 52549 12047 52607 12053
rect 53650 12044 53656 12056
rect 53708 12044 53714 12096
rect 54386 12084 54392 12096
rect 54347 12056 54392 12084
rect 54386 12044 54392 12056
rect 54444 12044 54450 12096
rect 56778 12084 56784 12096
rect 56739 12056 56784 12084
rect 56778 12044 56784 12056
rect 56836 12044 56842 12096
rect 58434 12044 58440 12096
rect 58492 12084 58498 12096
rect 58621 12087 58679 12093
rect 58621 12084 58633 12087
rect 58492 12056 58633 12084
rect 58492 12044 58498 12056
rect 58621 12053 58633 12056
rect 58667 12053 58679 12087
rect 58621 12047 58679 12053
rect 1104 11994 59340 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 59340 11994
rect 1104 11920 59340 11942
rect 4246 11880 4252 11892
rect 4207 11852 4252 11880
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 7742 11880 7748 11892
rect 7703 11852 7748 11880
rect 7742 11840 7748 11852
rect 7800 11840 7806 11892
rect 9766 11880 9772 11892
rect 9600 11852 9772 11880
rect 3136 11815 3194 11821
rect 3136 11781 3148 11815
rect 3182 11812 3194 11815
rect 5350 11812 5356 11824
rect 3182 11784 5356 11812
rect 3182 11781 3194 11784
rect 3136 11775 3194 11781
rect 5350 11772 5356 11784
rect 5408 11772 5414 11824
rect 6362 11772 6368 11824
rect 6420 11812 6426 11824
rect 6610 11815 6668 11821
rect 6610 11812 6622 11815
rect 6420 11784 6622 11812
rect 6420 11772 6426 11784
rect 6610 11781 6622 11784
rect 6656 11781 6668 11815
rect 6610 11775 6668 11781
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11744 2927 11747
rect 3878 11744 3884 11756
rect 2915 11716 3884 11744
rect 2915 11713 2927 11716
rect 2869 11707 2927 11713
rect 3878 11704 3884 11716
rect 3936 11704 3942 11756
rect 9401 11747 9459 11753
rect 9401 11713 9413 11747
rect 9447 11744 9459 11747
rect 9600 11744 9628 11852
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 13541 11883 13599 11889
rect 13541 11849 13553 11883
rect 13587 11849 13599 11883
rect 13541 11843 13599 11849
rect 9668 11815 9726 11821
rect 9668 11781 9680 11815
rect 9714 11812 9726 11815
rect 10778 11812 10784 11824
rect 9714 11784 10784 11812
rect 9714 11781 9726 11784
rect 9668 11775 9726 11781
rect 10778 11772 10784 11784
rect 10836 11772 10842 11824
rect 13556 11812 13584 11843
rect 22370 11840 22376 11892
rect 22428 11880 22434 11892
rect 23201 11883 23259 11889
rect 23201 11880 23213 11883
rect 22428 11852 23213 11880
rect 22428 11840 22434 11852
rect 23201 11849 23213 11852
rect 23247 11849 23259 11883
rect 23201 11843 23259 11849
rect 29086 11840 29092 11892
rect 29144 11880 29150 11892
rect 29273 11883 29331 11889
rect 29273 11880 29285 11883
rect 29144 11852 29285 11880
rect 29144 11840 29150 11852
rect 29273 11849 29285 11852
rect 29319 11849 29331 11883
rect 31110 11880 31116 11892
rect 31071 11852 31116 11880
rect 29273 11843 29331 11849
rect 31110 11840 31116 11852
rect 31168 11840 31174 11892
rect 33410 11840 33416 11892
rect 33468 11880 33474 11892
rect 33505 11883 33563 11889
rect 33505 11880 33517 11883
rect 33468 11852 33517 11880
rect 33468 11840 33474 11852
rect 33505 11849 33517 11852
rect 33551 11849 33563 11883
rect 38838 11880 38844 11892
rect 38799 11852 38844 11880
rect 33505 11843 33563 11849
rect 38838 11840 38844 11852
rect 38896 11840 38902 11892
rect 41874 11880 41880 11892
rect 41835 11852 41880 11880
rect 41874 11840 41880 11852
rect 41932 11840 41938 11892
rect 43809 11883 43867 11889
rect 43809 11849 43821 11883
rect 43855 11880 43867 11883
rect 45462 11880 45468 11892
rect 43855 11852 45468 11880
rect 43855 11849 43867 11852
rect 43809 11843 43867 11849
rect 45462 11840 45468 11852
rect 45520 11840 45526 11892
rect 45649 11883 45707 11889
rect 45649 11849 45661 11883
rect 45695 11880 45707 11883
rect 45738 11880 45744 11892
rect 45695 11852 45744 11880
rect 45695 11849 45707 11852
rect 45649 11843 45707 11849
rect 45738 11840 45744 11852
rect 45796 11840 45802 11892
rect 50154 11840 50160 11892
rect 50212 11880 50218 11892
rect 50341 11883 50399 11889
rect 50341 11880 50353 11883
rect 50212 11852 50353 11880
rect 50212 11840 50218 11852
rect 50341 11849 50353 11852
rect 50387 11849 50399 11883
rect 50341 11843 50399 11849
rect 55493 11883 55551 11889
rect 55493 11849 55505 11883
rect 55539 11880 55551 11883
rect 55582 11880 55588 11892
rect 55539 11852 55588 11880
rect 55539 11849 55551 11852
rect 55493 11843 55551 11849
rect 55582 11840 55588 11852
rect 55640 11840 55646 11892
rect 14246 11815 14304 11821
rect 14246 11812 14258 11815
rect 13556 11784 14258 11812
rect 14246 11781 14258 11784
rect 14292 11781 14304 11815
rect 14246 11775 14304 11781
rect 16936 11815 16994 11821
rect 16936 11781 16948 11815
rect 16982 11812 16994 11815
rect 17310 11812 17316 11824
rect 16982 11784 17316 11812
rect 16982 11781 16994 11784
rect 16936 11775 16994 11781
rect 17310 11772 17316 11784
rect 17368 11772 17374 11824
rect 22088 11815 22146 11821
rect 19904 11784 21864 11812
rect 9447 11716 9628 11744
rect 12428 11747 12486 11753
rect 9447 11713 9459 11716
rect 9401 11707 9459 11713
rect 12428 11713 12440 11747
rect 12474 11744 12486 11747
rect 15470 11744 15476 11756
rect 12474 11716 15476 11744
rect 12474 11713 12486 11716
rect 12428 11707 12486 11713
rect 15470 11704 15476 11716
rect 15528 11704 15534 11756
rect 19904 11688 19932 11784
rect 20156 11747 20214 11753
rect 20156 11713 20168 11747
rect 20202 11744 20214 11747
rect 21266 11744 21272 11756
rect 20202 11716 21272 11744
rect 20202 11713 20214 11716
rect 20156 11707 20214 11713
rect 21266 11704 21272 11716
rect 21324 11704 21330 11756
rect 21836 11753 21864 11784
rect 22088 11781 22100 11815
rect 22134 11812 22146 11815
rect 22186 11812 22192 11824
rect 22134 11784 22192 11812
rect 22134 11781 22146 11784
rect 22088 11775 22146 11781
rect 22186 11772 22192 11784
rect 22244 11772 22250 11824
rect 24388 11815 24446 11821
rect 24388 11781 24400 11815
rect 24434 11812 24446 11815
rect 25774 11812 25780 11824
rect 24434 11784 25780 11812
rect 24434 11781 24446 11784
rect 24388 11775 24446 11781
rect 25774 11772 25780 11784
rect 25832 11772 25838 11824
rect 28160 11815 28218 11821
rect 28160 11781 28172 11815
rect 28206 11812 28218 11815
rect 29362 11812 29368 11824
rect 28206 11784 29368 11812
rect 28206 11781 28218 11784
rect 28160 11775 28218 11781
rect 29362 11772 29368 11784
rect 29420 11772 29426 11824
rect 30000 11815 30058 11821
rect 30000 11781 30012 11815
rect 30046 11812 30058 11815
rect 30926 11812 30932 11824
rect 30046 11784 30932 11812
rect 30046 11781 30058 11784
rect 30000 11775 30058 11781
rect 30926 11772 30932 11784
rect 30984 11772 30990 11824
rect 42696 11815 42754 11821
rect 42696 11781 42708 11815
rect 42742 11812 42754 11815
rect 44266 11812 44272 11824
rect 42742 11784 44272 11812
rect 42742 11781 42754 11784
rect 42696 11775 42754 11781
rect 44266 11772 44272 11784
rect 44324 11772 44330 11824
rect 44542 11821 44548 11824
rect 44536 11812 44548 11821
rect 44503 11784 44548 11812
rect 44536 11775 44548 11784
rect 44542 11772 44548 11775
rect 44600 11772 44606 11824
rect 51166 11812 51172 11824
rect 50816 11784 51172 11812
rect 21821 11747 21879 11753
rect 21821 11713 21833 11747
rect 21867 11713 21879 11747
rect 24118 11744 24124 11756
rect 24079 11716 24124 11744
rect 21821 11707 21879 11713
rect 24118 11704 24124 11716
rect 24176 11704 24182 11756
rect 27430 11704 27436 11756
rect 27488 11744 27494 11756
rect 27893 11747 27951 11753
rect 27893 11744 27905 11747
rect 27488 11716 27905 11744
rect 27488 11704 27494 11716
rect 27893 11713 27905 11716
rect 27939 11744 27951 11747
rect 32122 11744 32128 11756
rect 27939 11716 29592 11744
rect 32083 11716 32128 11744
rect 27939 11713 27951 11716
rect 27893 11707 27951 11713
rect 29564 11688 29592 11716
rect 32122 11704 32128 11716
rect 32180 11704 32186 11756
rect 32398 11753 32404 11756
rect 32392 11744 32404 11753
rect 32359 11716 32404 11744
rect 32392 11707 32404 11716
rect 32398 11704 32404 11707
rect 32456 11704 32462 11756
rect 34238 11753 34244 11756
rect 34232 11744 34244 11753
rect 34199 11716 34244 11744
rect 34232 11707 34244 11716
rect 34238 11704 34244 11707
rect 34296 11704 34302 11756
rect 37461 11747 37519 11753
rect 37461 11713 37473 11747
rect 37507 11744 37519 11747
rect 37550 11744 37556 11756
rect 37507 11716 37556 11744
rect 37507 11713 37519 11716
rect 37461 11707 37519 11713
rect 37550 11704 37556 11716
rect 37608 11704 37614 11756
rect 37728 11747 37786 11753
rect 37728 11713 37740 11747
rect 37774 11744 37786 11747
rect 38746 11744 38752 11756
rect 37774 11716 38752 11744
rect 37774 11713 37786 11716
rect 37728 11707 37786 11713
rect 38746 11704 38752 11716
rect 38804 11704 38810 11756
rect 40494 11744 40500 11756
rect 40455 11716 40500 11744
rect 40494 11704 40500 11716
rect 40552 11704 40558 11756
rect 40764 11747 40822 11753
rect 40764 11713 40776 11747
rect 40810 11744 40822 11747
rect 41874 11744 41880 11756
rect 40810 11716 41880 11744
rect 40810 11713 40822 11716
rect 40764 11707 40822 11713
rect 41874 11704 41880 11716
rect 41932 11704 41938 11756
rect 42429 11747 42487 11753
rect 42429 11713 42441 11747
rect 42475 11744 42487 11747
rect 42518 11744 42524 11756
rect 42475 11716 42524 11744
rect 42475 11713 42487 11716
rect 42429 11707 42487 11713
rect 42518 11704 42524 11716
rect 42576 11744 42582 11756
rect 44910 11744 44916 11756
rect 42576 11716 44916 11744
rect 42576 11704 42582 11716
rect 6086 11636 6092 11688
rect 6144 11676 6150 11688
rect 6365 11679 6423 11685
rect 6365 11676 6377 11679
rect 6144 11648 6377 11676
rect 6144 11636 6150 11648
rect 6365 11645 6377 11648
rect 6411 11645 6423 11679
rect 12158 11676 12164 11688
rect 12119 11648 12164 11676
rect 6365 11639 6423 11645
rect 12158 11636 12164 11648
rect 12216 11636 12222 11688
rect 13998 11676 14004 11688
rect 13959 11648 14004 11676
rect 13998 11636 14004 11648
rect 14056 11636 14062 11688
rect 16666 11676 16672 11688
rect 16627 11648 16672 11676
rect 16666 11636 16672 11648
rect 16724 11636 16730 11688
rect 19886 11676 19892 11688
rect 19847 11648 19892 11676
rect 19886 11636 19892 11648
rect 19944 11636 19950 11688
rect 29546 11636 29552 11688
rect 29604 11676 29610 11688
rect 29733 11679 29791 11685
rect 29733 11676 29745 11679
rect 29604 11648 29745 11676
rect 29604 11636 29610 11648
rect 29733 11645 29745 11648
rect 29779 11645 29791 11679
rect 33962 11676 33968 11688
rect 33923 11648 33968 11676
rect 29733 11639 29791 11645
rect 33962 11636 33968 11648
rect 34020 11636 34026 11688
rect 44284 11685 44312 11716
rect 44910 11704 44916 11716
rect 44968 11704 44974 11756
rect 49228 11747 49286 11753
rect 49228 11713 49240 11747
rect 49274 11744 49286 11747
rect 49602 11744 49608 11756
rect 49274 11716 49608 11744
rect 49274 11713 49286 11716
rect 49228 11707 49286 11713
rect 49602 11704 49608 11716
rect 49660 11704 49666 11756
rect 50816 11753 50844 11784
rect 51166 11772 51172 11784
rect 51224 11772 51230 11824
rect 54380 11815 54438 11821
rect 54380 11781 54392 11815
rect 54426 11812 54438 11815
rect 56778 11812 56784 11824
rect 54426 11784 56784 11812
rect 54426 11781 54438 11784
rect 54380 11775 54438 11781
rect 56778 11772 56784 11784
rect 56836 11772 56842 11824
rect 58434 11812 58440 11824
rect 58395 11784 58440 11812
rect 58434 11772 58440 11784
rect 58492 11772 58498 11824
rect 50801 11747 50859 11753
rect 50801 11713 50813 11747
rect 50847 11713 50859 11747
rect 50801 11707 50859 11713
rect 51068 11747 51126 11753
rect 51068 11713 51080 11747
rect 51114 11744 51126 11747
rect 52086 11744 52092 11756
rect 51114 11716 52092 11744
rect 51114 11713 51126 11716
rect 51068 11707 51126 11713
rect 52086 11704 52092 11716
rect 52144 11704 52150 11756
rect 55398 11744 55404 11756
rect 54128 11716 55404 11744
rect 44269 11679 44327 11685
rect 44269 11645 44281 11679
rect 44315 11645 44327 11679
rect 44269 11639 44327 11645
rect 48590 11636 48596 11688
rect 48648 11676 48654 11688
rect 48961 11679 49019 11685
rect 48961 11676 48973 11679
rect 48648 11648 48973 11676
rect 48648 11636 48654 11648
rect 48961 11645 48973 11648
rect 49007 11645 49019 11679
rect 48961 11639 49019 11645
rect 53282 11636 53288 11688
rect 53340 11676 53346 11688
rect 54128 11685 54156 11716
rect 55398 11704 55404 11716
rect 55456 11744 55462 11756
rect 55953 11747 56011 11753
rect 55953 11744 55965 11747
rect 55456 11716 55965 11744
rect 55456 11704 55462 11716
rect 55953 11713 55965 11716
rect 55999 11713 56011 11747
rect 55953 11707 56011 11713
rect 56220 11747 56278 11753
rect 56220 11713 56232 11747
rect 56266 11744 56278 11747
rect 57238 11744 57244 11756
rect 56266 11716 57244 11744
rect 56266 11713 56278 11716
rect 56220 11707 56278 11713
rect 57238 11704 57244 11716
rect 57296 11704 57302 11756
rect 58618 11744 58624 11756
rect 58579 11716 58624 11744
rect 58618 11704 58624 11716
rect 58676 11704 58682 11756
rect 54113 11679 54171 11685
rect 54113 11676 54125 11679
rect 53340 11648 54125 11676
rect 53340 11636 53346 11648
rect 54113 11645 54125 11648
rect 54159 11645 54171 11679
rect 54113 11639 54171 11645
rect 10778 11540 10784 11552
rect 10739 11512 10784 11540
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 15378 11540 15384 11552
rect 15339 11512 15384 11540
rect 15378 11500 15384 11512
rect 15436 11500 15442 11552
rect 18046 11540 18052 11552
rect 18007 11512 18052 11540
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 21269 11543 21327 11549
rect 21269 11509 21281 11543
rect 21315 11540 21327 11543
rect 22094 11540 22100 11552
rect 21315 11512 22100 11540
rect 21315 11509 21327 11512
rect 21269 11503 21327 11509
rect 22094 11500 22100 11512
rect 22152 11500 22158 11552
rect 25498 11540 25504 11552
rect 25459 11512 25504 11540
rect 25498 11500 25504 11512
rect 25556 11500 25562 11552
rect 35342 11540 35348 11552
rect 35303 11512 35348 11540
rect 35342 11500 35348 11512
rect 35400 11500 35406 11552
rect 40402 11500 40408 11552
rect 40460 11540 40466 11552
rect 48406 11540 48412 11552
rect 40460 11512 48412 11540
rect 40460 11500 40466 11512
rect 48406 11500 48412 11512
rect 48464 11500 48470 11552
rect 51166 11500 51172 11552
rect 51224 11540 51230 11552
rect 52181 11543 52239 11549
rect 52181 11540 52193 11543
rect 51224 11512 52193 11540
rect 51224 11500 51230 11512
rect 52181 11509 52193 11512
rect 52227 11509 52239 11543
rect 52181 11503 52239 11509
rect 55950 11500 55956 11552
rect 56008 11540 56014 11552
rect 57333 11543 57391 11549
rect 57333 11540 57345 11543
rect 56008 11512 57345 11540
rect 56008 11500 56014 11512
rect 57333 11509 57345 11512
rect 57379 11509 57391 11543
rect 57333 11503 57391 11509
rect 1104 11450 59340 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 59340 11450
rect 1104 11376 59340 11398
rect 5810 11336 5816 11348
rect 5771 11308 5816 11336
rect 5810 11296 5816 11308
rect 5868 11296 5874 11348
rect 11146 11296 11152 11348
rect 11204 11336 11210 11348
rect 11517 11339 11575 11345
rect 11517 11336 11529 11339
rect 11204 11308 11529 11336
rect 11204 11296 11210 11308
rect 11517 11305 11529 11308
rect 11563 11305 11575 11339
rect 12158 11336 12164 11348
rect 12071 11308 12164 11336
rect 11517 11299 11575 11305
rect 11532 11268 11560 11299
rect 12158 11296 12164 11308
rect 12216 11336 12222 11348
rect 13998 11336 14004 11348
rect 12216 11308 14004 11336
rect 12216 11296 12222 11308
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 15470 11336 15476 11348
rect 15431 11308 15476 11336
rect 15470 11296 15476 11308
rect 15528 11296 15534 11348
rect 16666 11336 16672 11348
rect 15948 11308 16672 11336
rect 12066 11268 12072 11280
rect 11532 11240 12072 11268
rect 12066 11228 12072 11240
rect 12124 11228 12130 11280
rect 10962 11160 10968 11212
rect 11020 11200 11026 11212
rect 12176 11209 12204 11296
rect 13541 11271 13599 11277
rect 13541 11237 13553 11271
rect 13587 11268 13599 11271
rect 14090 11268 14096 11280
rect 13587 11240 14096 11268
rect 13587 11237 13599 11240
rect 13541 11231 13599 11237
rect 14090 11228 14096 11240
rect 14148 11228 14154 11280
rect 12161 11203 12219 11209
rect 12161 11200 12173 11203
rect 11020 11172 12173 11200
rect 11020 11160 11026 11172
rect 12161 11169 12173 11172
rect 12207 11169 12219 11203
rect 12161 11163 12219 11169
rect 13814 11160 13820 11212
rect 13872 11200 13878 11212
rect 15948 11209 15976 11308
rect 16666 11296 16672 11308
rect 16724 11296 16730 11348
rect 17218 11296 17224 11348
rect 17276 11336 17282 11348
rect 17313 11339 17371 11345
rect 17313 11336 17325 11339
rect 17276 11308 17325 11336
rect 17276 11296 17282 11308
rect 17313 11305 17325 11308
rect 17359 11305 17371 11339
rect 21266 11336 21272 11348
rect 21227 11308 21272 11336
rect 17313 11299 17371 11305
rect 21266 11296 21272 11308
rect 21324 11296 21330 11348
rect 23474 11336 23480 11348
rect 23435 11308 23480 11336
rect 23474 11296 23480 11308
rect 23532 11296 23538 11348
rect 31938 11336 31944 11348
rect 31899 11308 31944 11336
rect 31938 11296 31944 11308
rect 31996 11296 32002 11348
rect 33778 11336 33784 11348
rect 33739 11308 33784 11336
rect 33778 11296 33784 11308
rect 33836 11296 33842 11348
rect 35986 11296 35992 11348
rect 36044 11336 36050 11348
rect 36081 11339 36139 11345
rect 36081 11336 36093 11339
rect 36044 11308 36093 11336
rect 36044 11296 36050 11308
rect 36081 11305 36093 11308
rect 36127 11305 36139 11339
rect 38746 11336 38752 11348
rect 38707 11308 38752 11336
rect 36081 11299 36139 11305
rect 38746 11296 38752 11308
rect 38804 11296 38810 11348
rect 39850 11336 39856 11348
rect 39811 11308 39856 11336
rect 39850 11296 39856 11308
rect 39908 11296 39914 11348
rect 41874 11336 41880 11348
rect 41835 11308 41880 11336
rect 41874 11296 41880 11308
rect 41932 11296 41938 11348
rect 47946 11336 47952 11348
rect 46400 11308 47952 11336
rect 15933 11203 15991 11209
rect 13872 11172 14136 11200
rect 13872 11160 13878 11172
rect 4433 11135 4491 11141
rect 4433 11101 4445 11135
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 4700 11135 4758 11141
rect 4700 11101 4712 11135
rect 4746 11132 4758 11135
rect 7006 11132 7012 11144
rect 4746 11104 7012 11132
rect 4746 11101 4758 11104
rect 4700 11095 4758 11101
rect 4448 11064 4476 11095
rect 7006 11092 7012 11104
rect 7064 11092 7070 11144
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11101 9459 11135
rect 9401 11095 9459 11101
rect 9668 11135 9726 11141
rect 9668 11101 9680 11135
rect 9714 11132 9726 11135
rect 10778 11132 10784 11144
rect 9714 11104 10784 11132
rect 9714 11101 9726 11104
rect 9668 11095 9726 11101
rect 6086 11064 6092 11076
rect 4448 11036 6092 11064
rect 6086 11024 6092 11036
rect 6144 11024 6150 11076
rect 9416 11064 9444 11095
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 14108 11141 14136 11172
rect 15933 11169 15945 11203
rect 15979 11169 15991 11203
rect 40494 11200 40500 11212
rect 40455 11172 40500 11200
rect 15933 11163 15991 11169
rect 40494 11160 40500 11172
rect 40552 11160 40558 11212
rect 46400 11209 46428 11308
rect 47946 11296 47952 11308
rect 48004 11296 48010 11348
rect 49602 11336 49608 11348
rect 49563 11308 49608 11336
rect 49602 11296 49608 11308
rect 49660 11296 49666 11348
rect 52454 11296 52460 11348
rect 52512 11296 52518 11348
rect 52914 11336 52920 11348
rect 52875 11308 52920 11336
rect 52914 11296 52920 11308
rect 52972 11296 52978 11348
rect 52472 11268 52500 11296
rect 52472 11240 53420 11268
rect 53392 11209 53420 11240
rect 46385 11203 46443 11209
rect 46385 11169 46397 11203
rect 46431 11169 46443 11203
rect 46385 11163 46443 11169
rect 53377 11203 53435 11209
rect 53377 11169 53389 11203
rect 53423 11169 53435 11203
rect 56870 11200 56876 11212
rect 56831 11172 56876 11200
rect 53377 11163 53435 11169
rect 56870 11160 56876 11172
rect 56928 11160 56934 11212
rect 11701 11135 11759 11141
rect 11701 11101 11713 11135
rect 11747 11101 11759 11135
rect 14093 11135 14151 11141
rect 11701 11095 11759 11101
rect 12360 11104 14044 11132
rect 9858 11064 9864 11076
rect 9416 11036 9864 11064
rect 9858 11024 9864 11036
rect 9916 11064 9922 11076
rect 10962 11064 10968 11076
rect 9916 11036 10968 11064
rect 9916 11024 9922 11036
rect 10962 11024 10968 11036
rect 11020 11024 11026 11076
rect 11716 11064 11744 11095
rect 12360 11064 12388 11104
rect 11716 11036 12388 11064
rect 12428 11067 12486 11073
rect 12428 11033 12440 11067
rect 12474 11064 12486 11067
rect 13906 11064 13912 11076
rect 12474 11036 13912 11064
rect 12474 11033 12486 11036
rect 12428 11027 12486 11033
rect 13906 11024 13912 11036
rect 13964 11024 13970 11076
rect 14016 11064 14044 11104
rect 14093 11101 14105 11135
rect 14139 11101 14151 11135
rect 14093 11095 14151 11101
rect 14292 11104 15332 11132
rect 14292 11064 14320 11104
rect 14016 11036 14320 11064
rect 14360 11067 14418 11073
rect 14360 11033 14372 11067
rect 14406 11064 14418 11067
rect 15194 11064 15200 11076
rect 14406 11036 15200 11064
rect 14406 11033 14418 11036
rect 14360 11027 14418 11033
rect 15194 11024 15200 11036
rect 15252 11024 15258 11076
rect 15304 11064 15332 11104
rect 15378 11092 15384 11144
rect 15436 11132 15442 11144
rect 16189 11135 16247 11141
rect 16189 11132 16201 11135
rect 15436 11104 16201 11132
rect 15436 11092 15442 11104
rect 16189 11101 16201 11104
rect 16235 11101 16247 11135
rect 16189 11095 16247 11101
rect 19334 11092 19340 11144
rect 19392 11132 19398 11144
rect 19886 11132 19892 11144
rect 19392 11104 19892 11132
rect 19392 11092 19398 11104
rect 19886 11092 19892 11104
rect 19944 11092 19950 11144
rect 22097 11135 22155 11141
rect 22097 11101 22109 11135
rect 22143 11132 22155 11135
rect 24118 11132 24124 11144
rect 22143 11104 24124 11132
rect 22143 11101 22155 11104
rect 22097 11095 22155 11101
rect 24118 11092 24124 11104
rect 24176 11092 24182 11144
rect 24394 11132 24400 11144
rect 24355 11104 24400 11132
rect 24394 11092 24400 11104
rect 24452 11092 24458 11144
rect 24664 11135 24722 11141
rect 24664 11101 24676 11135
rect 24710 11132 24722 11135
rect 25498 11132 25504 11144
rect 24710 11104 25504 11132
rect 24710 11101 24722 11104
rect 24664 11095 24722 11101
rect 25498 11092 25504 11104
rect 25556 11092 25562 11144
rect 30561 11135 30619 11141
rect 30561 11101 30573 11135
rect 30607 11101 30619 11135
rect 30561 11095 30619 11101
rect 30828 11135 30886 11141
rect 30828 11101 30840 11135
rect 30874 11132 30886 11135
rect 31202 11132 31208 11144
rect 30874 11104 31208 11132
rect 30874 11101 30886 11104
rect 30828 11095 30886 11101
rect 19242 11064 19248 11076
rect 15304 11036 19248 11064
rect 19242 11024 19248 11036
rect 19300 11024 19306 11076
rect 20156 11067 20214 11073
rect 20156 11033 20168 11067
rect 20202 11064 20214 11067
rect 20990 11064 20996 11076
rect 20202 11036 20996 11064
rect 20202 11033 20214 11036
rect 20156 11027 20214 11033
rect 20990 11024 20996 11036
rect 21048 11024 21054 11076
rect 22364 11067 22422 11073
rect 22364 11033 22376 11067
rect 22410 11064 22422 11067
rect 23198 11064 23204 11076
rect 22410 11036 23204 11064
rect 22410 11033 22422 11036
rect 22364 11027 22422 11033
rect 23198 11024 23204 11036
rect 23256 11024 23262 11076
rect 30576 11064 30604 11095
rect 31202 11092 31208 11104
rect 31260 11092 31266 11144
rect 32401 11135 32459 11141
rect 32401 11101 32413 11135
rect 32447 11101 32459 11135
rect 32401 11095 32459 11101
rect 32668 11135 32726 11141
rect 32668 11101 32680 11135
rect 32714 11132 32726 11135
rect 33502 11132 33508 11144
rect 32714 11104 33508 11132
rect 32714 11101 32726 11104
rect 32668 11095 32726 11101
rect 32122 11064 32128 11076
rect 30576 11036 32128 11064
rect 32122 11024 32128 11036
rect 32180 11024 32186 11076
rect 32416 11064 32444 11095
rect 33502 11092 33508 11104
rect 33560 11092 33566 11144
rect 34701 11135 34759 11141
rect 34701 11101 34713 11135
rect 34747 11101 34759 11135
rect 34701 11095 34759 11101
rect 34968 11135 35026 11141
rect 34968 11101 34980 11135
rect 35014 11132 35026 11135
rect 35342 11132 35348 11144
rect 35014 11104 35348 11132
rect 35014 11101 35026 11104
rect 34968 11095 35026 11101
rect 33410 11064 33416 11076
rect 32416 11036 33416 11064
rect 33410 11024 33416 11036
rect 33468 11064 33474 11076
rect 33962 11064 33968 11076
rect 33468 11036 33968 11064
rect 33468 11024 33474 11036
rect 33962 11024 33968 11036
rect 34020 11064 34026 11076
rect 34716 11064 34744 11095
rect 35342 11092 35348 11104
rect 35400 11092 35406 11144
rect 37369 11135 37427 11141
rect 37369 11101 37381 11135
rect 37415 11132 37427 11135
rect 37458 11132 37464 11144
rect 37415 11104 37464 11132
rect 37415 11101 37427 11104
rect 37369 11095 37427 11101
rect 37458 11092 37464 11104
rect 37516 11092 37522 11144
rect 40037 11135 40095 11141
rect 40037 11101 40049 11135
rect 40083 11132 40095 11135
rect 40402 11132 40408 11144
rect 40083 11104 40408 11132
rect 40083 11101 40095 11104
rect 40037 11095 40095 11101
rect 40402 11092 40408 11104
rect 40460 11092 40466 11144
rect 46652 11135 46710 11141
rect 46652 11101 46664 11135
rect 46698 11132 46710 11135
rect 47762 11132 47768 11144
rect 46698 11104 47768 11132
rect 46698 11101 46710 11104
rect 46652 11095 46710 11101
rect 47762 11092 47768 11104
rect 47820 11092 47826 11144
rect 48225 11135 48283 11141
rect 48225 11101 48237 11135
rect 48271 11101 48283 11135
rect 48225 11095 48283 11101
rect 48492 11135 48550 11141
rect 48492 11101 48504 11135
rect 48538 11132 48550 11135
rect 50062 11132 50068 11144
rect 48538 11104 50068 11132
rect 48538 11101 48550 11104
rect 48492 11095 48550 11101
rect 34020 11036 34744 11064
rect 37636 11067 37694 11073
rect 34020 11024 34026 11036
rect 37636 11033 37648 11067
rect 37682 11064 37694 11067
rect 38654 11064 38660 11076
rect 37682 11036 38660 11064
rect 37682 11033 37694 11036
rect 37636 11027 37694 11033
rect 38654 11024 38660 11036
rect 38712 11024 38718 11076
rect 40764 11067 40822 11073
rect 40764 11033 40776 11067
rect 40810 11064 40822 11067
rect 41782 11064 41788 11076
rect 40810 11036 41788 11064
rect 40810 11033 40822 11036
rect 40764 11027 40822 11033
rect 41782 11024 41788 11036
rect 41840 11024 41846 11076
rect 45830 11024 45836 11076
rect 45888 11064 45894 11076
rect 48240 11064 48268 11095
rect 50062 11092 50068 11104
rect 50120 11092 50126 11144
rect 51537 11135 51595 11141
rect 51537 11101 51549 11135
rect 51583 11132 51595 11135
rect 53282 11132 53288 11144
rect 51583 11104 53288 11132
rect 51583 11101 51595 11104
rect 51537 11095 51595 11101
rect 53282 11092 53288 11104
rect 53340 11092 53346 11144
rect 53644 11135 53702 11141
rect 53644 11101 53656 11135
rect 53690 11132 53702 11135
rect 54386 11132 54392 11144
rect 53690 11104 54392 11132
rect 53690 11101 53702 11104
rect 53644 11095 53702 11101
rect 54386 11092 54392 11104
rect 54444 11092 54450 11144
rect 48590 11064 48596 11076
rect 45888 11036 48596 11064
rect 45888 11024 45894 11036
rect 48590 11024 48596 11036
rect 48648 11024 48654 11076
rect 51804 11067 51862 11073
rect 51804 11033 51816 11067
rect 51850 11064 51862 11067
rect 53742 11064 53748 11076
rect 51850 11036 53748 11064
rect 51850 11033 51862 11036
rect 51804 11027 51862 11033
rect 53742 11024 53748 11036
rect 53800 11024 53806 11076
rect 57140 11067 57198 11073
rect 57140 11033 57152 11067
rect 57186 11064 57198 11067
rect 57330 11064 57336 11076
rect 57186 11036 57336 11064
rect 57186 11033 57198 11036
rect 57140 11027 57198 11033
rect 57330 11024 57336 11036
rect 57388 11024 57394 11076
rect 10778 10996 10784 11008
rect 10739 10968 10784 10996
rect 10778 10956 10784 10968
rect 10836 10956 10842 11008
rect 25774 10996 25780 11008
rect 25735 10968 25780 10996
rect 25774 10956 25780 10968
rect 25832 10956 25838 11008
rect 47762 10996 47768 11008
rect 47723 10968 47768 10996
rect 47762 10956 47768 10968
rect 47820 10956 47826 11008
rect 54754 10996 54760 11008
rect 54715 10968 54760 10996
rect 54754 10956 54760 10968
rect 54812 10956 54818 11008
rect 58250 10996 58256 11008
rect 58211 10968 58256 10996
rect 58250 10956 58256 10968
rect 58308 10956 58314 11008
rect 1104 10906 59340 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 59340 10906
rect 1104 10832 59340 10854
rect 15194 10752 15200 10804
rect 15252 10792 15258 10804
rect 15473 10795 15531 10801
rect 15473 10792 15485 10795
rect 15252 10764 15485 10792
rect 15252 10752 15258 10764
rect 15473 10761 15485 10764
rect 15519 10761 15531 10795
rect 20990 10792 20996 10804
rect 20951 10764 20996 10792
rect 15473 10755 15531 10761
rect 20990 10752 20996 10764
rect 21048 10752 21054 10804
rect 23198 10792 23204 10804
rect 23159 10764 23204 10792
rect 23198 10752 23204 10764
rect 23256 10752 23262 10804
rect 33686 10752 33692 10804
rect 33744 10792 33750 10804
rect 33781 10795 33839 10801
rect 33781 10792 33793 10795
rect 33744 10764 33793 10792
rect 33744 10752 33750 10764
rect 33781 10761 33793 10764
rect 33827 10761 33839 10795
rect 38654 10792 38660 10804
rect 38615 10764 38660 10792
rect 33781 10755 33839 10761
rect 38654 10752 38660 10764
rect 38712 10752 38718 10804
rect 41782 10752 41788 10804
rect 41840 10792 41846 10804
rect 41877 10795 41935 10801
rect 41877 10792 41889 10795
rect 41840 10764 41889 10792
rect 41840 10752 41846 10764
rect 41877 10761 41889 10764
rect 41923 10761 41935 10795
rect 47029 10795 47087 10801
rect 47029 10792 47041 10795
rect 41877 10755 41935 10761
rect 45526 10764 47041 10792
rect 9576 10727 9634 10733
rect 9576 10693 9588 10727
rect 9622 10724 9634 10727
rect 10778 10724 10784 10736
rect 9622 10696 10784 10724
rect 9622 10693 9634 10696
rect 9576 10687 9634 10693
rect 10778 10684 10784 10696
rect 10836 10684 10842 10736
rect 14090 10684 14096 10736
rect 14148 10724 14154 10736
rect 14338 10727 14396 10733
rect 14338 10724 14350 10727
rect 14148 10696 14350 10724
rect 14148 10684 14154 10696
rect 14338 10693 14350 10696
rect 14384 10693 14396 10727
rect 14338 10687 14396 10693
rect 16936 10727 16994 10733
rect 16936 10693 16948 10727
rect 16982 10724 16994 10727
rect 18046 10724 18052 10736
rect 16982 10696 18052 10724
rect 16982 10693 16994 10696
rect 16936 10687 16994 10693
rect 18046 10684 18052 10696
rect 18104 10684 18110 10736
rect 19242 10684 19248 10736
rect 19300 10724 19306 10736
rect 20898 10724 20904 10736
rect 19300 10696 20904 10724
rect 19300 10684 19306 10696
rect 20898 10684 20904 10696
rect 20956 10684 20962 10736
rect 22094 10733 22100 10736
rect 22088 10724 22100 10733
rect 22055 10696 22100 10724
rect 22088 10687 22100 10696
rect 22094 10684 22100 10687
rect 22152 10684 22158 10736
rect 24296 10727 24354 10733
rect 24296 10693 24308 10727
rect 24342 10724 24354 10727
rect 25774 10724 25780 10736
rect 24342 10696 25780 10724
rect 24342 10693 24354 10696
rect 24296 10687 24354 10693
rect 25774 10684 25780 10696
rect 25832 10684 25838 10736
rect 29546 10724 29552 10736
rect 27632 10696 29552 10724
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10656 9367 10659
rect 9858 10656 9864 10668
rect 9355 10628 9864 10656
rect 9355 10625 9367 10628
rect 9309 10619 9367 10625
rect 9858 10616 9864 10628
rect 9916 10616 9922 10668
rect 11790 10665 11796 10668
rect 11784 10619 11796 10665
rect 11848 10656 11854 10668
rect 16669 10659 16727 10665
rect 11848 10628 11884 10656
rect 11790 10616 11796 10619
rect 11848 10616 11854 10628
rect 16669 10625 16681 10659
rect 16715 10656 16727 10659
rect 16758 10656 16764 10668
rect 16715 10628 16764 10656
rect 16715 10625 16727 10628
rect 16669 10619 16727 10625
rect 16758 10616 16764 10628
rect 16816 10616 16822 10668
rect 19161 10659 19219 10665
rect 19161 10625 19173 10659
rect 19207 10656 19219 10659
rect 19260 10656 19288 10684
rect 19207 10628 19288 10656
rect 19880 10659 19938 10665
rect 19207 10625 19219 10628
rect 19161 10619 19219 10625
rect 19880 10625 19892 10659
rect 19926 10656 19938 10659
rect 20714 10656 20720 10668
rect 19926 10628 20720 10656
rect 19926 10625 19938 10628
rect 19880 10619 19938 10625
rect 20714 10616 20720 10628
rect 20772 10616 20778 10668
rect 24029 10659 24087 10665
rect 24029 10625 24041 10659
rect 24075 10656 24087 10659
rect 24118 10656 24124 10668
rect 24075 10628 24124 10656
rect 24075 10625 24087 10628
rect 24029 10619 24087 10625
rect 24118 10616 24124 10628
rect 24176 10616 24182 10668
rect 27522 10616 27528 10668
rect 27580 10656 27586 10668
rect 27632 10665 27660 10696
rect 29546 10684 29552 10696
rect 29604 10684 29610 10736
rect 32668 10727 32726 10733
rect 32668 10693 32680 10727
rect 32714 10724 32726 10727
rect 34146 10724 34152 10736
rect 32714 10696 34152 10724
rect 32714 10693 32726 10696
rect 32668 10687 32726 10693
rect 34146 10684 34152 10696
rect 34204 10684 34210 10736
rect 34508 10727 34566 10733
rect 34508 10693 34520 10727
rect 34554 10724 34566 10727
rect 36078 10724 36084 10736
rect 34554 10696 36084 10724
rect 34554 10693 34566 10696
rect 34508 10687 34566 10693
rect 36078 10684 36084 10696
rect 36136 10684 36142 10736
rect 44076 10727 44134 10733
rect 44076 10693 44088 10727
rect 44122 10724 44134 10727
rect 45526 10724 45554 10764
rect 47029 10761 47041 10764
rect 47075 10761 47087 10795
rect 47029 10755 47087 10761
rect 48130 10752 48136 10804
rect 48188 10792 48194 10804
rect 48225 10795 48283 10801
rect 48225 10792 48237 10795
rect 48188 10764 48237 10792
rect 48188 10752 48194 10764
rect 48225 10761 48237 10764
rect 48271 10761 48283 10795
rect 48225 10755 48283 10761
rect 50341 10795 50399 10801
rect 50341 10761 50353 10795
rect 50387 10792 50399 10795
rect 50614 10792 50620 10804
rect 50387 10764 50620 10792
rect 50387 10761 50399 10764
rect 50341 10755 50399 10761
rect 50614 10752 50620 10764
rect 50672 10752 50678 10804
rect 51074 10752 51080 10804
rect 51132 10752 51138 10804
rect 55490 10792 55496 10804
rect 55451 10764 55496 10792
rect 55490 10752 55496 10764
rect 55548 10752 55554 10804
rect 57238 10752 57244 10804
rect 57296 10792 57302 10804
rect 57333 10795 57391 10801
rect 57333 10792 57345 10795
rect 57296 10764 57345 10792
rect 57296 10752 57302 10764
rect 57333 10761 57345 10764
rect 57379 10761 57391 10795
rect 57333 10755 57391 10761
rect 44122 10696 45554 10724
rect 45916 10727 45974 10733
rect 44122 10693 44134 10696
rect 44076 10687 44134 10693
rect 45916 10693 45928 10727
rect 45962 10724 45974 10727
rect 47762 10724 47768 10736
rect 45962 10696 47768 10724
rect 45962 10693 45974 10696
rect 45916 10687 45974 10693
rect 47762 10684 47768 10696
rect 47820 10684 47826 10736
rect 51092 10724 51120 10752
rect 50816 10696 51120 10724
rect 54380 10727 54438 10733
rect 27617 10659 27675 10665
rect 27617 10656 27629 10659
rect 27580 10628 27629 10656
rect 27580 10616 27586 10628
rect 27617 10625 27629 10628
rect 27663 10625 27675 10659
rect 27617 10619 27675 10625
rect 27884 10659 27942 10665
rect 27884 10625 27896 10659
rect 27930 10656 27942 10659
rect 30190 10656 30196 10668
rect 27930 10628 30196 10656
rect 27930 10625 27942 10628
rect 27884 10619 27942 10625
rect 30190 10616 30196 10628
rect 30248 10616 30254 10668
rect 32122 10616 32128 10668
rect 32180 10656 32186 10668
rect 32401 10659 32459 10665
rect 32401 10656 32413 10659
rect 32180 10628 32413 10656
rect 32180 10616 32186 10628
rect 32401 10625 32413 10628
rect 32447 10625 32459 10659
rect 32401 10619 32459 10625
rect 37544 10659 37602 10665
rect 37544 10625 37556 10659
rect 37590 10656 37602 10659
rect 38562 10656 38568 10668
rect 37590 10628 38568 10656
rect 37590 10625 37602 10628
rect 37544 10619 37602 10625
rect 38562 10616 38568 10628
rect 38620 10616 38626 10668
rect 40494 10656 40500 10668
rect 40455 10628 40500 10656
rect 40494 10616 40500 10628
rect 40552 10616 40558 10668
rect 40764 10659 40822 10665
rect 40764 10625 40776 10659
rect 40810 10656 40822 10659
rect 41874 10656 41880 10668
rect 40810 10628 41880 10656
rect 40810 10625 40822 10628
rect 40764 10619 40822 10625
rect 41874 10616 41880 10628
rect 41932 10616 41938 10668
rect 43809 10659 43867 10665
rect 43809 10625 43821 10659
rect 43855 10656 43867 10659
rect 45649 10659 45707 10665
rect 45649 10656 45661 10659
rect 43855 10628 45661 10656
rect 43855 10625 43867 10628
rect 43809 10619 43867 10625
rect 45649 10625 45661 10628
rect 45695 10656 45707 10659
rect 45738 10656 45744 10668
rect 45695 10628 45744 10656
rect 45695 10625 45707 10628
rect 45649 10619 45707 10625
rect 45738 10616 45744 10628
rect 45796 10616 45802 10668
rect 48406 10656 48412 10668
rect 48367 10628 48412 10656
rect 48406 10616 48412 10628
rect 48464 10616 48470 10668
rect 49228 10659 49286 10665
rect 49228 10625 49240 10659
rect 49274 10656 49286 10659
rect 50154 10656 50160 10668
rect 49274 10628 50160 10656
rect 49274 10625 49286 10628
rect 49228 10619 49286 10625
rect 50154 10616 50160 10628
rect 50212 10616 50218 10668
rect 50816 10665 50844 10696
rect 54380 10693 54392 10727
rect 54426 10724 54438 10727
rect 55950 10724 55956 10736
rect 54426 10696 55956 10724
rect 54426 10693 54438 10696
rect 54380 10687 54438 10693
rect 55950 10684 55956 10696
rect 56008 10684 56014 10736
rect 56220 10727 56278 10733
rect 56220 10693 56232 10727
rect 56266 10724 56278 10727
rect 58250 10724 58256 10736
rect 56266 10696 58256 10724
rect 56266 10693 56278 10696
rect 56220 10687 56278 10693
rect 58250 10684 58256 10696
rect 58308 10684 58314 10736
rect 50801 10659 50859 10665
rect 50801 10625 50813 10659
rect 50847 10625 50859 10659
rect 50801 10619 50859 10625
rect 51068 10659 51126 10665
rect 51068 10625 51080 10659
rect 51114 10656 51126 10659
rect 52914 10656 52920 10668
rect 51114 10628 52920 10656
rect 51114 10625 51126 10628
rect 51068 10619 51126 10625
rect 52914 10616 52920 10628
rect 52972 10616 52978 10668
rect 53282 10616 53288 10668
rect 53340 10656 53346 10668
rect 54113 10659 54171 10665
rect 54113 10656 54125 10659
rect 53340 10628 54125 10656
rect 53340 10616 53346 10628
rect 54113 10625 54125 10628
rect 54159 10656 54171 10659
rect 54159 10628 55996 10656
rect 54159 10625 54171 10628
rect 54113 10619 54171 10625
rect 10778 10548 10784 10600
rect 10836 10588 10842 10600
rect 11517 10591 11575 10597
rect 11517 10588 11529 10591
rect 10836 10560 11529 10588
rect 10836 10548 10842 10560
rect 11517 10557 11529 10560
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 13814 10548 13820 10600
rect 13872 10588 13878 10600
rect 14093 10591 14151 10597
rect 14093 10588 14105 10591
rect 13872 10560 14105 10588
rect 13872 10548 13878 10560
rect 14093 10557 14105 10560
rect 14139 10557 14151 10591
rect 14093 10551 14151 10557
rect 19334 10548 19340 10600
rect 19392 10588 19398 10600
rect 19613 10591 19671 10597
rect 19613 10588 19625 10591
rect 19392 10560 19625 10588
rect 19392 10548 19398 10560
rect 19613 10557 19625 10560
rect 19659 10557 19671 10591
rect 19613 10551 19671 10557
rect 20622 10548 20628 10600
rect 20680 10588 20686 10600
rect 21821 10591 21879 10597
rect 21821 10588 21833 10591
rect 20680 10560 21833 10588
rect 20680 10548 20686 10560
rect 21821 10557 21833 10560
rect 21867 10557 21879 10591
rect 21821 10551 21879 10557
rect 33410 10548 33416 10600
rect 33468 10588 33474 10600
rect 34241 10591 34299 10597
rect 34241 10588 34253 10591
rect 33468 10560 34253 10588
rect 33468 10548 33474 10560
rect 34241 10557 34253 10560
rect 34287 10557 34299 10591
rect 37274 10588 37280 10600
rect 37235 10560 37280 10588
rect 34241 10551 34299 10557
rect 37274 10548 37280 10560
rect 37332 10548 37338 10600
rect 48958 10588 48964 10600
rect 48919 10560 48964 10588
rect 48958 10548 48964 10560
rect 49016 10548 49022 10600
rect 55968 10597 55996 10628
rect 55953 10591 56011 10597
rect 55953 10557 55965 10591
rect 55999 10557 56011 10591
rect 55953 10551 56011 10557
rect 10686 10452 10692 10464
rect 10647 10424 10692 10452
rect 10686 10412 10692 10424
rect 10744 10412 10750 10464
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10452 12955 10455
rect 14366 10452 14372 10464
rect 12943 10424 14372 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 14366 10412 14372 10424
rect 14424 10412 14430 10464
rect 18046 10452 18052 10464
rect 18007 10424 18052 10452
rect 18046 10412 18052 10424
rect 18104 10412 18110 10464
rect 18598 10412 18604 10464
rect 18656 10452 18662 10464
rect 18969 10455 19027 10461
rect 18969 10452 18981 10455
rect 18656 10424 18981 10452
rect 18656 10412 18662 10424
rect 18969 10421 18981 10424
rect 19015 10421 19027 10455
rect 25406 10452 25412 10464
rect 25367 10424 25412 10452
rect 18969 10415 19027 10421
rect 25406 10412 25412 10424
rect 25464 10412 25470 10464
rect 28997 10455 29055 10461
rect 28997 10421 29009 10455
rect 29043 10452 29055 10455
rect 29822 10452 29828 10464
rect 29043 10424 29828 10452
rect 29043 10421 29055 10424
rect 28997 10415 29055 10421
rect 29822 10412 29828 10424
rect 29880 10412 29886 10464
rect 35618 10452 35624 10464
rect 35579 10424 35624 10452
rect 35618 10412 35624 10424
rect 35676 10412 35682 10464
rect 43346 10412 43352 10464
rect 43404 10452 43410 10464
rect 45189 10455 45247 10461
rect 45189 10452 45201 10455
rect 43404 10424 45201 10452
rect 43404 10412 43410 10424
rect 45189 10421 45201 10424
rect 45235 10421 45247 10455
rect 52178 10452 52184 10464
rect 52139 10424 52184 10452
rect 45189 10415 45247 10421
rect 52178 10412 52184 10424
rect 52236 10412 52242 10464
rect 55968 10452 55996 10551
rect 56870 10452 56876 10464
rect 55968 10424 56876 10452
rect 56870 10412 56876 10424
rect 56928 10412 56934 10464
rect 1104 10362 59340 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 59340 10362
rect 1104 10288 59340 10310
rect 9858 10248 9864 10260
rect 9140 10220 9864 10248
rect 6086 10112 6092 10124
rect 6047 10084 6092 10112
rect 6086 10072 6092 10084
rect 6144 10072 6150 10124
rect 9030 10072 9036 10124
rect 9088 10112 9094 10124
rect 9140 10121 9168 10220
rect 9858 10208 9864 10220
rect 9916 10208 9922 10260
rect 13906 10208 13912 10260
rect 13964 10248 13970 10260
rect 16117 10251 16175 10257
rect 16117 10248 16129 10251
rect 13964 10220 16129 10248
rect 13964 10208 13970 10220
rect 16117 10217 16129 10220
rect 16163 10217 16175 10251
rect 17954 10248 17960 10260
rect 17915 10220 17960 10248
rect 16117 10211 16175 10217
rect 17954 10208 17960 10220
rect 18012 10208 18018 10260
rect 19334 10208 19340 10260
rect 19392 10248 19398 10260
rect 20622 10248 20628 10260
rect 19392 10220 20628 10248
rect 19392 10208 19398 10220
rect 20622 10208 20628 10220
rect 20680 10248 20686 10260
rect 20901 10251 20959 10257
rect 20901 10248 20913 10251
rect 20680 10220 20913 10248
rect 20680 10208 20686 10220
rect 20901 10217 20913 10220
rect 20947 10217 20959 10251
rect 26234 10248 26240 10260
rect 20901 10211 20959 10217
rect 21008 10220 26240 10248
rect 21008 10180 21036 10220
rect 26234 10208 26240 10220
rect 26292 10208 26298 10260
rect 37458 10248 37464 10260
rect 37200 10220 37464 10248
rect 19628 10152 21036 10180
rect 9125 10115 9183 10121
rect 9125 10112 9137 10115
rect 9088 10084 9137 10112
rect 9088 10072 9094 10084
rect 9125 10081 9137 10084
rect 9171 10081 9183 10115
rect 10962 10112 10968 10124
rect 10923 10084 10968 10112
rect 9125 10075 9183 10081
rect 10962 10072 10968 10084
rect 11020 10072 11026 10124
rect 9392 10047 9450 10053
rect 9392 10013 9404 10047
rect 9438 10044 9450 10047
rect 10686 10044 10692 10056
rect 9438 10016 10692 10044
rect 9438 10013 9450 10016
rect 9392 10007 9450 10013
rect 10686 10004 10692 10016
rect 10744 10004 10750 10056
rect 14090 10004 14096 10056
rect 14148 10044 14154 10056
rect 14737 10047 14795 10053
rect 14737 10044 14749 10047
rect 14148 10016 14749 10044
rect 14148 10004 14154 10016
rect 14737 10013 14749 10016
rect 14783 10013 14795 10047
rect 14737 10007 14795 10013
rect 16577 10047 16635 10053
rect 16577 10013 16589 10047
rect 16623 10044 16635 10047
rect 16666 10044 16672 10056
rect 16623 10016 16672 10044
rect 16623 10013 16635 10016
rect 16577 10007 16635 10013
rect 16666 10004 16672 10016
rect 16724 10004 16730 10056
rect 16844 10047 16902 10053
rect 16844 10013 16856 10047
rect 16890 10044 16902 10047
rect 18046 10044 18052 10056
rect 16890 10016 18052 10044
rect 16890 10013 16902 10016
rect 16844 10007 16902 10013
rect 18046 10004 18052 10016
rect 18104 10004 18110 10056
rect 18598 10004 18604 10056
rect 18656 10044 18662 10056
rect 19426 10044 19432 10056
rect 18656 10016 19432 10044
rect 18656 10004 18662 10016
rect 19426 10004 19432 10016
rect 19484 10044 19490 10056
rect 19628 10053 19656 10152
rect 28445 10115 28503 10121
rect 28445 10081 28457 10115
rect 28491 10112 28503 10115
rect 29546 10112 29552 10124
rect 28491 10084 29552 10112
rect 28491 10081 28503 10084
rect 28445 10075 28503 10081
rect 29546 10072 29552 10084
rect 29604 10072 29610 10124
rect 37200 10121 37228 10220
rect 37458 10208 37464 10220
rect 37516 10208 37522 10260
rect 38562 10248 38568 10260
rect 38523 10220 38568 10248
rect 38562 10208 38568 10220
rect 38620 10208 38626 10260
rect 44453 10251 44511 10257
rect 44453 10217 44465 10251
rect 44499 10248 44511 10251
rect 47854 10248 47860 10260
rect 44499 10220 47860 10248
rect 44499 10217 44511 10220
rect 44453 10211 44511 10217
rect 47854 10208 47860 10220
rect 47912 10208 47918 10260
rect 48590 10248 48596 10260
rect 48551 10220 48596 10248
rect 48590 10208 48596 10220
rect 48648 10208 48654 10260
rect 52914 10248 52920 10260
rect 52875 10220 52920 10248
rect 52914 10208 52920 10220
rect 52972 10208 52978 10260
rect 53742 10208 53748 10260
rect 53800 10248 53806 10260
rect 54757 10251 54815 10257
rect 54757 10248 54769 10251
rect 53800 10220 54769 10248
rect 53800 10208 53806 10220
rect 54757 10217 54769 10220
rect 54803 10217 54815 10251
rect 54757 10211 54815 10217
rect 37185 10115 37243 10121
rect 37185 10081 37197 10115
rect 37231 10081 37243 10115
rect 37185 10075 37243 10081
rect 53282 10072 53288 10124
rect 53340 10112 53346 10124
rect 53377 10115 53435 10121
rect 53377 10112 53389 10115
rect 53340 10084 53389 10112
rect 53340 10072 53346 10084
rect 53377 10081 53389 10084
rect 53423 10081 53435 10115
rect 56870 10112 56876 10124
rect 56831 10084 56876 10112
rect 53377 10075 53435 10081
rect 56870 10072 56876 10084
rect 56928 10072 56934 10124
rect 19613 10047 19671 10053
rect 19613 10044 19625 10047
rect 19484 10016 19625 10044
rect 19484 10004 19490 10016
rect 19613 10013 19625 10016
rect 19659 10013 19671 10047
rect 24394 10044 24400 10056
rect 24355 10016 24400 10044
rect 19613 10007 19671 10013
rect 24394 10004 24400 10016
rect 24452 10004 24458 10056
rect 24664 10047 24722 10053
rect 24664 10013 24676 10047
rect 24710 10044 24722 10047
rect 25406 10044 25412 10056
rect 24710 10016 25412 10044
rect 24710 10013 24722 10016
rect 24664 10007 24722 10013
rect 25406 10004 25412 10016
rect 25464 10004 25470 10056
rect 26234 10004 26240 10056
rect 26292 10044 26298 10056
rect 26697 10047 26755 10053
rect 26697 10044 26709 10047
rect 26292 10016 26709 10044
rect 26292 10004 26298 10016
rect 26697 10013 26709 10016
rect 26743 10013 26755 10047
rect 26697 10007 26755 10013
rect 32769 10047 32827 10053
rect 32769 10013 32781 10047
rect 32815 10044 32827 10047
rect 33410 10044 33416 10056
rect 32815 10016 33416 10044
rect 32815 10013 32827 10016
rect 32769 10007 32827 10013
rect 33410 10004 33416 10016
rect 33468 10004 33474 10056
rect 43073 10047 43131 10053
rect 43073 10013 43085 10047
rect 43119 10044 43131 10047
rect 45005 10047 45063 10053
rect 45005 10044 45017 10047
rect 43119 10016 45017 10044
rect 43119 10013 43131 10016
rect 43073 10007 43131 10013
rect 45005 10013 45017 10016
rect 45051 10044 45063 10047
rect 45738 10044 45744 10056
rect 45051 10016 45744 10044
rect 45051 10013 45063 10016
rect 45005 10007 45063 10013
rect 45738 10004 45744 10016
rect 45796 10004 45802 10056
rect 47305 10047 47363 10053
rect 47305 10013 47317 10047
rect 47351 10044 47363 10047
rect 48130 10044 48136 10056
rect 47351 10016 48136 10044
rect 47351 10013 47363 10016
rect 47305 10007 47363 10013
rect 48130 10004 48136 10016
rect 48188 10004 48194 10056
rect 51534 10044 51540 10056
rect 51495 10016 51540 10044
rect 51534 10004 51540 10016
rect 51592 10004 51598 10056
rect 53644 10047 53702 10053
rect 53644 10013 53656 10047
rect 53690 10044 53702 10047
rect 54754 10044 54760 10056
rect 53690 10016 54760 10044
rect 53690 10013 53702 10016
rect 53644 10007 53702 10013
rect 54754 10004 54760 10016
rect 54812 10004 54818 10056
rect 6356 9979 6414 9985
rect 6356 9945 6368 9979
rect 6402 9976 6414 9979
rect 7282 9976 7288 9988
rect 6402 9948 7288 9976
rect 6402 9945 6414 9948
rect 6356 9939 6414 9945
rect 7282 9936 7288 9948
rect 7340 9936 7346 9988
rect 11054 9936 11060 9988
rect 11112 9976 11118 9988
rect 11210 9979 11268 9985
rect 11210 9976 11222 9979
rect 11112 9948 11222 9976
rect 11112 9936 11118 9948
rect 11210 9945 11222 9948
rect 11256 9945 11268 9979
rect 11210 9939 11268 9945
rect 15004 9979 15062 9985
rect 15004 9945 15016 9979
rect 15050 9976 15062 9979
rect 15470 9976 15476 9988
rect 15050 9948 15476 9976
rect 15050 9945 15062 9948
rect 15004 9939 15062 9945
rect 15470 9936 15476 9948
rect 15528 9936 15534 9988
rect 29816 9979 29874 9985
rect 29816 9945 29828 9979
rect 29862 9976 29874 9979
rect 30834 9976 30840 9988
rect 29862 9948 30840 9976
rect 29862 9945 29874 9948
rect 29816 9939 29874 9945
rect 30834 9936 30840 9948
rect 30892 9936 30898 9988
rect 33036 9979 33094 9985
rect 33036 9945 33048 9979
rect 33082 9976 33094 9979
rect 34054 9976 34060 9988
rect 33082 9948 34060 9976
rect 33082 9945 33094 9948
rect 33036 9939 33094 9945
rect 34054 9936 34060 9948
rect 34112 9936 34118 9988
rect 37452 9979 37510 9985
rect 37452 9945 37464 9979
rect 37498 9976 37510 9979
rect 38654 9976 38660 9988
rect 37498 9948 38660 9976
rect 37498 9945 37510 9948
rect 37452 9939 37510 9945
rect 38654 9936 38660 9948
rect 38712 9936 38718 9988
rect 43346 9985 43352 9988
rect 43340 9976 43352 9985
rect 43307 9948 43352 9976
rect 43340 9939 43352 9948
rect 43346 9936 43352 9939
rect 43404 9936 43410 9988
rect 45272 9979 45330 9985
rect 45272 9945 45284 9979
rect 45318 9976 45330 9979
rect 45646 9976 45652 9988
rect 45318 9948 45652 9976
rect 45318 9945 45330 9948
rect 45272 9939 45330 9945
rect 45646 9936 45652 9948
rect 45704 9936 45710 9988
rect 51804 9979 51862 9985
rect 51804 9945 51816 9979
rect 51850 9976 51862 9979
rect 53742 9976 53748 9988
rect 51850 9948 53748 9976
rect 51850 9945 51862 9948
rect 51804 9939 51862 9945
rect 53742 9936 53748 9948
rect 53800 9936 53806 9988
rect 57140 9979 57198 9985
rect 57140 9945 57152 9979
rect 57186 9976 57198 9979
rect 59449 9979 59507 9985
rect 59449 9976 59461 9979
rect 57186 9948 59461 9976
rect 57186 9945 57198 9948
rect 57140 9939 57198 9945
rect 59449 9945 59461 9948
rect 59495 9945 59507 9979
rect 59449 9939 59507 9945
rect 7466 9908 7472 9920
rect 7427 9880 7472 9908
rect 7466 9868 7472 9880
rect 7524 9868 7530 9920
rect 10502 9908 10508 9920
rect 10463 9880 10508 9908
rect 10502 9868 10508 9880
rect 10560 9868 10566 9920
rect 10594 9868 10600 9920
rect 10652 9908 10658 9920
rect 12345 9911 12403 9917
rect 12345 9908 12357 9911
rect 10652 9880 12357 9908
rect 10652 9868 10658 9880
rect 12345 9877 12357 9880
rect 12391 9877 12403 9911
rect 12345 9871 12403 9877
rect 25130 9868 25136 9920
rect 25188 9908 25194 9920
rect 25777 9911 25835 9917
rect 25777 9908 25789 9911
rect 25188 9880 25789 9908
rect 25188 9868 25194 9880
rect 25777 9877 25789 9880
rect 25823 9877 25835 9911
rect 25777 9871 25835 9877
rect 30929 9911 30987 9917
rect 30929 9877 30941 9911
rect 30975 9908 30987 9911
rect 32214 9908 32220 9920
rect 30975 9880 32220 9908
rect 30975 9877 30987 9880
rect 30929 9871 30987 9877
rect 32214 9868 32220 9880
rect 32272 9868 32278 9920
rect 34146 9908 34152 9920
rect 34107 9880 34152 9908
rect 34146 9868 34152 9880
rect 34204 9868 34210 9920
rect 45370 9868 45376 9920
rect 45428 9908 45434 9920
rect 46385 9911 46443 9917
rect 46385 9908 46397 9911
rect 45428 9880 46397 9908
rect 45428 9868 45434 9880
rect 46385 9877 46397 9880
rect 46431 9877 46443 9911
rect 58250 9908 58256 9920
rect 58211 9880 58256 9908
rect 46385 9871 46443 9877
rect 58250 9868 58256 9880
rect 58308 9868 58314 9920
rect 1104 9818 59340 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 59340 9818
rect 1104 9744 59340 9766
rect 20714 9704 20720 9716
rect 20675 9676 20720 9704
rect 20714 9664 20720 9676
rect 20772 9664 20778 9716
rect 30190 9704 30196 9716
rect 30151 9676 30196 9704
rect 30190 9664 30196 9676
rect 30248 9664 30254 9716
rect 38654 9704 38660 9716
rect 38615 9676 38660 9704
rect 38654 9664 38660 9676
rect 38712 9664 38718 9716
rect 41874 9704 41880 9716
rect 41835 9676 41880 9704
rect 41874 9664 41880 9676
rect 41932 9664 41938 9716
rect 45646 9704 45652 9716
rect 45607 9676 45652 9704
rect 45646 9664 45652 9676
rect 45704 9664 45710 9716
rect 50154 9664 50160 9716
rect 50212 9704 50218 9716
rect 50341 9707 50399 9713
rect 50341 9704 50353 9707
rect 50212 9676 50353 9704
rect 50212 9664 50218 9676
rect 50341 9673 50353 9676
rect 50387 9673 50399 9707
rect 50341 9667 50399 9673
rect 6632 9639 6690 9645
rect 6632 9605 6644 9639
rect 6678 9636 6690 9639
rect 9300 9639 9358 9645
rect 6678 9608 6914 9636
rect 6678 9605 6690 9608
rect 6632 9599 6690 9605
rect 6886 9568 6914 9608
rect 9300 9605 9312 9639
rect 9346 9636 9358 9639
rect 10502 9636 10508 9648
rect 9346 9608 10508 9636
rect 9346 9605 9358 9608
rect 9300 9599 9358 9605
rect 10502 9596 10508 9608
rect 10560 9596 10566 9648
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 12897 9639 12955 9645
rect 12897 9636 12909 9639
rect 12492 9608 12909 9636
rect 12492 9596 12498 9608
rect 12897 9605 12909 9608
rect 12943 9605 12955 9639
rect 12897 9599 12955 9605
rect 16936 9639 16994 9645
rect 16936 9605 16948 9639
rect 16982 9636 16994 9639
rect 18138 9636 18144 9648
rect 16982 9608 18144 9636
rect 16982 9605 16994 9608
rect 16936 9599 16994 9605
rect 18138 9596 18144 9608
rect 18196 9596 18202 9648
rect 24394 9636 24400 9648
rect 23216 9608 24400 9636
rect 12802 9568 12808 9580
rect 6886 9540 12808 9568
rect 12802 9528 12808 9540
rect 12860 9528 12866 9580
rect 16666 9568 16672 9580
rect 16627 9540 16672 9568
rect 16666 9528 16672 9540
rect 16724 9528 16730 9580
rect 19604 9571 19662 9577
rect 19604 9537 19616 9571
rect 19650 9568 19662 9571
rect 20530 9568 20536 9580
rect 19650 9540 20536 9568
rect 19650 9537 19662 9540
rect 19604 9531 19662 9537
rect 20530 9528 20536 9540
rect 20588 9528 20594 9580
rect 23216 9577 23244 9608
rect 24394 9596 24400 9608
rect 24452 9636 24458 9648
rect 26234 9636 26240 9648
rect 24452 9608 26240 9636
rect 24452 9596 24458 9608
rect 23201 9571 23259 9577
rect 23201 9537 23213 9571
rect 23247 9537 23259 9571
rect 23201 9531 23259 9537
rect 23468 9571 23526 9577
rect 23468 9537 23480 9571
rect 23514 9568 23526 9571
rect 24946 9568 24952 9580
rect 23514 9540 24952 9568
rect 23514 9537 23526 9540
rect 23468 9531 23526 9537
rect 24946 9528 24952 9540
rect 25004 9528 25010 9580
rect 25056 9577 25084 9608
rect 26234 9596 26240 9608
rect 26292 9636 26298 9648
rect 27522 9636 27528 9648
rect 26292 9608 27528 9636
rect 26292 9596 26298 9608
rect 25041 9571 25099 9577
rect 25041 9537 25053 9571
rect 25087 9537 25099 9571
rect 25041 9531 25099 9537
rect 25308 9571 25366 9577
rect 25308 9537 25320 9571
rect 25354 9568 25366 9571
rect 25774 9568 25780 9580
rect 25354 9540 25780 9568
rect 25354 9537 25366 9540
rect 25308 9531 25366 9537
rect 25774 9528 25780 9540
rect 25832 9528 25838 9580
rect 26988 9577 27016 9608
rect 27522 9596 27528 9608
rect 27580 9596 27586 9648
rect 34048 9639 34106 9645
rect 34048 9605 34060 9639
rect 34094 9636 34106 9639
rect 35618 9636 35624 9648
rect 34094 9608 35624 9636
rect 34094 9605 34106 9608
rect 34048 9599 34106 9605
rect 35618 9596 35624 9608
rect 35676 9596 35682 9648
rect 49228 9639 49286 9645
rect 37292 9608 44312 9636
rect 37292 9580 37320 9608
rect 40512 9580 40540 9608
rect 26973 9571 27031 9577
rect 26973 9537 26985 9571
rect 27019 9537 27031 9571
rect 26973 9531 27031 9537
rect 27240 9571 27298 9577
rect 27240 9537 27252 9571
rect 27286 9568 27298 9571
rect 27614 9568 27620 9580
rect 27286 9540 27620 9568
rect 27286 9537 27298 9540
rect 27240 9531 27298 9537
rect 27614 9528 27620 9540
rect 27672 9528 27678 9580
rect 29086 9577 29092 9580
rect 29080 9531 29092 9577
rect 29144 9568 29150 9580
rect 37274 9568 37280 9580
rect 29144 9540 29180 9568
rect 37235 9540 37280 9568
rect 29086 9528 29092 9531
rect 29144 9528 29150 9540
rect 37274 9528 37280 9540
rect 37332 9528 37338 9580
rect 37366 9528 37372 9580
rect 37424 9568 37430 9580
rect 37533 9571 37591 9577
rect 37533 9568 37545 9571
rect 37424 9540 37545 9568
rect 37424 9528 37430 9540
rect 37533 9537 37545 9540
rect 37579 9537 37591 9571
rect 40494 9568 40500 9580
rect 40407 9540 40500 9568
rect 37533 9531 37591 9537
rect 40494 9528 40500 9540
rect 40552 9528 40558 9580
rect 40764 9571 40822 9577
rect 40764 9537 40776 9571
rect 40810 9568 40822 9571
rect 42058 9568 42064 9580
rect 40810 9540 42064 9568
rect 40810 9537 40822 9540
rect 40764 9531 40822 9537
rect 42058 9528 42064 9540
rect 42116 9528 42122 9580
rect 42444 9577 42472 9608
rect 42429 9571 42487 9577
rect 42429 9537 42441 9571
rect 42475 9537 42487 9571
rect 42429 9531 42487 9537
rect 42696 9571 42754 9577
rect 42696 9537 42708 9571
rect 42742 9568 42754 9571
rect 43898 9568 43904 9580
rect 42742 9540 43904 9568
rect 42742 9537 42754 9540
rect 42696 9531 42754 9537
rect 43898 9528 43904 9540
rect 43956 9528 43962 9580
rect 44284 9577 44312 9608
rect 49228 9605 49240 9639
rect 49274 9636 49286 9639
rect 51166 9636 51172 9648
rect 49274 9608 51172 9636
rect 49274 9605 49286 9608
rect 49228 9599 49286 9605
rect 51166 9596 51172 9608
rect 51224 9596 51230 9648
rect 53650 9645 53656 9648
rect 53644 9636 53656 9645
rect 53611 9608 53656 9636
rect 53644 9599 53656 9608
rect 53650 9596 53656 9599
rect 53708 9596 53714 9648
rect 56220 9639 56278 9645
rect 56220 9605 56232 9639
rect 56266 9636 56278 9639
rect 58250 9636 58256 9648
rect 56266 9608 58256 9636
rect 56266 9605 56278 9608
rect 56220 9599 56278 9605
rect 58250 9596 58256 9608
rect 58308 9596 58314 9648
rect 44269 9571 44327 9577
rect 44269 9537 44281 9571
rect 44315 9537 44327 9571
rect 44269 9531 44327 9537
rect 44536 9571 44594 9577
rect 44536 9537 44548 9571
rect 44582 9568 44594 9571
rect 45646 9568 45652 9580
rect 44582 9540 45652 9568
rect 44582 9537 44594 9540
rect 44536 9531 44594 9537
rect 45646 9528 45652 9540
rect 45704 9528 45710 9580
rect 48958 9568 48964 9580
rect 48919 9540 48964 9568
rect 48958 9528 48964 9540
rect 49016 9568 49022 9580
rect 50801 9571 50859 9577
rect 50801 9568 50813 9571
rect 49016 9540 50813 9568
rect 49016 9528 49022 9540
rect 50801 9537 50813 9540
rect 50847 9537 50859 9571
rect 50801 9531 50859 9537
rect 51068 9571 51126 9577
rect 51068 9537 51080 9571
rect 51114 9568 51126 9571
rect 52546 9568 52552 9580
rect 51114 9540 52552 9568
rect 51114 9537 51126 9540
rect 51068 9531 51126 9537
rect 5902 9460 5908 9512
rect 5960 9500 5966 9512
rect 6365 9503 6423 9509
rect 6365 9500 6377 9503
rect 5960 9472 6377 9500
rect 5960 9460 5966 9472
rect 6365 9469 6377 9472
rect 6411 9469 6423 9503
rect 9030 9500 9036 9512
rect 8991 9472 9036 9500
rect 6365 9463 6423 9469
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 19334 9500 19340 9512
rect 19295 9472 19340 9500
rect 19334 9460 19340 9472
rect 19392 9460 19398 9512
rect 28813 9503 28871 9509
rect 28813 9469 28825 9503
rect 28859 9469 28871 9503
rect 28813 9463 28871 9469
rect 18049 9435 18107 9441
rect 18049 9401 18061 9435
rect 18095 9432 18107 9435
rect 18230 9432 18236 9444
rect 18095 9404 18236 9432
rect 18095 9401 18107 9404
rect 18049 9395 18107 9401
rect 18230 9392 18236 9404
rect 18288 9392 18294 9444
rect 7742 9364 7748 9376
rect 7703 9336 7748 9364
rect 7742 9324 7748 9336
rect 7800 9324 7806 9376
rect 9214 9324 9220 9376
rect 9272 9364 9278 9376
rect 10413 9367 10471 9373
rect 10413 9364 10425 9367
rect 9272 9336 10425 9364
rect 9272 9324 9278 9336
rect 10413 9333 10425 9336
rect 10459 9333 10471 9367
rect 10413 9327 10471 9333
rect 14090 9324 14096 9376
rect 14148 9364 14154 9376
rect 14185 9367 14243 9373
rect 14185 9364 14197 9367
rect 14148 9336 14197 9364
rect 14148 9324 14154 9336
rect 14185 9333 14197 9336
rect 14231 9333 14243 9367
rect 24578 9364 24584 9376
rect 24539 9336 24584 9364
rect 14185 9327 14243 9333
rect 24578 9324 24584 9336
rect 24636 9324 24642 9376
rect 26421 9367 26479 9373
rect 26421 9333 26433 9367
rect 26467 9364 26479 9367
rect 26510 9364 26516 9376
rect 26467 9336 26516 9364
rect 26467 9333 26479 9336
rect 26421 9327 26479 9333
rect 26510 9324 26516 9336
rect 26568 9324 26574 9376
rect 28350 9364 28356 9376
rect 28311 9336 28356 9364
rect 28350 9324 28356 9336
rect 28408 9324 28414 9376
rect 28828 9364 28856 9463
rect 33410 9460 33416 9512
rect 33468 9500 33474 9512
rect 33781 9503 33839 9509
rect 33781 9500 33793 9503
rect 33468 9472 33793 9500
rect 33468 9460 33474 9472
rect 33781 9469 33793 9472
rect 33827 9469 33839 9503
rect 33781 9463 33839 9469
rect 28994 9364 29000 9376
rect 28828 9336 29000 9364
rect 28994 9324 29000 9336
rect 29052 9324 29058 9376
rect 34054 9324 34060 9376
rect 34112 9364 34118 9376
rect 35161 9367 35219 9373
rect 35161 9364 35173 9367
rect 34112 9336 35173 9364
rect 34112 9324 34118 9336
rect 35161 9333 35173 9336
rect 35207 9333 35219 9367
rect 43806 9364 43812 9376
rect 43767 9336 43812 9364
rect 35161 9327 35219 9333
rect 43806 9324 43812 9336
rect 43864 9324 43870 9376
rect 50816 9364 50844 9531
rect 52546 9528 52552 9540
rect 52604 9528 52610 9580
rect 53006 9460 53012 9512
rect 53064 9500 53070 9512
rect 53377 9503 53435 9509
rect 53377 9500 53389 9503
rect 53064 9472 53389 9500
rect 53064 9460 53070 9472
rect 53377 9469 53389 9472
rect 53423 9469 53435 9503
rect 53377 9463 53435 9469
rect 55306 9460 55312 9512
rect 55364 9500 55370 9512
rect 55953 9503 56011 9509
rect 55953 9500 55965 9503
rect 55364 9472 55965 9500
rect 55364 9460 55370 9472
rect 55953 9469 55965 9472
rect 55999 9469 56011 9503
rect 55953 9463 56011 9469
rect 52086 9392 52092 9444
rect 52144 9432 52150 9444
rect 52181 9435 52239 9441
rect 52181 9432 52193 9435
rect 52144 9404 52193 9432
rect 52144 9392 52150 9404
rect 52181 9401 52193 9404
rect 52227 9401 52239 9435
rect 57330 9432 57336 9444
rect 57291 9404 57336 9432
rect 52181 9395 52239 9401
rect 57330 9392 57336 9404
rect 57388 9392 57394 9444
rect 51166 9364 51172 9376
rect 50816 9336 51172 9364
rect 51166 9324 51172 9336
rect 51224 9364 51230 9376
rect 51534 9364 51540 9376
rect 51224 9336 51540 9364
rect 51224 9324 51230 9336
rect 51534 9324 51540 9336
rect 51592 9324 51598 9376
rect 53742 9324 53748 9376
rect 53800 9364 53806 9376
rect 54757 9367 54815 9373
rect 54757 9364 54769 9367
rect 53800 9336 54769 9364
rect 53800 9324 53806 9336
rect 54757 9333 54769 9336
rect 54803 9333 54815 9367
rect 54757 9327 54815 9333
rect 1104 9274 59340 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 59340 9274
rect 1104 9200 59340 9222
rect 7282 9160 7288 9172
rect 7243 9132 7288 9160
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 10321 9163 10379 9169
rect 10321 9129 10333 9163
rect 10367 9160 10379 9163
rect 11054 9160 11060 9172
rect 10367 9132 11060 9160
rect 10367 9129 10379 9132
rect 10321 9123 10379 9129
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 15470 9160 15476 9172
rect 15431 9132 15476 9160
rect 15470 9120 15476 9132
rect 15528 9120 15534 9172
rect 25774 9160 25780 9172
rect 25735 9132 25780 9160
rect 25774 9120 25780 9132
rect 25832 9120 25838 9172
rect 27614 9160 27620 9172
rect 27575 9132 27620 9160
rect 27614 9120 27620 9132
rect 27672 9120 27678 9172
rect 42058 9160 42064 9172
rect 42019 9132 42064 9160
rect 42058 9120 42064 9132
rect 42116 9120 42122 9172
rect 43898 9160 43904 9172
rect 43859 9132 43904 9160
rect 43898 9120 43904 9132
rect 43956 9120 43962 9172
rect 52546 9160 52552 9172
rect 52507 9132 52552 9160
rect 52546 9120 52552 9132
rect 52604 9120 52610 9172
rect 5350 8984 5356 9036
rect 5408 9024 5414 9036
rect 5902 9024 5908 9036
rect 5408 8996 5908 9024
rect 5408 8984 5414 8996
rect 5902 8984 5908 8996
rect 5960 8984 5966 9036
rect 19334 8984 19340 9036
rect 19392 9024 19398 9036
rect 20349 9027 20407 9033
rect 20349 9024 20361 9027
rect 19392 8996 20361 9024
rect 19392 8984 19398 8996
rect 20349 8993 20361 8996
rect 20395 8993 20407 9027
rect 20349 8987 20407 8993
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8956 4123 8959
rect 5368 8956 5396 8984
rect 4111 8928 5396 8956
rect 6172 8959 6230 8965
rect 4111 8925 4123 8928
rect 4065 8919 4123 8925
rect 6172 8925 6184 8959
rect 6218 8956 6230 8959
rect 7742 8956 7748 8968
rect 6218 8928 7748 8956
rect 6218 8925 6230 8928
rect 6172 8919 6230 8925
rect 7742 8916 7748 8928
rect 7800 8916 7806 8968
rect 8662 8916 8668 8968
rect 8720 8956 8726 8968
rect 9214 8965 9220 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8720 8928 8953 8956
rect 8720 8916 8726 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 9208 8956 9220 8965
rect 9175 8928 9220 8956
rect 8941 8919 8999 8925
rect 9208 8919 9220 8928
rect 9214 8916 9220 8919
rect 9272 8916 9278 8968
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8956 10839 8959
rect 10870 8956 10876 8968
rect 10827 8928 10876 8956
rect 10827 8925 10839 8928
rect 10781 8919 10839 8925
rect 10870 8916 10876 8928
rect 10928 8916 10934 8968
rect 14090 8956 14096 8968
rect 14051 8928 14096 8956
rect 14090 8916 14096 8928
rect 14148 8916 14154 8968
rect 14366 8965 14372 8968
rect 14360 8956 14372 8965
rect 14327 8928 14372 8956
rect 14360 8919 14372 8928
rect 14366 8916 14372 8919
rect 14424 8916 14430 8968
rect 20364 8956 20392 8987
rect 26234 8984 26240 9036
rect 26292 9024 26298 9036
rect 26292 8996 26337 9024
rect 26292 8984 26298 8996
rect 40494 8984 40500 9036
rect 40552 9024 40558 9036
rect 40681 9027 40739 9033
rect 40681 9024 40693 9027
rect 40552 8996 40693 9024
rect 40552 8984 40558 8996
rect 40681 8993 40693 8996
rect 40727 8993 40739 9027
rect 51166 9024 51172 9036
rect 51127 8996 51172 9024
rect 40681 8987 40739 8993
rect 22189 8959 22247 8965
rect 22189 8956 22201 8959
rect 20364 8928 22201 8956
rect 22189 8925 22201 8928
rect 22235 8925 22247 8959
rect 22189 8919 22247 8925
rect 23842 8916 23848 8968
rect 23900 8956 23906 8968
rect 24394 8956 24400 8968
rect 23900 8928 24400 8956
rect 23900 8916 23906 8928
rect 24394 8916 24400 8928
rect 24452 8916 24458 8968
rect 24664 8959 24722 8965
rect 24664 8925 24676 8959
rect 24710 8956 24722 8959
rect 25130 8956 25136 8968
rect 24710 8928 25136 8956
rect 24710 8925 24722 8928
rect 24664 8919 24722 8925
rect 25130 8916 25136 8928
rect 25188 8916 25194 8968
rect 26510 8965 26516 8968
rect 26504 8956 26516 8965
rect 26471 8928 26516 8956
rect 26504 8919 26516 8928
rect 26510 8916 26516 8919
rect 26568 8916 26574 8968
rect 29549 8959 29607 8965
rect 29549 8925 29561 8959
rect 29595 8956 29607 8959
rect 29638 8956 29644 8968
rect 29595 8928 29644 8956
rect 29595 8925 29607 8928
rect 29549 8919 29607 8925
rect 29638 8916 29644 8928
rect 29696 8916 29702 8968
rect 32306 8916 32312 8968
rect 32364 8956 32370 8968
rect 32401 8959 32459 8965
rect 32401 8956 32413 8959
rect 32364 8928 32413 8956
rect 32364 8916 32370 8928
rect 32401 8925 32413 8928
rect 32447 8925 32459 8959
rect 34422 8956 34428 8968
rect 32401 8919 32459 8925
rect 33704 8928 34428 8956
rect 4332 8891 4390 8897
rect 4332 8857 4344 8891
rect 4378 8888 4390 8891
rect 5626 8888 5632 8900
rect 4378 8860 5632 8888
rect 4378 8857 4390 8860
rect 4332 8851 4390 8857
rect 5626 8848 5632 8860
rect 5684 8848 5690 8900
rect 10410 8848 10416 8900
rect 10468 8888 10474 8900
rect 11026 8891 11084 8897
rect 11026 8888 11038 8891
rect 10468 8860 11038 8888
rect 10468 8848 10474 8860
rect 11026 8857 11038 8860
rect 11072 8857 11084 8891
rect 11026 8851 11084 8857
rect 20616 8891 20674 8897
rect 20616 8857 20628 8891
rect 20662 8888 20674 8891
rect 22002 8888 22008 8900
rect 20662 8860 22008 8888
rect 20662 8857 20674 8860
rect 20616 8851 20674 8857
rect 22002 8848 22008 8860
rect 22060 8848 22066 8900
rect 22456 8891 22514 8897
rect 22456 8857 22468 8891
rect 22502 8888 22514 8891
rect 23382 8888 23388 8900
rect 22502 8860 23388 8888
rect 22502 8857 22514 8860
rect 22456 8851 22514 8857
rect 23382 8848 23388 8860
rect 23440 8848 23446 8900
rect 29816 8891 29874 8897
rect 29816 8857 29828 8891
rect 29862 8888 29874 8891
rect 30466 8888 30472 8900
rect 29862 8860 30472 8888
rect 29862 8857 29874 8860
rect 29816 8851 29874 8857
rect 30466 8848 30472 8860
rect 30524 8848 30530 8900
rect 5442 8820 5448 8832
rect 5403 8792 5448 8820
rect 5442 8780 5448 8792
rect 5500 8780 5506 8832
rect 12158 8820 12164 8832
rect 12119 8792 12164 8820
rect 12158 8780 12164 8792
rect 12216 8780 12222 8832
rect 21726 8820 21732 8832
rect 21687 8792 21732 8820
rect 21726 8780 21732 8792
rect 21784 8780 21790 8832
rect 22186 8780 22192 8832
rect 22244 8820 22250 8832
rect 23569 8823 23627 8829
rect 23569 8820 23581 8823
rect 22244 8792 23581 8820
rect 22244 8780 22250 8792
rect 23569 8789 23581 8792
rect 23615 8789 23627 8823
rect 30926 8820 30932 8832
rect 30887 8792 30932 8820
rect 23569 8783 23627 8789
rect 30926 8780 30932 8792
rect 30984 8780 30990 8832
rect 33410 8780 33416 8832
rect 33468 8820 33474 8832
rect 33704 8829 33732 8928
rect 34422 8916 34428 8928
rect 34480 8956 34486 8968
rect 34701 8959 34759 8965
rect 34701 8956 34713 8959
rect 34480 8928 34713 8956
rect 34480 8916 34486 8928
rect 34701 8925 34713 8928
rect 34747 8925 34759 8959
rect 34701 8919 34759 8925
rect 35802 8916 35808 8968
rect 35860 8956 35866 8968
rect 36541 8959 36599 8965
rect 36541 8956 36553 8959
rect 35860 8928 36553 8956
rect 35860 8916 35866 8928
rect 36541 8925 36553 8928
rect 36587 8925 36599 8959
rect 40696 8956 40724 8987
rect 51166 8984 51172 8996
rect 51224 8984 51230 9036
rect 42521 8959 42579 8965
rect 42521 8956 42533 8959
rect 40696 8928 42533 8956
rect 36541 8919 36599 8925
rect 42521 8925 42533 8928
rect 42567 8925 42579 8959
rect 42521 8919 42579 8925
rect 45005 8959 45063 8965
rect 45005 8925 45017 8959
rect 45051 8956 45063 8959
rect 45738 8956 45744 8968
rect 45051 8928 45744 8956
rect 45051 8925 45063 8928
rect 45005 8919 45063 8925
rect 45738 8916 45744 8928
rect 45796 8956 45802 8968
rect 46842 8956 46848 8968
rect 45796 8928 46848 8956
rect 45796 8916 45802 8928
rect 46842 8916 46848 8928
rect 46900 8916 46906 8968
rect 34790 8848 34796 8900
rect 34848 8888 34854 8900
rect 34946 8891 35004 8897
rect 34946 8888 34958 8891
rect 34848 8860 34958 8888
rect 34848 8848 34854 8860
rect 34946 8857 34958 8860
rect 34992 8857 35004 8891
rect 34946 8851 35004 8857
rect 36630 8848 36636 8900
rect 36688 8888 36694 8900
rect 36786 8891 36844 8897
rect 36786 8888 36798 8891
rect 36688 8860 36798 8888
rect 36688 8848 36694 8860
rect 36786 8857 36798 8860
rect 36832 8857 36844 8891
rect 36786 8851 36844 8857
rect 40948 8891 41006 8897
rect 40948 8857 40960 8891
rect 40994 8888 41006 8891
rect 41874 8888 41880 8900
rect 40994 8860 41880 8888
rect 40994 8857 41006 8860
rect 40948 8851 41006 8857
rect 41874 8848 41880 8860
rect 41932 8848 41938 8900
rect 41966 8848 41972 8900
rect 42024 8888 42030 8900
rect 42766 8891 42824 8897
rect 42766 8888 42778 8891
rect 42024 8860 42778 8888
rect 42024 8848 42030 8860
rect 42766 8857 42778 8860
rect 42812 8857 42824 8891
rect 42766 8851 42824 8857
rect 44174 8848 44180 8900
rect 44232 8888 44238 8900
rect 47118 8897 47124 8900
rect 45250 8891 45308 8897
rect 45250 8888 45262 8891
rect 44232 8860 45262 8888
rect 44232 8848 44238 8860
rect 45250 8857 45262 8860
rect 45296 8857 45308 8891
rect 45250 8851 45308 8857
rect 47112 8851 47124 8897
rect 47176 8888 47182 8900
rect 51184 8888 51212 8984
rect 51436 8959 51494 8965
rect 51436 8925 51448 8959
rect 51482 8956 51494 8959
rect 52178 8956 52184 8968
rect 51482 8928 52184 8956
rect 51482 8925 51494 8928
rect 51436 8919 51494 8925
rect 52178 8916 52184 8928
rect 52236 8916 52242 8968
rect 53006 8956 53012 8968
rect 52919 8928 53012 8956
rect 53006 8916 53012 8928
rect 53064 8916 53070 8968
rect 55306 8956 55312 8968
rect 55267 8928 55312 8956
rect 55306 8916 55312 8928
rect 55364 8956 55370 8968
rect 57149 8959 57207 8965
rect 57149 8956 57161 8959
rect 55364 8928 57161 8956
rect 55364 8916 55370 8928
rect 57149 8925 57161 8928
rect 57195 8925 57207 8959
rect 57149 8919 57207 8925
rect 52638 8888 52644 8900
rect 47176 8860 47212 8888
rect 51184 8860 52644 8888
rect 47118 8848 47124 8851
rect 47176 8848 47182 8860
rect 52638 8848 52644 8860
rect 52696 8888 52702 8900
rect 53024 8888 53052 8916
rect 52696 8860 53052 8888
rect 53276 8891 53334 8897
rect 52696 8848 52702 8860
rect 53276 8857 53288 8891
rect 53322 8888 53334 8891
rect 54110 8888 54116 8900
rect 53322 8860 54116 8888
rect 53322 8857 53334 8860
rect 53276 8851 53334 8857
rect 54110 8848 54116 8860
rect 54168 8848 54174 8900
rect 55576 8891 55634 8897
rect 55576 8857 55588 8891
rect 55622 8888 55634 8891
rect 56594 8888 56600 8900
rect 55622 8860 56600 8888
rect 55622 8857 55634 8860
rect 55576 8851 55634 8857
rect 56594 8848 56600 8860
rect 56652 8848 56658 8900
rect 57416 8891 57474 8897
rect 57416 8857 57428 8891
rect 57462 8888 57474 8891
rect 58434 8888 58440 8900
rect 57462 8860 58440 8888
rect 57462 8857 57474 8860
rect 57416 8851 57474 8857
rect 58434 8848 58440 8860
rect 58492 8848 58498 8900
rect 33689 8823 33747 8829
rect 33689 8820 33701 8823
rect 33468 8792 33701 8820
rect 33468 8780 33474 8792
rect 33689 8789 33701 8792
rect 33735 8789 33747 8823
rect 36078 8820 36084 8832
rect 36039 8792 36084 8820
rect 33689 8783 33747 8789
rect 36078 8780 36084 8792
rect 36136 8780 36142 8832
rect 37918 8820 37924 8832
rect 37879 8792 37924 8820
rect 37918 8780 37924 8792
rect 37976 8780 37982 8832
rect 46382 8820 46388 8832
rect 46343 8792 46388 8820
rect 46382 8780 46388 8792
rect 46440 8780 46446 8832
rect 47394 8780 47400 8832
rect 47452 8820 47458 8832
rect 48225 8823 48283 8829
rect 48225 8820 48237 8823
rect 47452 8792 48237 8820
rect 47452 8780 47458 8792
rect 48225 8789 48237 8792
rect 48271 8789 48283 8823
rect 54386 8820 54392 8832
rect 54347 8792 54392 8820
rect 48225 8783 48283 8789
rect 54386 8780 54392 8792
rect 54444 8780 54450 8832
rect 55858 8780 55864 8832
rect 55916 8820 55922 8832
rect 56689 8823 56747 8829
rect 56689 8820 56701 8823
rect 55916 8792 56701 8820
rect 55916 8780 55922 8792
rect 56689 8789 56701 8792
rect 56735 8789 56747 8823
rect 58526 8820 58532 8832
rect 58487 8792 58532 8820
rect 56689 8783 56747 8789
rect 58526 8780 58532 8792
rect 58584 8780 58590 8832
rect 1104 8730 59340 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 59340 8730
rect 1104 8656 59340 8678
rect 10410 8616 10416 8628
rect 10371 8588 10416 8616
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 12802 8576 12808 8628
rect 12860 8616 12866 8628
rect 13633 8619 13691 8625
rect 13633 8616 13645 8619
rect 12860 8588 13645 8616
rect 12860 8576 12866 8588
rect 13633 8585 13645 8588
rect 13679 8585 13691 8619
rect 19334 8616 19340 8628
rect 13633 8579 13691 8585
rect 19168 8588 19340 8616
rect 4700 8551 4758 8557
rect 4700 8517 4712 8551
rect 4746 8548 4758 8551
rect 5442 8548 5448 8560
rect 4746 8520 5448 8548
rect 4746 8517 4758 8520
rect 4700 8511 4758 8517
rect 5442 8508 5448 8520
rect 5500 8508 5506 8560
rect 6632 8551 6690 8557
rect 6632 8517 6644 8551
rect 6678 8548 6690 8551
rect 7466 8548 7472 8560
rect 6678 8520 7472 8548
rect 6678 8517 6690 8520
rect 6632 8511 6690 8517
rect 7466 8508 7472 8520
rect 7524 8508 7530 8560
rect 9300 8551 9358 8557
rect 9300 8517 9312 8551
rect 9346 8548 9358 8551
rect 10594 8548 10600 8560
rect 9346 8520 10600 8548
rect 9346 8517 9358 8520
rect 9300 8511 9358 8517
rect 10594 8508 10600 8520
rect 10652 8508 10658 8560
rect 12158 8508 12164 8560
rect 12216 8548 12222 8560
rect 12498 8551 12556 8557
rect 12498 8548 12510 8551
rect 12216 8520 12510 8548
rect 12216 8508 12222 8520
rect 12498 8517 12510 8520
rect 12544 8517 12556 8551
rect 12498 8511 12556 8517
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8480 4491 8483
rect 5258 8480 5264 8492
rect 4479 8452 5264 8480
rect 4479 8449 4491 8452
rect 4433 8443 4491 8449
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 14544 8483 14602 8489
rect 14544 8449 14556 8483
rect 14590 8480 14602 8483
rect 16022 8480 16028 8492
rect 14590 8452 16028 8480
rect 14590 8449 14602 8452
rect 14544 8443 14602 8449
rect 16022 8440 16028 8452
rect 16080 8440 16086 8492
rect 5902 8372 5908 8424
rect 5960 8412 5966 8424
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 5960 8384 6377 8412
rect 5960 8372 5966 8384
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 6365 8375 6423 8381
rect 8662 8372 8668 8424
rect 8720 8412 8726 8424
rect 9033 8415 9091 8421
rect 9033 8412 9045 8415
rect 8720 8384 9045 8412
rect 8720 8372 8726 8384
rect 9033 8381 9045 8384
rect 9079 8381 9091 8415
rect 9033 8375 9091 8381
rect 12158 8372 12164 8424
rect 12216 8412 12222 8424
rect 12253 8415 12311 8421
rect 12253 8412 12265 8415
rect 12216 8384 12265 8412
rect 12216 8372 12222 8384
rect 12253 8381 12265 8384
rect 12299 8381 12311 8415
rect 12253 8375 12311 8381
rect 14090 8372 14096 8424
rect 14148 8412 14154 8424
rect 14277 8415 14335 8421
rect 14277 8412 14289 8415
rect 14148 8384 14289 8412
rect 14148 8372 14154 8384
rect 14277 8381 14289 8384
rect 14323 8381 14335 8415
rect 14277 8375 14335 8381
rect 17310 8372 17316 8424
rect 17368 8412 17374 8424
rect 19168 8421 19196 8588
rect 19334 8576 19340 8588
rect 19392 8576 19398 8628
rect 20530 8616 20536 8628
rect 20491 8588 20536 8616
rect 20530 8576 20536 8588
rect 20588 8576 20594 8628
rect 23382 8616 23388 8628
rect 23343 8588 23388 8616
rect 23382 8576 23388 8588
rect 23440 8576 23446 8628
rect 24946 8576 24952 8628
rect 25004 8616 25010 8628
rect 25225 8619 25283 8625
rect 25225 8616 25237 8619
rect 25004 8588 25237 8616
rect 25004 8576 25010 8588
rect 25225 8585 25237 8588
rect 25271 8585 25283 8619
rect 25225 8579 25283 8585
rect 28353 8619 28411 8625
rect 28353 8585 28365 8619
rect 28399 8585 28411 8619
rect 28353 8579 28411 8585
rect 19420 8551 19478 8557
rect 19420 8517 19432 8551
rect 19466 8548 19478 8551
rect 21726 8548 21732 8560
rect 19466 8520 21732 8548
rect 19466 8517 19478 8520
rect 19420 8511 19478 8517
rect 21726 8508 21732 8520
rect 21784 8508 21790 8560
rect 22272 8551 22330 8557
rect 22272 8517 22284 8551
rect 22318 8548 22330 8551
rect 24578 8548 24584 8560
rect 22318 8520 24584 8548
rect 22318 8517 22330 8520
rect 22272 8511 22330 8517
rect 24578 8508 24584 8520
rect 24636 8508 24642 8560
rect 28368 8548 28396 8579
rect 28534 8576 28540 8628
rect 28592 8616 28598 8628
rect 30193 8619 30251 8625
rect 30193 8616 30205 8619
rect 28592 8588 30205 8616
rect 28592 8576 28598 8588
rect 30193 8585 30205 8588
rect 30239 8585 30251 8619
rect 34790 8616 34796 8628
rect 34751 8588 34796 8616
rect 30193 8579 30251 8585
rect 34790 8576 34796 8588
rect 34848 8576 34854 8628
rect 36630 8616 36636 8628
rect 36591 8588 36636 8616
rect 36630 8576 36636 8588
rect 36688 8576 36694 8628
rect 45646 8616 45652 8628
rect 45607 8588 45652 8616
rect 45646 8576 45652 8588
rect 45704 8576 45710 8628
rect 48961 8619 49019 8625
rect 48961 8585 48973 8619
rect 49007 8585 49019 8619
rect 54110 8616 54116 8628
rect 54071 8588 54116 8616
rect 48961 8579 49019 8585
rect 29058 8551 29116 8557
rect 29058 8548 29070 8551
rect 28368 8520 29070 8548
rect 29058 8517 29070 8520
rect 29104 8517 29116 8551
rect 29058 8511 29116 8517
rect 33680 8551 33738 8557
rect 33680 8517 33692 8551
rect 33726 8548 33738 8551
rect 34146 8548 34152 8560
rect 33726 8520 34152 8548
rect 33726 8517 33738 8520
rect 33680 8511 33738 8517
rect 34146 8508 34152 8520
rect 34204 8508 34210 8560
rect 37544 8551 37602 8557
rect 37544 8517 37556 8551
rect 37590 8548 37602 8551
rect 37918 8548 37924 8560
rect 37590 8520 37924 8548
rect 37590 8517 37602 8520
rect 37544 8511 37602 8517
rect 37918 8508 37924 8520
rect 37976 8508 37982 8560
rect 44536 8551 44594 8557
rect 44536 8517 44548 8551
rect 44582 8548 44594 8551
rect 46382 8548 46388 8560
rect 44582 8520 46388 8548
rect 44582 8517 44594 8520
rect 44536 8511 44594 8517
rect 46382 8508 46388 8520
rect 46440 8508 46446 8560
rect 48976 8548 49004 8579
rect 54110 8576 54116 8588
rect 54168 8576 54174 8628
rect 49666 8551 49724 8557
rect 49666 8548 49678 8551
rect 48976 8520 49678 8548
rect 49666 8517 49678 8520
rect 49712 8517 49724 8551
rect 49666 8511 49724 8517
rect 53834 8508 53840 8560
rect 53892 8548 53898 8560
rect 54849 8551 54907 8557
rect 54849 8548 54861 8551
rect 53892 8520 54861 8548
rect 53892 8508 53898 8520
rect 54849 8517 54861 8520
rect 54895 8517 54907 8551
rect 54849 8511 54907 8517
rect 24112 8483 24170 8489
rect 24112 8449 24124 8483
rect 24158 8480 24170 8483
rect 25774 8480 25780 8492
rect 24158 8452 25780 8480
rect 24158 8449 24170 8452
rect 24112 8443 24170 8449
rect 25774 8440 25780 8452
rect 25832 8440 25838 8492
rect 26234 8440 26240 8492
rect 26292 8480 26298 8492
rect 26973 8483 27031 8489
rect 26973 8480 26985 8483
rect 26292 8452 26985 8480
rect 26292 8440 26298 8452
rect 26973 8449 26985 8452
rect 27019 8449 27031 8483
rect 26973 8443 27031 8449
rect 27240 8483 27298 8489
rect 27240 8449 27252 8483
rect 27286 8480 27298 8483
rect 27614 8480 27620 8492
rect 27286 8452 27620 8480
rect 27286 8449 27298 8452
rect 27240 8443 27298 8449
rect 27614 8440 27620 8452
rect 27672 8440 27678 8492
rect 34422 8440 34428 8492
rect 34480 8480 34486 8492
rect 35253 8483 35311 8489
rect 35253 8480 35265 8483
rect 34480 8452 35265 8480
rect 34480 8440 34486 8452
rect 35253 8449 35265 8452
rect 35299 8449 35311 8483
rect 35253 8443 35311 8449
rect 35520 8483 35578 8489
rect 35520 8449 35532 8483
rect 35566 8480 35578 8483
rect 35986 8480 35992 8492
rect 35566 8452 35992 8480
rect 35566 8449 35578 8452
rect 35520 8443 35578 8449
rect 35986 8440 35992 8452
rect 36044 8440 36050 8492
rect 37274 8480 37280 8492
rect 37235 8452 37280 8480
rect 37274 8440 37280 8452
rect 37332 8480 37338 8492
rect 37332 8452 38792 8480
rect 37332 8440 37338 8452
rect 19153 8415 19211 8421
rect 19153 8412 19165 8415
rect 17368 8384 19165 8412
rect 17368 8372 17374 8384
rect 19153 8381 19165 8384
rect 19199 8381 19211 8415
rect 19153 8375 19211 8381
rect 21634 8372 21640 8424
rect 21692 8412 21698 8424
rect 22005 8415 22063 8421
rect 22005 8412 22017 8415
rect 21692 8384 22017 8412
rect 21692 8372 21698 8384
rect 22005 8381 22017 8384
rect 22051 8381 22063 8415
rect 23842 8412 23848 8424
rect 23803 8384 23848 8412
rect 22005 8375 22063 8381
rect 23842 8372 23848 8384
rect 23900 8372 23906 8424
rect 28718 8372 28724 8424
rect 28776 8412 28782 8424
rect 28813 8415 28871 8421
rect 28813 8412 28825 8415
rect 28776 8384 28825 8412
rect 28776 8372 28782 8384
rect 28813 8381 28825 8384
rect 28859 8381 28871 8415
rect 33410 8412 33416 8424
rect 33371 8384 33416 8412
rect 28813 8375 28871 8381
rect 33410 8372 33416 8384
rect 33468 8372 33474 8424
rect 38764 8412 38792 8452
rect 38838 8440 38844 8492
rect 38896 8480 38902 8492
rect 39373 8483 39431 8489
rect 39373 8480 39385 8483
rect 38896 8452 39385 8480
rect 38896 8440 38902 8452
rect 39373 8449 39385 8452
rect 39419 8449 39431 8483
rect 39373 8443 39431 8449
rect 41414 8440 41420 8492
rect 41472 8480 41478 8492
rect 42685 8483 42743 8489
rect 42685 8480 42697 8483
rect 41472 8452 42697 8480
rect 41472 8440 41478 8452
rect 42685 8449 42697 8452
rect 42731 8449 42743 8483
rect 42685 8443 42743 8449
rect 44269 8483 44327 8489
rect 44269 8449 44281 8483
rect 44315 8480 44327 8483
rect 45738 8480 45744 8492
rect 44315 8452 45744 8480
rect 44315 8449 44327 8452
rect 44269 8443 44327 8449
rect 45738 8440 45744 8452
rect 45796 8440 45802 8492
rect 46842 8440 46848 8492
rect 46900 8480 46906 8492
rect 47581 8483 47639 8489
rect 47581 8480 47593 8483
rect 46900 8452 47593 8480
rect 46900 8440 46906 8452
rect 47581 8449 47593 8452
rect 47627 8449 47639 8483
rect 47581 8443 47639 8449
rect 47848 8483 47906 8489
rect 47848 8449 47860 8483
rect 47894 8480 47906 8483
rect 48222 8480 48228 8492
rect 47894 8452 48228 8480
rect 47894 8449 47906 8452
rect 47848 8443 47906 8449
rect 48222 8440 48228 8452
rect 48280 8440 48286 8492
rect 49421 8483 49479 8489
rect 49421 8449 49433 8483
rect 49467 8480 49479 8483
rect 50154 8480 50160 8492
rect 49467 8452 50160 8480
rect 49467 8449 49479 8452
rect 49421 8443 49479 8449
rect 50154 8440 50160 8452
rect 50212 8480 50218 8492
rect 52730 8480 52736 8492
rect 50212 8452 52736 8480
rect 50212 8440 50218 8452
rect 52730 8440 52736 8452
rect 52788 8440 52794 8492
rect 53000 8483 53058 8489
rect 53000 8449 53012 8483
rect 53046 8480 53058 8483
rect 54110 8480 54116 8492
rect 53046 8452 54116 8480
rect 53046 8449 53058 8452
rect 53000 8443 53058 8449
rect 54110 8440 54116 8452
rect 54168 8440 54174 8492
rect 39117 8415 39175 8421
rect 39117 8412 39129 8415
rect 38764 8384 39129 8412
rect 39117 8381 39129 8384
rect 39163 8381 39175 8415
rect 39117 8375 39175 8381
rect 40494 8372 40500 8424
rect 40552 8412 40558 8424
rect 42429 8415 42487 8421
rect 42429 8412 42441 8415
rect 40552 8384 42441 8412
rect 40552 8372 40558 8384
rect 42429 8381 42441 8384
rect 42475 8381 42487 8415
rect 42429 8375 42487 8381
rect 5442 8304 5448 8356
rect 5500 8344 5506 8356
rect 5813 8347 5871 8353
rect 5813 8344 5825 8347
rect 5500 8316 5825 8344
rect 5500 8304 5506 8316
rect 5813 8313 5825 8316
rect 5859 8313 5871 8347
rect 15657 8347 15715 8353
rect 15657 8344 15669 8347
rect 5813 8307 5871 8313
rect 15212 8316 15669 8344
rect 7742 8276 7748 8288
rect 7703 8248 7748 8276
rect 7742 8236 7748 8248
rect 7800 8236 7806 8288
rect 13814 8236 13820 8288
rect 13872 8276 13878 8288
rect 15212 8276 15240 8316
rect 15657 8313 15669 8316
rect 15703 8313 15715 8347
rect 15657 8307 15715 8313
rect 38654 8276 38660 8288
rect 13872 8248 15240 8276
rect 38615 8248 38660 8276
rect 13872 8236 13878 8248
rect 38654 8236 38660 8248
rect 38712 8236 38718 8288
rect 40494 8276 40500 8288
rect 40455 8248 40500 8276
rect 40494 8236 40500 8248
rect 40552 8236 40558 8288
rect 42444 8276 42472 8375
rect 43622 8304 43628 8356
rect 43680 8344 43686 8356
rect 43809 8347 43867 8353
rect 43809 8344 43821 8347
rect 43680 8316 43821 8344
rect 43680 8304 43686 8316
rect 43809 8313 43821 8316
rect 43855 8313 43867 8347
rect 43809 8307 43867 8313
rect 42794 8276 42800 8288
rect 42444 8248 42800 8276
rect 42794 8236 42800 8248
rect 42852 8236 42858 8288
rect 50798 8276 50804 8288
rect 50759 8248 50804 8276
rect 50798 8236 50804 8248
rect 50856 8236 50862 8288
rect 55306 8236 55312 8288
rect 55364 8276 55370 8288
rect 56137 8279 56195 8285
rect 56137 8276 56149 8279
rect 55364 8248 56149 8276
rect 55364 8236 55370 8248
rect 56137 8245 56149 8248
rect 56183 8245 56195 8279
rect 56137 8239 56195 8245
rect 1104 8186 59340 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 59340 8186
rect 1104 8112 59340 8134
rect 5626 8032 5632 8084
rect 5684 8072 5690 8084
rect 7285 8075 7343 8081
rect 7285 8072 7297 8075
rect 5684 8044 7297 8072
rect 5684 8032 5690 8044
rect 7285 8041 7297 8044
rect 7331 8041 7343 8075
rect 7285 8035 7343 8041
rect 11701 8075 11759 8081
rect 11701 8041 11713 8075
rect 11747 8072 11759 8075
rect 11790 8072 11796 8084
rect 11747 8044 11796 8072
rect 11747 8041 11759 8044
rect 11701 8035 11759 8041
rect 11790 8032 11796 8044
rect 11848 8032 11854 8084
rect 22002 8032 22008 8084
rect 22060 8072 22066 8084
rect 23017 8075 23075 8081
rect 23017 8072 23029 8075
rect 22060 8044 23029 8072
rect 22060 8032 22066 8044
rect 23017 8041 23029 8044
rect 23063 8041 23075 8075
rect 25774 8072 25780 8084
rect 25735 8044 25780 8072
rect 23017 8035 23075 8041
rect 25774 8032 25780 8044
rect 25832 8032 25838 8084
rect 27614 8072 27620 8084
rect 27575 8044 27620 8072
rect 27614 8032 27620 8044
rect 27672 8032 27678 8084
rect 30466 8032 30472 8084
rect 30524 8072 30530 8084
rect 30929 8075 30987 8081
rect 30929 8072 30941 8075
rect 30524 8044 30941 8072
rect 30524 8032 30530 8044
rect 30929 8041 30941 8044
rect 30975 8041 30987 8075
rect 30929 8035 30987 8041
rect 35986 8032 35992 8084
rect 36044 8072 36050 8084
rect 36081 8075 36139 8081
rect 36081 8072 36093 8075
rect 36044 8044 36093 8072
rect 36044 8032 36050 8044
rect 36081 8041 36093 8044
rect 36127 8041 36139 8075
rect 38838 8072 38844 8084
rect 38799 8044 38844 8072
rect 36081 8035 36139 8041
rect 38838 8032 38844 8044
rect 38896 8032 38902 8084
rect 42794 8032 42800 8084
rect 42852 8072 42858 8084
rect 43073 8075 43131 8081
rect 43073 8072 43085 8075
rect 42852 8044 43085 8072
rect 42852 8032 42858 8044
rect 43073 8041 43085 8044
rect 43119 8041 43131 8075
rect 43073 8035 43131 8041
rect 46385 8075 46443 8081
rect 46385 8041 46397 8075
rect 46431 8072 46443 8075
rect 47118 8072 47124 8084
rect 46431 8044 47124 8072
rect 46431 8041 46443 8044
rect 46385 8035 46443 8041
rect 47118 8032 47124 8044
rect 47176 8032 47182 8084
rect 48222 8072 48228 8084
rect 48183 8044 48228 8072
rect 48222 8032 48228 8044
rect 48280 8032 48286 8084
rect 54110 8072 54116 8084
rect 54071 8044 54116 8072
rect 54110 8032 54116 8044
rect 54168 8032 54174 8084
rect 56594 8032 56600 8084
rect 56652 8072 56658 8084
rect 56689 8075 56747 8081
rect 56689 8072 56701 8075
rect 56652 8044 56701 8072
rect 56652 8032 56658 8044
rect 56689 8041 56701 8044
rect 56735 8041 56747 8075
rect 56689 8035 56747 8041
rect 58434 8032 58440 8084
rect 58492 8072 58498 8084
rect 58529 8075 58587 8081
rect 58529 8072 58541 8075
rect 58492 8044 58541 8072
rect 58492 8032 58498 8044
rect 58529 8041 58541 8044
rect 58575 8041 58587 8075
rect 58529 8035 58587 8041
rect 26234 7896 26240 7948
rect 26292 7936 26298 7948
rect 46842 7936 46848 7948
rect 26292 7908 26337 7936
rect 46803 7908 46848 7936
rect 26292 7896 26298 7908
rect 46842 7896 46848 7908
rect 46900 7896 46906 7948
rect 50154 7936 50160 7948
rect 50115 7908 50160 7936
rect 50154 7896 50160 7908
rect 50212 7896 50218 7948
rect 52638 7896 52644 7948
rect 52696 7936 52702 7948
rect 52733 7939 52791 7945
rect 52733 7936 52745 7939
rect 52696 7908 52745 7936
rect 52696 7896 52702 7908
rect 52733 7905 52745 7908
rect 52779 7905 52791 7939
rect 52733 7899 52791 7905
rect 1854 7868 1860 7880
rect 1815 7840 1860 7868
rect 1854 7828 1860 7840
rect 1912 7828 1918 7880
rect 4065 7871 4123 7877
rect 4065 7837 4077 7871
rect 4111 7868 4123 7871
rect 4154 7868 4160 7880
rect 4111 7840 4160 7868
rect 4111 7837 4123 7840
rect 4065 7831 4123 7837
rect 4154 7828 4160 7840
rect 4212 7868 4218 7880
rect 5350 7868 5356 7880
rect 4212 7840 5356 7868
rect 4212 7828 4218 7840
rect 5350 7828 5356 7840
rect 5408 7828 5414 7880
rect 5902 7868 5908 7880
rect 5863 7840 5908 7868
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 6172 7871 6230 7877
rect 6172 7837 6184 7871
rect 6218 7868 6230 7871
rect 7742 7868 7748 7880
rect 6218 7840 7748 7868
rect 6218 7837 6230 7840
rect 6172 7831 6230 7837
rect 7742 7828 7748 7840
rect 7800 7828 7806 7880
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7868 10379 7871
rect 12158 7868 12164 7880
rect 10367 7840 12164 7868
rect 10367 7837 10379 7840
rect 10321 7831 10379 7837
rect 12158 7828 12164 7840
rect 12216 7828 12222 7880
rect 14461 7871 14519 7877
rect 14461 7837 14473 7871
rect 14507 7868 14519 7871
rect 16301 7871 16359 7877
rect 16301 7868 16313 7871
rect 14507 7840 16313 7868
rect 14507 7837 14519 7840
rect 14461 7831 14519 7837
rect 14844 7812 14872 7840
rect 16301 7837 16313 7840
rect 16347 7868 16359 7871
rect 16850 7868 16856 7880
rect 16347 7840 16856 7868
rect 16347 7837 16359 7840
rect 16301 7831 16359 7837
rect 16850 7828 16856 7840
rect 16908 7868 16914 7880
rect 17310 7868 17316 7880
rect 16908 7840 17316 7868
rect 16908 7828 16914 7840
rect 17310 7828 17316 7840
rect 17368 7828 17374 7880
rect 19337 7871 19395 7877
rect 19337 7837 19349 7871
rect 19383 7868 19395 7871
rect 21634 7868 21640 7880
rect 19383 7840 21640 7868
rect 19383 7837 19395 7840
rect 19337 7831 19395 7837
rect 21634 7828 21640 7840
rect 21692 7828 21698 7880
rect 21904 7871 21962 7877
rect 21904 7837 21916 7871
rect 21950 7868 21962 7871
rect 22186 7868 22192 7880
rect 21950 7840 22192 7868
rect 21950 7837 21962 7840
rect 21904 7831 21962 7837
rect 22186 7828 22192 7840
rect 22244 7828 22250 7880
rect 24302 7828 24308 7880
rect 24360 7868 24366 7880
rect 24397 7871 24455 7877
rect 24397 7868 24409 7871
rect 24360 7840 24409 7868
rect 24360 7828 24366 7840
rect 24397 7837 24409 7840
rect 24443 7837 24455 7871
rect 24397 7831 24455 7837
rect 2124 7803 2182 7809
rect 2124 7769 2136 7803
rect 2170 7800 2182 7803
rect 4332 7803 4390 7809
rect 2170 7772 3832 7800
rect 2170 7769 2182 7772
rect 2124 7763 2182 7769
rect 3234 7732 3240 7744
rect 3195 7704 3240 7732
rect 3234 7692 3240 7704
rect 3292 7692 3298 7744
rect 3804 7732 3832 7772
rect 4332 7769 4344 7803
rect 4378 7800 4390 7803
rect 6546 7800 6552 7812
rect 4378 7772 6552 7800
rect 4378 7769 4390 7772
rect 4332 7763 4390 7769
rect 6546 7760 6552 7772
rect 6604 7760 6610 7812
rect 10588 7803 10646 7809
rect 10588 7769 10600 7803
rect 10634 7800 10646 7803
rect 12250 7800 12256 7812
rect 10634 7772 12256 7800
rect 10634 7769 10646 7772
rect 10588 7763 10646 7769
rect 12250 7760 12256 7772
rect 12308 7760 12314 7812
rect 12428 7803 12486 7809
rect 12428 7769 12440 7803
rect 12474 7800 12486 7803
rect 13078 7800 13084 7812
rect 12474 7772 13084 7800
rect 12474 7769 12486 7772
rect 12428 7763 12486 7769
rect 13078 7760 13084 7772
rect 13136 7760 13142 7812
rect 14728 7803 14786 7809
rect 14728 7769 14740 7803
rect 14774 7769 14786 7803
rect 14728 7763 14786 7769
rect 5445 7735 5503 7741
rect 5445 7732 5457 7735
rect 3804 7704 5457 7732
rect 5445 7701 5457 7704
rect 5491 7701 5503 7735
rect 13538 7732 13544 7744
rect 13499 7704 13544 7732
rect 5445 7695 5503 7701
rect 13538 7692 13544 7704
rect 13596 7692 13602 7744
rect 14752 7732 14780 7763
rect 14826 7760 14832 7812
rect 14884 7760 14890 7812
rect 16206 7800 16212 7812
rect 15672 7772 16212 7800
rect 15672 7732 15700 7772
rect 16206 7760 16212 7772
rect 16264 7760 16270 7812
rect 16568 7803 16626 7809
rect 16568 7769 16580 7803
rect 16614 7800 16626 7803
rect 18322 7800 18328 7812
rect 16614 7772 18328 7800
rect 16614 7769 16626 7772
rect 16568 7763 16626 7769
rect 18322 7760 18328 7772
rect 18380 7760 18386 7812
rect 19604 7803 19662 7809
rect 19604 7769 19616 7803
rect 19650 7800 19662 7803
rect 21082 7800 21088 7812
rect 19650 7772 21088 7800
rect 19650 7769 19662 7772
rect 19604 7763 19662 7769
rect 21082 7760 21088 7772
rect 21140 7760 21146 7812
rect 21652 7800 21680 7828
rect 22002 7800 22008 7812
rect 21652 7772 22008 7800
rect 22002 7760 22008 7772
rect 22060 7760 22066 7812
rect 24664 7803 24722 7809
rect 24664 7769 24676 7803
rect 24710 7800 24722 7803
rect 25222 7800 25228 7812
rect 24710 7772 25228 7800
rect 24710 7769 24722 7772
rect 24664 7763 24722 7769
rect 25222 7760 25228 7772
rect 25280 7760 25286 7812
rect 26252 7800 26280 7896
rect 26504 7871 26562 7877
rect 26504 7837 26516 7871
rect 26550 7868 26562 7871
rect 28350 7868 28356 7880
rect 26550 7840 28356 7868
rect 26550 7837 26562 7840
rect 26504 7831 26562 7837
rect 28350 7828 28356 7840
rect 28408 7828 28414 7880
rect 29822 7877 29828 7880
rect 29549 7871 29607 7877
rect 29549 7837 29561 7871
rect 29595 7837 29607 7871
rect 29816 7868 29828 7877
rect 29783 7840 29828 7868
rect 29549 7831 29607 7837
rect 29816 7831 29828 7840
rect 26970 7800 26976 7812
rect 26252 7772 26976 7800
rect 26970 7760 26976 7772
rect 27028 7800 27034 7812
rect 29564 7800 29592 7831
rect 29822 7828 29828 7831
rect 29880 7828 29886 7880
rect 32122 7868 32128 7880
rect 32083 7840 32128 7868
rect 32122 7828 32128 7840
rect 32180 7828 32186 7880
rect 32214 7828 32220 7880
rect 32272 7868 32278 7880
rect 32381 7871 32439 7877
rect 32381 7868 32393 7871
rect 32272 7840 32393 7868
rect 32272 7828 32278 7840
rect 32381 7837 32393 7840
rect 32427 7837 32439 7871
rect 32381 7831 32439 7837
rect 34701 7871 34759 7877
rect 34701 7837 34713 7871
rect 34747 7837 34759 7871
rect 34701 7831 34759 7837
rect 34968 7871 35026 7877
rect 34968 7837 34980 7871
rect 35014 7868 35026 7871
rect 36078 7868 36084 7880
rect 35014 7840 36084 7868
rect 35014 7837 35026 7840
rect 34968 7831 35026 7837
rect 27028 7772 29592 7800
rect 32140 7800 32168 7828
rect 33410 7800 33416 7812
rect 32140 7772 33416 7800
rect 27028 7760 27034 7772
rect 33410 7760 33416 7772
rect 33468 7760 33474 7812
rect 34716 7800 34744 7831
rect 36078 7828 36084 7840
rect 36136 7828 36142 7880
rect 37461 7871 37519 7877
rect 37461 7837 37473 7871
rect 37507 7837 37519 7871
rect 37461 7831 37519 7837
rect 37728 7871 37786 7877
rect 37728 7837 37740 7871
rect 37774 7868 37786 7871
rect 38654 7868 38660 7880
rect 37774 7840 38660 7868
rect 37774 7837 37786 7840
rect 37728 7831 37786 7837
rect 35802 7800 35808 7812
rect 34716 7772 35808 7800
rect 35802 7760 35808 7772
rect 35860 7800 35866 7812
rect 37476 7800 37504 7831
rect 38654 7828 38660 7840
rect 38712 7828 38718 7880
rect 41690 7828 41696 7880
rect 41748 7868 41754 7880
rect 41785 7871 41843 7877
rect 41785 7868 41797 7871
rect 41748 7840 41797 7868
rect 41748 7828 41754 7840
rect 41785 7837 41797 7840
rect 41831 7837 41843 7871
rect 41785 7831 41843 7837
rect 45005 7871 45063 7877
rect 45005 7837 45017 7871
rect 45051 7868 45063 7871
rect 45738 7868 45744 7880
rect 45051 7840 45744 7868
rect 45051 7837 45063 7840
rect 45005 7831 45063 7837
rect 45738 7828 45744 7840
rect 45796 7828 45802 7880
rect 47112 7871 47170 7877
rect 47112 7837 47124 7871
rect 47158 7868 47170 7871
rect 47394 7868 47400 7880
rect 47158 7840 47400 7868
rect 47158 7837 47170 7840
rect 47112 7831 47170 7837
rect 47394 7828 47400 7840
rect 47452 7828 47458 7880
rect 55306 7868 55312 7880
rect 55267 7840 55312 7868
rect 55306 7828 55312 7840
rect 55364 7868 55370 7880
rect 57149 7871 57207 7877
rect 57149 7868 57161 7871
rect 55364 7840 57161 7868
rect 55364 7828 55370 7840
rect 57149 7837 57161 7840
rect 57195 7837 57207 7871
rect 57149 7831 57207 7837
rect 35860 7772 37504 7800
rect 45272 7803 45330 7809
rect 35860 7760 35866 7772
rect 45272 7769 45284 7803
rect 45318 7800 45330 7803
rect 45370 7800 45376 7812
rect 45318 7772 45376 7800
rect 45318 7769 45330 7772
rect 45272 7763 45330 7769
rect 45370 7760 45376 7772
rect 45428 7760 45434 7812
rect 50424 7803 50482 7809
rect 50424 7769 50436 7803
rect 50470 7800 50482 7803
rect 50614 7800 50620 7812
rect 50470 7772 50620 7800
rect 50470 7769 50482 7772
rect 50424 7763 50482 7769
rect 50614 7760 50620 7772
rect 50672 7760 50678 7812
rect 53000 7803 53058 7809
rect 53000 7769 53012 7803
rect 53046 7800 53058 7803
rect 54018 7800 54024 7812
rect 53046 7772 54024 7800
rect 53046 7769 53058 7772
rect 53000 7763 53058 7769
rect 54018 7760 54024 7772
rect 54076 7760 54082 7812
rect 55576 7803 55634 7809
rect 55576 7769 55588 7803
rect 55622 7800 55634 7803
rect 55950 7800 55956 7812
rect 55622 7772 55956 7800
rect 55622 7769 55634 7772
rect 55576 7763 55634 7769
rect 55950 7760 55956 7772
rect 56008 7760 56014 7812
rect 56778 7760 56784 7812
rect 56836 7800 56842 7812
rect 57394 7803 57452 7809
rect 57394 7800 57406 7803
rect 56836 7772 57406 7800
rect 56836 7760 56842 7772
rect 57394 7769 57406 7772
rect 57440 7769 57452 7803
rect 57394 7763 57452 7769
rect 15838 7732 15844 7744
rect 14752 7704 15700 7732
rect 15799 7704 15844 7732
rect 15838 7692 15844 7704
rect 15896 7692 15902 7744
rect 17678 7732 17684 7744
rect 17639 7704 17684 7732
rect 17678 7692 17684 7704
rect 17736 7692 17742 7744
rect 20714 7732 20720 7744
rect 20675 7704 20720 7732
rect 20714 7692 20720 7704
rect 20772 7692 20778 7744
rect 33502 7732 33508 7744
rect 33463 7704 33508 7732
rect 33502 7692 33508 7704
rect 33560 7692 33566 7744
rect 51166 7692 51172 7744
rect 51224 7732 51230 7744
rect 51537 7735 51595 7741
rect 51537 7732 51549 7735
rect 51224 7704 51549 7732
rect 51224 7692 51230 7704
rect 51537 7701 51549 7704
rect 51583 7701 51595 7735
rect 51537 7695 51595 7701
rect 1104 7642 59340 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 59340 7642
rect 1104 7568 59340 7590
rect 5350 7528 5356 7540
rect 5311 7500 5356 7528
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 21082 7528 21088 7540
rect 21043 7500 21088 7528
rect 21082 7488 21088 7500
rect 21140 7488 21146 7540
rect 25222 7528 25228 7540
rect 25183 7500 25228 7528
rect 25222 7488 25228 7500
rect 25280 7488 25286 7540
rect 28353 7531 28411 7537
rect 28353 7497 28365 7531
rect 28399 7528 28411 7531
rect 29086 7528 29092 7540
rect 28399 7500 29092 7528
rect 28399 7497 28411 7500
rect 28353 7491 28411 7497
rect 29086 7488 29092 7500
rect 29144 7488 29150 7540
rect 36725 7531 36783 7537
rect 36725 7497 36737 7531
rect 36771 7528 36783 7531
rect 37366 7528 37372 7540
rect 36771 7500 37372 7528
rect 36771 7497 36783 7500
rect 36725 7491 36783 7497
rect 37366 7488 37372 7500
rect 37424 7488 37430 7540
rect 40037 7531 40095 7537
rect 40037 7497 40049 7531
rect 40083 7528 40095 7531
rect 41414 7528 41420 7540
rect 40083 7500 41420 7528
rect 40083 7497 40095 7500
rect 40037 7491 40095 7497
rect 41414 7488 41420 7500
rect 41472 7488 41478 7540
rect 41874 7528 41880 7540
rect 41835 7500 41880 7528
rect 41874 7488 41880 7500
rect 41932 7488 41938 7540
rect 44174 7528 44180 7540
rect 44135 7500 44180 7528
rect 44174 7488 44180 7500
rect 44232 7488 44238 7540
rect 50341 7531 50399 7537
rect 50341 7497 50353 7531
rect 50387 7528 50399 7531
rect 50614 7528 50620 7540
rect 50387 7500 50620 7528
rect 50387 7497 50399 7500
rect 50341 7491 50399 7497
rect 50614 7488 50620 7500
rect 50672 7488 50678 7540
rect 54018 7488 54024 7540
rect 54076 7528 54082 7540
rect 54113 7531 54171 7537
rect 54113 7528 54125 7531
rect 54076 7500 54125 7528
rect 54076 7488 54082 7500
rect 54113 7497 54125 7500
rect 54159 7497 54171 7531
rect 55950 7528 55956 7540
rect 55911 7500 55956 7528
rect 54113 7491 54171 7497
rect 55950 7488 55956 7500
rect 56008 7488 56014 7540
rect 2308 7463 2366 7469
rect 2308 7429 2320 7463
rect 2354 7460 2366 7463
rect 3234 7460 3240 7472
rect 2354 7432 3240 7460
rect 2354 7429 2366 7432
rect 2308 7423 2366 7429
rect 3234 7420 3240 7432
rect 3292 7420 3298 7472
rect 4065 7463 4123 7469
rect 4065 7429 4077 7463
rect 4111 7460 4123 7463
rect 7190 7460 7196 7472
rect 4111 7432 7196 7460
rect 4111 7429 4123 7432
rect 4065 7423 4123 7429
rect 7190 7420 7196 7432
rect 7248 7420 7254 7472
rect 13164 7463 13222 7469
rect 13164 7429 13176 7463
rect 13210 7460 13222 7463
rect 13814 7460 13820 7472
rect 13210 7432 13820 7460
rect 13210 7429 13222 7432
rect 13164 7423 13222 7429
rect 13814 7420 13820 7432
rect 13872 7420 13878 7472
rect 15004 7463 15062 7469
rect 15004 7429 15016 7463
rect 15050 7460 15062 7463
rect 17678 7460 17684 7472
rect 15050 7432 17684 7460
rect 15050 7429 15062 7432
rect 15004 7423 15062 7429
rect 17678 7420 17684 7432
rect 17736 7420 17742 7472
rect 18132 7463 18190 7469
rect 18132 7429 18144 7463
rect 18178 7460 18190 7463
rect 20714 7460 20720 7472
rect 18178 7432 20720 7460
rect 18178 7429 18190 7432
rect 18132 7423 18190 7429
rect 20714 7420 20720 7432
rect 20772 7420 20778 7472
rect 24394 7460 24400 7472
rect 24044 7432 24400 7460
rect 1854 7352 1860 7404
rect 1912 7392 1918 7404
rect 2041 7395 2099 7401
rect 2041 7392 2053 7395
rect 1912 7364 2053 7392
rect 1912 7352 1918 7364
rect 2041 7361 2053 7364
rect 2087 7361 2099 7395
rect 2041 7355 2099 7361
rect 7000 7395 7058 7401
rect 7000 7361 7012 7395
rect 7046 7392 7058 7395
rect 8386 7392 8392 7404
rect 7046 7364 8392 7392
rect 7046 7361 7058 7364
rect 7000 7355 7058 7361
rect 8386 7352 8392 7364
rect 8444 7352 8450 7404
rect 8573 7395 8631 7401
rect 8573 7361 8585 7395
rect 8619 7392 8631 7395
rect 8662 7392 8668 7404
rect 8619 7364 8668 7392
rect 8619 7361 8631 7364
rect 8573 7355 8631 7361
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 8840 7395 8898 7401
rect 8840 7361 8852 7395
rect 8886 7392 8898 7395
rect 10778 7392 10784 7404
rect 8886 7364 10784 7392
rect 8886 7361 8898 7364
rect 8840 7355 8898 7361
rect 10778 7352 10784 7364
rect 10836 7352 10842 7404
rect 14737 7395 14795 7401
rect 14737 7361 14749 7395
rect 14783 7392 14795 7395
rect 14826 7392 14832 7404
rect 14783 7364 14832 7392
rect 14783 7361 14795 7364
rect 14737 7355 14795 7361
rect 14826 7352 14832 7364
rect 14884 7352 14890 7404
rect 17310 7352 17316 7404
rect 17368 7392 17374 7404
rect 17865 7395 17923 7401
rect 17865 7392 17877 7395
rect 17368 7364 17877 7392
rect 17368 7352 17374 7364
rect 17865 7361 17877 7364
rect 17911 7361 17923 7395
rect 17865 7355 17923 7361
rect 19972 7395 20030 7401
rect 19972 7361 19984 7395
rect 20018 7392 20030 7395
rect 21174 7392 21180 7404
rect 20018 7364 21180 7392
rect 20018 7361 20030 7364
rect 19972 7355 20030 7361
rect 21174 7352 21180 7364
rect 21232 7352 21238 7404
rect 24044 7392 24072 7432
rect 24394 7420 24400 7432
rect 24452 7420 24458 7472
rect 27240 7463 27298 7469
rect 27240 7429 27252 7463
rect 27286 7460 27298 7463
rect 28534 7460 28540 7472
rect 27286 7432 28540 7460
rect 27286 7429 27298 7432
rect 27240 7423 27298 7429
rect 28534 7420 28540 7432
rect 28592 7420 28598 7472
rect 29816 7463 29874 7469
rect 29816 7429 29828 7463
rect 29862 7460 29874 7463
rect 30926 7460 30932 7472
rect 29862 7432 30932 7460
rect 29862 7429 29874 7432
rect 29816 7423 29874 7429
rect 30926 7420 30932 7432
rect 30984 7420 30990 7472
rect 32392 7463 32450 7469
rect 32392 7429 32404 7463
rect 32438 7460 32450 7463
rect 33502 7460 33508 7472
rect 32438 7432 33508 7460
rect 32438 7429 32450 7432
rect 32392 7423 32450 7429
rect 33502 7420 33508 7432
rect 33560 7420 33566 7472
rect 35802 7460 35808 7472
rect 35360 7432 35808 7460
rect 35360 7404 35388 7432
rect 35802 7420 35808 7432
rect 35860 7420 35866 7472
rect 38924 7463 38982 7469
rect 38924 7429 38936 7463
rect 38970 7460 38982 7463
rect 40494 7460 40500 7472
rect 38970 7432 40500 7460
rect 38970 7429 38982 7432
rect 38924 7423 38982 7429
rect 40494 7420 40500 7432
rect 40552 7420 40558 7472
rect 43064 7463 43122 7469
rect 43064 7429 43076 7463
rect 43110 7460 43122 7463
rect 43806 7460 43812 7472
rect 43110 7432 43812 7460
rect 43110 7429 43122 7432
rect 43064 7423 43122 7429
rect 43806 7420 43812 7432
rect 43864 7420 43870 7472
rect 49228 7463 49286 7469
rect 49228 7429 49240 7463
rect 49274 7460 49286 7463
rect 50798 7460 50804 7472
rect 49274 7432 50804 7460
rect 49274 7429 49286 7432
rect 49228 7423 49286 7429
rect 50798 7420 50804 7432
rect 50856 7420 50862 7472
rect 52638 7420 52644 7472
rect 52696 7460 52702 7472
rect 52696 7432 54340 7460
rect 52696 7420 52702 7432
rect 23952 7364 24072 7392
rect 24112 7395 24170 7401
rect 5902 7284 5908 7336
rect 5960 7324 5966 7336
rect 6730 7324 6736 7336
rect 5960 7296 6736 7324
rect 5960 7284 5966 7296
rect 6730 7284 6736 7296
rect 6788 7284 6794 7336
rect 12897 7327 12955 7333
rect 12897 7293 12909 7327
rect 12943 7293 12955 7327
rect 19702 7324 19708 7336
rect 19663 7296 19708 7324
rect 12897 7287 12955 7293
rect 3421 7191 3479 7197
rect 3421 7157 3433 7191
rect 3467 7188 3479 7191
rect 4062 7188 4068 7200
rect 3467 7160 4068 7188
rect 3467 7157 3479 7160
rect 3421 7151 3479 7157
rect 4062 7148 4068 7160
rect 4120 7148 4126 7200
rect 8113 7191 8171 7197
rect 8113 7157 8125 7191
rect 8159 7188 8171 7191
rect 8846 7188 8852 7200
rect 8159 7160 8852 7188
rect 8159 7157 8171 7160
rect 8113 7151 8171 7157
rect 8846 7148 8852 7160
rect 8904 7148 8910 7200
rect 9950 7188 9956 7200
rect 9911 7160 9956 7188
rect 9950 7148 9956 7160
rect 10008 7148 10014 7200
rect 12158 7148 12164 7200
rect 12216 7188 12222 7200
rect 12912 7188 12940 7287
rect 19702 7284 19708 7296
rect 19760 7284 19766 7336
rect 23842 7324 23848 7336
rect 23755 7296 23848 7324
rect 23842 7284 23848 7296
rect 23900 7324 23906 7336
rect 23952 7324 23980 7364
rect 24112 7361 24124 7395
rect 24158 7392 24170 7395
rect 25774 7392 25780 7404
rect 24158 7364 25780 7392
rect 24158 7361 24170 7364
rect 24112 7355 24170 7361
rect 25774 7352 25780 7364
rect 25832 7352 25838 7404
rect 26970 7392 26976 7404
rect 26931 7364 26976 7392
rect 26970 7352 26976 7364
rect 27028 7352 27034 7404
rect 35342 7392 35348 7404
rect 35255 7364 35348 7392
rect 35342 7352 35348 7364
rect 35400 7352 35406 7404
rect 35612 7395 35670 7401
rect 35612 7361 35624 7395
rect 35658 7392 35670 7395
rect 39206 7392 39212 7404
rect 35658 7364 39212 7392
rect 35658 7361 35670 7364
rect 35612 7355 35670 7361
rect 39206 7352 39212 7364
rect 39264 7352 39270 7404
rect 40764 7395 40822 7401
rect 40764 7361 40776 7395
rect 40810 7392 40822 7395
rect 43530 7392 43536 7404
rect 40810 7364 43536 7392
rect 40810 7361 40822 7364
rect 40764 7355 40822 7361
rect 43530 7352 43536 7364
rect 43588 7352 43594 7404
rect 45916 7395 45974 7401
rect 45916 7361 45928 7395
rect 45962 7392 45974 7395
rect 47118 7392 47124 7404
rect 45962 7364 47124 7392
rect 45962 7361 45974 7364
rect 45916 7355 45974 7361
rect 47118 7352 47124 7364
rect 47176 7352 47182 7404
rect 51068 7395 51126 7401
rect 51068 7361 51080 7395
rect 51114 7392 51126 7395
rect 51534 7392 51540 7404
rect 51114 7364 51540 7392
rect 51114 7361 51126 7364
rect 51068 7355 51126 7361
rect 51534 7352 51540 7364
rect 51592 7352 51598 7404
rect 52730 7392 52736 7404
rect 52691 7364 52736 7392
rect 52730 7352 52736 7364
rect 52788 7352 52794 7404
rect 53000 7395 53058 7401
rect 53000 7361 53012 7395
rect 53046 7392 53058 7395
rect 54202 7392 54208 7404
rect 53046 7364 54208 7392
rect 53046 7361 53058 7364
rect 53000 7355 53058 7361
rect 54202 7352 54208 7364
rect 54260 7352 54266 7404
rect 54312 7392 54340 7432
rect 54386 7420 54392 7472
rect 54444 7460 54450 7472
rect 54818 7463 54876 7469
rect 54818 7460 54830 7463
rect 54444 7432 54830 7460
rect 54444 7420 54450 7432
rect 54818 7429 54830 7432
rect 54864 7429 54876 7463
rect 54818 7423 54876 7429
rect 54573 7395 54631 7401
rect 54573 7392 54585 7395
rect 54312 7364 54585 7392
rect 54573 7361 54585 7364
rect 54619 7392 54631 7395
rect 55306 7392 55312 7404
rect 54619 7364 55312 7392
rect 54619 7361 54631 7364
rect 54573 7355 54631 7361
rect 55306 7352 55312 7364
rect 55364 7352 55370 7404
rect 23900 7296 23980 7324
rect 23900 7284 23906 7296
rect 29178 7284 29184 7336
rect 29236 7324 29242 7336
rect 29549 7327 29607 7333
rect 29549 7324 29561 7327
rect 29236 7296 29561 7324
rect 29236 7284 29242 7296
rect 29549 7293 29561 7296
rect 29595 7293 29607 7327
rect 32122 7324 32128 7336
rect 32083 7296 32128 7324
rect 29549 7287 29607 7293
rect 32122 7284 32128 7296
rect 32180 7284 32186 7336
rect 38654 7324 38660 7336
rect 38615 7296 38660 7324
rect 38654 7284 38660 7296
rect 38712 7284 38718 7336
rect 40402 7284 40408 7336
rect 40460 7324 40466 7336
rect 40497 7327 40555 7333
rect 40497 7324 40509 7327
rect 40460 7296 40509 7324
rect 40460 7284 40466 7296
rect 40497 7293 40509 7296
rect 40543 7293 40555 7327
rect 42794 7324 42800 7336
rect 42755 7296 42800 7324
rect 40497 7287 40555 7293
rect 42794 7284 42800 7296
rect 42852 7284 42858 7336
rect 45646 7324 45652 7336
rect 45607 7296 45652 7324
rect 45646 7284 45652 7296
rect 45704 7284 45710 7336
rect 46842 7284 46848 7336
rect 46900 7324 46906 7336
rect 47486 7324 47492 7336
rect 46900 7296 47492 7324
rect 46900 7284 46906 7296
rect 47486 7284 47492 7296
rect 47544 7324 47550 7336
rect 48961 7327 49019 7333
rect 48961 7324 48973 7327
rect 47544 7296 48973 7324
rect 47544 7284 47550 7296
rect 48961 7293 48973 7296
rect 49007 7293 49019 7327
rect 48961 7287 49019 7293
rect 50154 7284 50160 7336
rect 50212 7324 50218 7336
rect 50801 7327 50859 7333
rect 50801 7324 50813 7327
rect 50212 7296 50813 7324
rect 50212 7284 50218 7296
rect 50801 7293 50813 7296
rect 50847 7293 50859 7327
rect 50801 7287 50859 7293
rect 30834 7216 30840 7268
rect 30892 7256 30898 7268
rect 30929 7259 30987 7265
rect 30929 7256 30941 7259
rect 30892 7228 30941 7256
rect 30892 7216 30898 7228
rect 30929 7225 30941 7228
rect 30975 7225 30987 7259
rect 30929 7219 30987 7225
rect 14090 7188 14096 7200
rect 12216 7160 14096 7188
rect 12216 7148 12222 7160
rect 14090 7148 14096 7160
rect 14148 7148 14154 7200
rect 14274 7188 14280 7200
rect 14235 7160 14280 7188
rect 14274 7148 14280 7160
rect 14332 7148 14338 7200
rect 16114 7188 16120 7200
rect 16075 7160 16120 7188
rect 16114 7148 16120 7160
rect 16172 7148 16178 7200
rect 19242 7188 19248 7200
rect 19203 7160 19248 7188
rect 19242 7148 19248 7160
rect 19300 7148 19306 7200
rect 32306 7148 32312 7200
rect 32364 7188 32370 7200
rect 33505 7191 33563 7197
rect 33505 7188 33517 7191
rect 32364 7160 33517 7188
rect 32364 7148 32370 7160
rect 33505 7157 33517 7160
rect 33551 7157 33563 7191
rect 33505 7151 33563 7157
rect 47029 7191 47087 7197
rect 47029 7157 47041 7191
rect 47075 7188 47087 7191
rect 47670 7188 47676 7200
rect 47075 7160 47676 7188
rect 47075 7157 47087 7160
rect 47029 7151 47087 7157
rect 47670 7148 47676 7160
rect 47728 7148 47734 7200
rect 52178 7188 52184 7200
rect 52139 7160 52184 7188
rect 52178 7148 52184 7160
rect 52236 7148 52242 7200
rect 1104 7098 59340 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 59340 7098
rect 1104 7024 59340 7046
rect 6546 6984 6552 6996
rect 6507 6956 6552 6984
rect 6546 6944 6552 6956
rect 6604 6944 6610 6996
rect 8386 6984 8392 6996
rect 8347 6956 8392 6984
rect 8386 6944 8392 6956
rect 8444 6944 8450 6996
rect 13078 6944 13084 6996
rect 13136 6984 13142 6996
rect 13541 6987 13599 6993
rect 13541 6984 13553 6987
rect 13136 6956 13553 6984
rect 13136 6944 13142 6956
rect 13541 6953 13553 6956
rect 13587 6953 13599 6987
rect 21174 6984 21180 6996
rect 21135 6956 21180 6984
rect 13541 6947 13599 6953
rect 21174 6944 21180 6956
rect 21232 6944 21238 6996
rect 25774 6984 25780 6996
rect 25735 6956 25780 6984
rect 25774 6944 25780 6956
rect 25832 6944 25838 6996
rect 39206 6984 39212 6996
rect 39167 6956 39212 6984
rect 39206 6944 39212 6956
rect 39264 6944 39270 6996
rect 47118 6984 47124 6996
rect 47079 6956 47124 6984
rect 47118 6944 47124 6956
rect 47176 6944 47182 6996
rect 51534 6984 51540 6996
rect 51495 6956 51540 6984
rect 51534 6944 51540 6956
rect 51592 6944 51598 6996
rect 54202 6984 54208 6996
rect 54163 6956 54208 6984
rect 54202 6944 54208 6956
rect 54260 6944 54266 6996
rect 56689 6987 56747 6993
rect 56689 6953 56701 6987
rect 56735 6984 56747 6987
rect 56778 6984 56784 6996
rect 56735 6956 56784 6984
rect 56735 6953 56747 6956
rect 56689 6947 56747 6953
rect 56778 6944 56784 6956
rect 56836 6944 56842 6996
rect 58529 6987 58587 6993
rect 58529 6953 58541 6987
rect 58575 6984 58587 6987
rect 59449 6987 59507 6993
rect 59449 6984 59461 6987
rect 58575 6956 59461 6984
rect 58575 6953 58587 6956
rect 58529 6947 58587 6953
rect 59449 6953 59461 6956
rect 59495 6953 59507 6987
rect 59449 6947 59507 6953
rect 14090 6808 14096 6860
rect 14148 6848 14154 6860
rect 14734 6848 14740 6860
rect 14148 6820 14740 6848
rect 14148 6808 14154 6820
rect 14734 6808 14740 6820
rect 14792 6848 14798 6860
rect 15105 6851 15163 6857
rect 15105 6848 15117 6851
rect 14792 6820 15117 6848
rect 14792 6808 14798 6820
rect 15105 6817 15117 6820
rect 15151 6817 15163 6851
rect 17310 6848 17316 6860
rect 17271 6820 17316 6848
rect 15105 6811 15163 6817
rect 17310 6808 17316 6820
rect 17368 6808 17374 6860
rect 24394 6848 24400 6860
rect 24355 6820 24400 6848
rect 24394 6808 24400 6820
rect 24452 6808 24458 6860
rect 28718 6808 28724 6860
rect 28776 6848 28782 6860
rect 29638 6848 29644 6860
rect 28776 6820 29644 6848
rect 28776 6808 28782 6820
rect 29638 6808 29644 6820
rect 29696 6808 29702 6860
rect 32122 6808 32128 6860
rect 32180 6848 32186 6860
rect 32677 6851 32735 6857
rect 32677 6848 32689 6851
rect 32180 6820 32689 6848
rect 32180 6808 32186 6820
rect 32677 6817 32689 6820
rect 32723 6817 32735 6851
rect 40586 6848 40592 6860
rect 40547 6820 40592 6848
rect 32677 6811 32735 6817
rect 40586 6808 40592 6820
rect 40644 6808 40650 6860
rect 52730 6808 52736 6860
rect 52788 6848 52794 6860
rect 52825 6851 52883 6857
rect 52825 6848 52837 6851
rect 52788 6820 52837 6848
rect 52788 6808 52794 6820
rect 52825 6817 52837 6820
rect 52871 6817 52883 6851
rect 52825 6811 52883 6817
rect 1857 6783 1915 6789
rect 1857 6749 1869 6783
rect 1903 6780 1915 6783
rect 1946 6780 1952 6792
rect 1903 6752 1952 6780
rect 1903 6749 1915 6752
rect 1857 6743 1915 6749
rect 1946 6740 1952 6752
rect 2004 6740 2010 6792
rect 5442 6789 5448 6792
rect 5169 6783 5227 6789
rect 5169 6749 5181 6783
rect 5215 6780 5227 6783
rect 5215 6752 5396 6780
rect 5215 6749 5227 6752
rect 5169 6743 5227 6749
rect 2124 6715 2182 6721
rect 2124 6681 2136 6715
rect 2170 6712 2182 6715
rect 5258 6712 5264 6724
rect 2170 6684 5264 6712
rect 2170 6681 2182 6684
rect 2124 6675 2182 6681
rect 5258 6672 5264 6684
rect 5316 6672 5322 6724
rect 5368 6712 5396 6752
rect 5436 6743 5448 6789
rect 5500 6780 5506 6792
rect 5500 6752 5536 6780
rect 5442 6740 5448 6743
rect 5500 6740 5506 6752
rect 6730 6740 6736 6792
rect 6788 6780 6794 6792
rect 7009 6783 7067 6789
rect 7009 6780 7021 6783
rect 6788 6752 7021 6780
rect 6788 6740 6794 6752
rect 7009 6749 7021 6752
rect 7055 6780 7067 6783
rect 8662 6780 8668 6792
rect 7055 6752 8668 6780
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 8662 6740 8668 6752
rect 8720 6740 8726 6792
rect 8938 6780 8944 6792
rect 8899 6752 8944 6780
rect 8938 6740 8944 6752
rect 8996 6780 9002 6792
rect 10686 6780 10692 6792
rect 8996 6752 10692 6780
rect 8996 6740 9002 6752
rect 10686 6740 10692 6752
rect 10744 6740 10750 6792
rect 11882 6740 11888 6792
rect 11940 6780 11946 6792
rect 12158 6780 12164 6792
rect 11940 6752 12164 6780
rect 11940 6740 11946 6752
rect 12158 6740 12164 6752
rect 12216 6740 12222 6792
rect 12428 6783 12486 6789
rect 12428 6749 12440 6783
rect 12474 6780 12486 6783
rect 14274 6780 14280 6792
rect 12474 6752 14280 6780
rect 12474 6749 12486 6752
rect 12428 6743 12486 6749
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 15372 6783 15430 6789
rect 15372 6749 15384 6783
rect 15418 6780 15430 6783
rect 16114 6780 16120 6792
rect 15418 6752 16120 6780
rect 15418 6749 15430 6752
rect 15372 6743 15430 6749
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 17580 6783 17638 6789
rect 17580 6749 17592 6783
rect 17626 6780 17638 6783
rect 19242 6780 19248 6792
rect 17626 6752 19248 6780
rect 17626 6749 17638 6752
rect 17580 6743 17638 6749
rect 19242 6740 19248 6752
rect 19300 6740 19306 6792
rect 19702 6740 19708 6792
rect 19760 6780 19766 6792
rect 19797 6783 19855 6789
rect 19797 6780 19809 6783
rect 19760 6752 19809 6780
rect 19760 6740 19766 6752
rect 19797 6749 19809 6752
rect 19843 6780 19855 6783
rect 22002 6780 22008 6792
rect 19843 6752 22008 6780
rect 19843 6749 19855 6752
rect 19797 6743 19855 6749
rect 22002 6740 22008 6752
rect 22060 6780 22066 6792
rect 22465 6783 22523 6789
rect 22465 6780 22477 6783
rect 22060 6752 22477 6780
rect 22060 6740 22066 6752
rect 22465 6749 22477 6752
rect 22511 6780 22523 6783
rect 24302 6780 24308 6792
rect 22511 6752 24308 6780
rect 22511 6749 22523 6752
rect 22465 6743 22523 6749
rect 24302 6740 24308 6752
rect 24360 6740 24366 6792
rect 27617 6783 27675 6789
rect 27617 6749 27629 6783
rect 27663 6780 27675 6783
rect 28810 6780 28816 6792
rect 27663 6752 28816 6780
rect 27663 6749 27675 6752
rect 27617 6743 27675 6749
rect 28810 6740 28816 6752
rect 28868 6780 28874 6792
rect 29178 6780 29184 6792
rect 28868 6752 29184 6780
rect 28868 6740 28874 6752
rect 29178 6740 29184 6752
rect 29236 6780 29242 6792
rect 30282 6780 30288 6792
rect 29236 6752 30288 6780
rect 29236 6740 29242 6752
rect 30282 6740 30288 6752
rect 30340 6780 30346 6792
rect 30837 6783 30895 6789
rect 30837 6780 30849 6783
rect 30340 6752 30849 6780
rect 30340 6740 30346 6752
rect 30837 6749 30849 6752
rect 30883 6749 30895 6783
rect 30837 6743 30895 6749
rect 31104 6783 31162 6789
rect 31104 6749 31116 6783
rect 31150 6780 31162 6783
rect 32306 6780 32312 6792
rect 31150 6752 32312 6780
rect 31150 6749 31162 6752
rect 31104 6743 31162 6749
rect 32306 6740 32312 6752
rect 32364 6740 32370 6792
rect 35802 6740 35808 6792
rect 35860 6780 35866 6792
rect 35989 6783 36047 6789
rect 35989 6780 36001 6783
rect 35860 6752 36001 6780
rect 35860 6740 35866 6752
rect 35989 6749 36001 6752
rect 36035 6749 36047 6783
rect 35989 6743 36047 6749
rect 37734 6740 37740 6792
rect 37792 6780 37798 6792
rect 37829 6783 37887 6789
rect 37829 6780 37841 6783
rect 37792 6752 37841 6780
rect 37792 6740 37798 6752
rect 37829 6749 37841 6752
rect 37875 6780 37887 6783
rect 38654 6780 38660 6792
rect 37875 6752 38660 6780
rect 37875 6749 37887 6752
rect 37829 6743 37887 6749
rect 38654 6740 38660 6752
rect 38712 6740 38718 6792
rect 43070 6780 43076 6792
rect 43031 6752 43076 6780
rect 43070 6740 43076 6752
rect 43128 6740 43134 6792
rect 43622 6780 43628 6792
rect 43272 6752 43628 6780
rect 5810 6712 5816 6724
rect 5368 6684 5816 6712
rect 5810 6672 5816 6684
rect 5868 6712 5874 6724
rect 6748 6712 6776 6740
rect 5868 6684 6776 6712
rect 7276 6715 7334 6721
rect 5868 6672 5874 6684
rect 7276 6681 7288 6715
rect 7322 6712 7334 6715
rect 7742 6712 7748 6724
rect 7322 6684 7748 6712
rect 7322 6681 7334 6684
rect 7276 6675 7334 6681
rect 7742 6672 7748 6684
rect 7800 6672 7806 6724
rect 9208 6715 9266 6721
rect 9208 6681 9220 6715
rect 9254 6712 9266 6715
rect 10226 6712 10232 6724
rect 9254 6684 10232 6712
rect 9254 6681 9266 6684
rect 9208 6675 9266 6681
rect 10226 6672 10232 6684
rect 10284 6672 10290 6724
rect 20064 6715 20122 6721
rect 20064 6681 20076 6715
rect 20110 6712 20122 6715
rect 20898 6712 20904 6724
rect 20110 6684 20904 6712
rect 20110 6681 20122 6684
rect 20064 6675 20122 6681
rect 20898 6672 20904 6684
rect 20956 6672 20962 6724
rect 22732 6715 22790 6721
rect 22732 6681 22744 6715
rect 22778 6712 22790 6715
rect 23474 6712 23480 6724
rect 22778 6684 23480 6712
rect 22778 6681 22790 6684
rect 22732 6675 22790 6681
rect 23474 6672 23480 6684
rect 23532 6672 23538 6724
rect 24664 6715 24722 6721
rect 24664 6681 24676 6715
rect 24710 6712 24722 6715
rect 25774 6712 25780 6724
rect 24710 6684 25780 6712
rect 24710 6681 24722 6684
rect 24664 6675 24722 6681
rect 25774 6672 25780 6684
rect 25832 6672 25838 6724
rect 27884 6715 27942 6721
rect 27884 6681 27896 6715
rect 27930 6712 27942 6715
rect 31018 6712 31024 6724
rect 27930 6684 31024 6712
rect 27930 6681 27942 6684
rect 27884 6675 27942 6681
rect 31018 6672 31024 6684
rect 31076 6672 31082 6724
rect 32922 6715 32980 6721
rect 32922 6712 32934 6715
rect 32232 6684 32934 6712
rect 3234 6644 3240 6656
rect 3195 6616 3240 6644
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 10318 6644 10324 6656
rect 10279 6616 10324 6644
rect 10318 6604 10324 6616
rect 10376 6604 10382 6656
rect 16485 6647 16543 6653
rect 16485 6613 16497 6647
rect 16531 6644 16543 6647
rect 16574 6644 16580 6656
rect 16531 6616 16580 6644
rect 16531 6613 16543 6616
rect 16485 6607 16543 6613
rect 16574 6604 16580 6616
rect 16632 6604 16638 6656
rect 18690 6644 18696 6656
rect 18651 6616 18696 6644
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 23842 6644 23848 6656
rect 23803 6616 23848 6644
rect 23842 6604 23848 6616
rect 23900 6604 23906 6656
rect 28994 6644 29000 6656
rect 28955 6616 29000 6644
rect 28994 6604 29000 6616
rect 29052 6604 29058 6656
rect 32232 6653 32260 6684
rect 32922 6681 32934 6684
rect 32968 6681 32980 6715
rect 32922 6675 32980 6681
rect 36256 6715 36314 6721
rect 36256 6681 36268 6715
rect 36302 6712 36314 6715
rect 36722 6712 36728 6724
rect 36302 6684 36728 6712
rect 36302 6681 36314 6684
rect 36256 6675 36314 6681
rect 36722 6672 36728 6684
rect 36780 6672 36786 6724
rect 38074 6715 38132 6721
rect 38074 6712 38086 6715
rect 37384 6684 38086 6712
rect 32217 6647 32275 6653
rect 32217 6613 32229 6647
rect 32263 6613 32275 6647
rect 34054 6644 34060 6656
rect 34015 6616 34060 6644
rect 32217 6607 32275 6613
rect 34054 6604 34060 6616
rect 34112 6604 34118 6656
rect 37384 6653 37412 6684
rect 38074 6681 38086 6684
rect 38120 6681 38132 6715
rect 38074 6675 38132 6681
rect 40856 6715 40914 6721
rect 40856 6681 40868 6715
rect 40902 6712 40914 6715
rect 43272 6712 43300 6752
rect 43622 6740 43628 6752
rect 43680 6740 43686 6792
rect 43898 6740 43904 6792
rect 43956 6780 43962 6792
rect 45646 6780 45652 6792
rect 43956 6752 45652 6780
rect 43956 6740 43962 6752
rect 45646 6740 45652 6752
rect 45704 6740 45710 6792
rect 45741 6783 45799 6789
rect 45741 6749 45753 6783
rect 45787 6780 45799 6783
rect 47486 6780 47492 6792
rect 45787 6752 47492 6780
rect 45787 6749 45799 6752
rect 45741 6743 45799 6749
rect 47486 6740 47492 6752
rect 47544 6780 47550 6792
rect 47854 6789 47860 6792
rect 47581 6783 47639 6789
rect 47581 6780 47593 6783
rect 47544 6752 47593 6780
rect 47544 6740 47550 6752
rect 47581 6749 47593 6752
rect 47627 6749 47639 6783
rect 47581 6743 47639 6749
rect 47848 6743 47860 6789
rect 47912 6780 47918 6792
rect 47912 6752 47948 6780
rect 47854 6740 47860 6743
rect 47912 6740 47918 6752
rect 49786 6740 49792 6792
rect 49844 6780 49850 6792
rect 50154 6780 50160 6792
rect 49844 6752 50160 6780
rect 49844 6740 49850 6752
rect 50154 6740 50160 6752
rect 50212 6740 50218 6792
rect 50424 6783 50482 6789
rect 50424 6749 50436 6783
rect 50470 6780 50482 6783
rect 51166 6780 51172 6792
rect 50470 6752 51172 6780
rect 50470 6749 50482 6752
rect 50424 6743 50482 6749
rect 51166 6740 51172 6752
rect 51224 6740 51230 6792
rect 55306 6780 55312 6792
rect 55219 6752 55312 6780
rect 55306 6740 55312 6752
rect 55364 6740 55370 6792
rect 55576 6783 55634 6789
rect 55576 6749 55588 6783
rect 55622 6780 55634 6783
rect 55858 6780 55864 6792
rect 55622 6752 55864 6780
rect 55622 6749 55634 6752
rect 55576 6743 55634 6749
rect 55858 6740 55864 6752
rect 55916 6740 55922 6792
rect 57149 6783 57207 6789
rect 57149 6749 57161 6783
rect 57195 6749 57207 6783
rect 57149 6743 57207 6749
rect 57416 6783 57474 6789
rect 57416 6749 57428 6783
rect 57462 6780 57474 6783
rect 58526 6780 58532 6792
rect 57462 6752 58532 6780
rect 57462 6749 57474 6752
rect 57416 6743 57474 6749
rect 40902 6684 43300 6712
rect 43340 6715 43398 6721
rect 40902 6681 40914 6684
rect 40856 6675 40914 6681
rect 43340 6681 43352 6715
rect 43386 6712 43398 6715
rect 45278 6712 45284 6724
rect 43386 6684 45284 6712
rect 43386 6681 43398 6684
rect 43340 6675 43398 6681
rect 45278 6672 45284 6684
rect 45336 6672 45342 6724
rect 46008 6715 46066 6721
rect 46008 6681 46020 6715
rect 46054 6712 46066 6715
rect 49326 6712 49332 6724
rect 46054 6684 49332 6712
rect 46054 6681 46066 6684
rect 46008 6675 46066 6681
rect 49326 6672 49332 6684
rect 49384 6672 49390 6724
rect 53092 6715 53150 6721
rect 53092 6681 53104 6715
rect 53138 6712 53150 6715
rect 54662 6712 54668 6724
rect 53138 6684 54668 6712
rect 53138 6681 53150 6684
rect 53092 6675 53150 6681
rect 54662 6672 54668 6684
rect 54720 6672 54726 6724
rect 55324 6712 55352 6740
rect 57164 6712 57192 6743
rect 58526 6740 58532 6752
rect 58584 6740 58590 6792
rect 55324 6684 57192 6712
rect 37369 6647 37427 6653
rect 37369 6613 37381 6647
rect 37415 6613 37427 6647
rect 41966 6644 41972 6656
rect 41927 6616 41972 6644
rect 37369 6607 37427 6613
rect 41966 6604 41972 6616
rect 42024 6604 42030 6656
rect 44450 6644 44456 6656
rect 44411 6616 44456 6644
rect 44450 6604 44456 6616
rect 44508 6604 44514 6656
rect 48958 6644 48964 6656
rect 48919 6616 48964 6644
rect 48958 6604 48964 6616
rect 49016 6604 49022 6656
rect 1104 6554 59340 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 59340 6554
rect 1104 6480 59340 6502
rect 5258 6440 5264 6452
rect 5219 6412 5264 6440
rect 5258 6400 5264 6412
rect 5316 6400 5322 6452
rect 8662 6440 8668 6452
rect 8623 6412 8668 6440
rect 8662 6400 8668 6412
rect 8720 6400 8726 6452
rect 10778 6440 10784 6452
rect 10739 6412 10784 6440
rect 10778 6400 10784 6412
rect 10836 6400 10842 6452
rect 12250 6400 12256 6452
rect 12308 6440 12314 6452
rect 13265 6443 13323 6449
rect 13265 6440 13277 6443
rect 12308 6412 13277 6440
rect 12308 6400 12314 6412
rect 13265 6409 13277 6412
rect 13311 6409 13323 6443
rect 13265 6403 13323 6409
rect 16022 6400 16028 6452
rect 16080 6440 16086 6452
rect 16117 6443 16175 6449
rect 16117 6440 16129 6443
rect 16080 6412 16129 6440
rect 16080 6400 16086 6412
rect 16117 6409 16129 6412
rect 16163 6409 16175 6443
rect 18322 6440 18328 6452
rect 18283 6412 18328 6440
rect 16117 6403 16175 6409
rect 18322 6400 18328 6412
rect 18380 6400 18386 6452
rect 20898 6440 20904 6452
rect 20859 6412 20904 6440
rect 20898 6400 20904 6412
rect 20956 6400 20962 6452
rect 23474 6440 23480 6452
rect 23435 6412 23480 6440
rect 23474 6400 23480 6412
rect 23532 6400 23538 6452
rect 25774 6440 25780 6452
rect 25735 6412 25780 6440
rect 25774 6400 25780 6412
rect 25832 6400 25838 6452
rect 36722 6440 36728 6452
rect 36683 6412 36728 6440
rect 36722 6400 36728 6412
rect 36780 6400 36786 6452
rect 41233 6443 41291 6449
rect 41233 6409 41245 6443
rect 41279 6409 41291 6443
rect 49326 6440 49332 6452
rect 49287 6412 49332 6440
rect 41233 6403 41291 6409
rect 2308 6375 2366 6381
rect 2308 6341 2320 6375
rect 2354 6372 2366 6375
rect 3234 6372 3240 6384
rect 2354 6344 3240 6372
rect 2354 6341 2366 6344
rect 2308 6335 2366 6341
rect 3234 6332 3240 6344
rect 3292 6332 3298 6384
rect 4154 6381 4160 6384
rect 4148 6335 4160 6381
rect 4212 6372 4218 6384
rect 4212 6344 4248 6372
rect 4154 6332 4160 6335
rect 4212 6332 4218 6344
rect 8846 6332 8852 6384
rect 8904 6372 8910 6384
rect 9646 6375 9704 6381
rect 9646 6372 9658 6375
rect 8904 6344 9658 6372
rect 8904 6332 8910 6344
rect 9646 6341 9658 6344
rect 9692 6341 9704 6375
rect 12152 6375 12210 6381
rect 9646 6335 9704 6341
rect 9784 6344 12020 6372
rect 1946 6264 1952 6316
rect 2004 6304 2010 6316
rect 2041 6307 2099 6313
rect 2041 6304 2053 6307
rect 2004 6276 2053 6304
rect 2004 6264 2010 6276
rect 2041 6273 2053 6276
rect 2087 6304 2099 6307
rect 3881 6307 3939 6313
rect 3881 6304 3893 6307
rect 2087 6276 3893 6304
rect 2087 6273 2099 6276
rect 2041 6267 2099 6273
rect 3881 6273 3893 6276
rect 3927 6304 3939 6307
rect 3970 6304 3976 6316
rect 3927 6276 3976 6304
rect 3927 6273 3939 6276
rect 3881 6267 3939 6273
rect 3970 6264 3976 6276
rect 4028 6264 4034 6316
rect 7190 6304 7196 6316
rect 7103 6276 7196 6304
rect 7190 6264 7196 6276
rect 7248 6304 7254 6316
rect 9784 6304 9812 6344
rect 11882 6304 11888 6316
rect 7248 6276 9812 6304
rect 11843 6276 11888 6304
rect 7248 6264 7254 6276
rect 11882 6264 11888 6276
rect 11940 6264 11946 6316
rect 11992 6304 12020 6344
rect 12152 6341 12164 6375
rect 12198 6372 12210 6375
rect 13538 6372 13544 6384
rect 12198 6344 13544 6372
rect 12198 6341 12210 6344
rect 12152 6335 12210 6341
rect 13538 6332 13544 6344
rect 13596 6332 13602 6384
rect 15004 6375 15062 6381
rect 15004 6341 15016 6375
rect 15050 6372 15062 6375
rect 15838 6372 15844 6384
rect 15050 6344 15844 6372
rect 15050 6341 15062 6344
rect 15004 6335 15062 6341
rect 15838 6332 15844 6344
rect 15896 6332 15902 6384
rect 17212 6375 17270 6381
rect 17212 6341 17224 6375
rect 17258 6372 17270 6375
rect 18690 6372 18696 6384
rect 17258 6344 18696 6372
rect 17258 6341 17270 6344
rect 17212 6335 17270 6341
rect 18690 6332 18696 6344
rect 18748 6332 18754 6384
rect 23842 6332 23848 6384
rect 23900 6372 23906 6384
rect 24642 6375 24700 6381
rect 24642 6372 24654 6375
rect 23900 6344 24654 6372
rect 23900 6332 23906 6344
rect 24642 6341 24654 6344
rect 24688 6341 24700 6375
rect 24642 6335 24700 6341
rect 30282 6332 30288 6384
rect 30340 6372 30346 6384
rect 32392 6375 32450 6381
rect 30340 6344 31064 6372
rect 30340 6332 30346 6344
rect 12434 6304 12440 6316
rect 11992 6276 12440 6304
rect 12434 6264 12440 6276
rect 12492 6264 12498 6316
rect 14734 6304 14740 6316
rect 14695 6276 14740 6304
rect 14734 6264 14740 6276
rect 14792 6264 14798 6316
rect 19788 6307 19846 6313
rect 19788 6273 19800 6307
rect 19834 6304 19846 6307
rect 20622 6304 20628 6316
rect 19834 6276 20628 6304
rect 19834 6273 19846 6276
rect 19788 6267 19846 6273
rect 20622 6264 20628 6276
rect 20680 6264 20686 6316
rect 22002 6264 22008 6316
rect 22060 6304 22066 6316
rect 22097 6307 22155 6313
rect 22097 6304 22109 6307
rect 22060 6276 22109 6304
rect 22060 6264 22066 6276
rect 22097 6273 22109 6276
rect 22143 6273 22155 6307
rect 22097 6267 22155 6273
rect 22364 6307 22422 6313
rect 22364 6273 22376 6307
rect 22410 6304 22422 6307
rect 23198 6304 23204 6316
rect 22410 6276 23204 6304
rect 22410 6273 22422 6276
rect 22364 6267 22422 6273
rect 23198 6264 23204 6276
rect 23256 6264 23262 6316
rect 27240 6307 27298 6313
rect 27240 6273 27252 6307
rect 27286 6304 27298 6307
rect 28902 6304 28908 6316
rect 27286 6276 28908 6304
rect 27286 6273 27298 6276
rect 27240 6267 27298 6273
rect 28902 6264 28908 6276
rect 28960 6264 28966 6316
rect 29638 6264 29644 6316
rect 29696 6304 29702 6316
rect 29733 6307 29791 6313
rect 29733 6304 29745 6307
rect 29696 6276 29745 6304
rect 29696 6264 29702 6276
rect 29733 6273 29745 6276
rect 29779 6273 29791 6307
rect 29733 6267 29791 6273
rect 30000 6307 30058 6313
rect 30000 6273 30012 6307
rect 30046 6304 30058 6307
rect 30926 6304 30932 6316
rect 30046 6276 30932 6304
rect 30046 6273 30058 6276
rect 30000 6267 30058 6273
rect 30926 6264 30932 6276
rect 30984 6264 30990 6316
rect 8938 6196 8944 6248
rect 8996 6236 9002 6248
rect 9401 6239 9459 6245
rect 9401 6236 9413 6239
rect 8996 6208 9413 6236
rect 8996 6196 9002 6208
rect 9401 6205 9413 6208
rect 9447 6205 9459 6239
rect 9401 6199 9459 6205
rect 16298 6196 16304 6248
rect 16356 6236 16362 6248
rect 16945 6239 17003 6245
rect 16945 6236 16957 6239
rect 16356 6208 16957 6236
rect 16356 6196 16362 6208
rect 16945 6205 16957 6208
rect 16991 6205 17003 6239
rect 16945 6199 17003 6205
rect 19426 6196 19432 6248
rect 19484 6236 19490 6248
rect 19521 6239 19579 6245
rect 19521 6236 19533 6239
rect 19484 6208 19533 6236
rect 19484 6196 19490 6208
rect 19521 6205 19533 6208
rect 19567 6205 19579 6239
rect 19521 6199 19579 6205
rect 24302 6196 24308 6248
rect 24360 6236 24366 6248
rect 24397 6239 24455 6245
rect 24397 6236 24409 6239
rect 24360 6208 24409 6236
rect 24360 6196 24366 6208
rect 24397 6205 24409 6208
rect 24443 6205 24455 6239
rect 26970 6236 26976 6248
rect 26931 6208 26976 6236
rect 24397 6199 24455 6205
rect 3421 6103 3479 6109
rect 3421 6069 3433 6103
rect 3467 6100 3479 6103
rect 4062 6100 4068 6112
rect 3467 6072 4068 6100
rect 3467 6069 3479 6072
rect 3421 6063 3479 6069
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 24412 6100 24440 6199
rect 26970 6196 26976 6208
rect 27028 6196 27034 6248
rect 31036 6236 31064 6344
rect 32392 6341 32404 6375
rect 32438 6372 32450 6375
rect 34054 6372 34060 6384
rect 32438 6344 34060 6372
rect 32438 6341 32450 6344
rect 32392 6335 32450 6341
rect 34054 6332 34060 6344
rect 34112 6332 34118 6384
rect 38280 6375 38338 6381
rect 38280 6341 38292 6375
rect 38326 6372 38338 6375
rect 41248 6372 41276 6403
rect 49326 6400 49332 6412
rect 49384 6400 49390 6452
rect 54662 6440 54668 6452
rect 54623 6412 54668 6440
rect 54662 6400 54668 6412
rect 54720 6400 54726 6452
rect 38326 6344 41276 6372
rect 48216 6375 48274 6381
rect 38326 6341 38338 6344
rect 38280 6335 38338 6341
rect 48216 6341 48228 6375
rect 48262 6372 48274 6375
rect 48958 6372 48964 6384
rect 48262 6344 48964 6372
rect 48262 6341 48274 6344
rect 48216 6335 48274 6341
rect 48958 6332 48964 6344
rect 49016 6332 49022 6384
rect 50056 6375 50114 6381
rect 50056 6341 50068 6375
rect 50102 6372 50114 6375
rect 52178 6372 52184 6384
rect 50102 6344 52184 6372
rect 50102 6341 50114 6344
rect 50056 6335 50114 6341
rect 52178 6332 52184 6344
rect 52236 6332 52242 6384
rect 35612 6307 35670 6313
rect 35612 6273 35624 6307
rect 35658 6304 35670 6307
rect 36722 6304 36728 6316
rect 35658 6276 36728 6304
rect 35658 6273 35670 6276
rect 35612 6267 35670 6273
rect 36722 6264 36728 6276
rect 36780 6264 36786 6316
rect 40120 6307 40178 6313
rect 40120 6273 40132 6307
rect 40166 6304 40178 6307
rect 41690 6304 41696 6316
rect 40166 6276 41696 6304
rect 40166 6273 40178 6276
rect 40120 6267 40178 6273
rect 41690 6264 41696 6276
rect 41748 6264 41754 6316
rect 43070 6264 43076 6316
rect 43128 6304 43134 6316
rect 43809 6307 43867 6313
rect 43809 6304 43821 6307
rect 43128 6276 43821 6304
rect 43128 6264 43134 6276
rect 43809 6273 43821 6276
rect 43855 6304 43867 6307
rect 43898 6304 43904 6316
rect 43855 6276 43904 6304
rect 43855 6273 43867 6276
rect 43809 6267 43867 6273
rect 43898 6264 43904 6276
rect 43956 6264 43962 6316
rect 44076 6307 44134 6313
rect 44076 6273 44088 6307
rect 44122 6304 44134 6307
rect 45370 6304 45376 6316
rect 44122 6276 45376 6304
rect 44122 6273 44134 6276
rect 44076 6267 44134 6273
rect 45370 6264 45376 6276
rect 45428 6264 45434 6316
rect 45916 6307 45974 6313
rect 45916 6273 45928 6307
rect 45962 6304 45974 6307
rect 47394 6304 47400 6316
rect 45962 6276 47400 6304
rect 45962 6273 45974 6276
rect 45916 6267 45974 6273
rect 47394 6264 47400 6276
rect 47452 6264 47458 6316
rect 47486 6264 47492 6316
rect 47544 6304 47550 6316
rect 47949 6307 48007 6313
rect 47949 6304 47961 6307
rect 47544 6276 47961 6304
rect 47544 6264 47550 6276
rect 47949 6273 47961 6276
rect 47995 6273 48007 6307
rect 49786 6304 49792 6316
rect 47949 6267 48007 6273
rect 48056 6276 49792 6304
rect 32122 6236 32128 6248
rect 31036 6208 32128 6236
rect 32122 6196 32128 6208
rect 32180 6196 32186 6248
rect 35342 6236 35348 6248
rect 35303 6208 35348 6236
rect 35342 6196 35348 6208
rect 35400 6196 35406 6248
rect 37734 6196 37740 6248
rect 37792 6236 37798 6248
rect 38013 6239 38071 6245
rect 38013 6236 38025 6239
rect 37792 6208 38025 6236
rect 37792 6196 37798 6208
rect 38013 6205 38025 6208
rect 38059 6205 38071 6239
rect 38013 6199 38071 6205
rect 39853 6239 39911 6245
rect 39853 6205 39865 6239
rect 39899 6205 39911 6239
rect 39853 6199 39911 6205
rect 45649 6239 45707 6245
rect 45649 6205 45661 6239
rect 45695 6205 45707 6239
rect 48056 6236 48084 6276
rect 49786 6264 49792 6276
rect 49844 6264 49850 6316
rect 53552 6307 53610 6313
rect 53552 6273 53564 6307
rect 53598 6304 53610 6307
rect 54110 6304 54116 6316
rect 53598 6276 54116 6304
rect 53598 6273 53610 6276
rect 53552 6267 53610 6273
rect 54110 6264 54116 6276
rect 54168 6264 54174 6316
rect 45649 6199 45707 6205
rect 46860 6208 48084 6236
rect 24670 6100 24676 6112
rect 24412 6072 24676 6100
rect 24670 6060 24676 6072
rect 24728 6060 24734 6112
rect 26050 6060 26056 6112
rect 26108 6100 26114 6112
rect 28353 6103 28411 6109
rect 28353 6100 28365 6103
rect 26108 6072 28365 6100
rect 26108 6060 26114 6072
rect 28353 6069 28365 6072
rect 28399 6069 28411 6103
rect 31110 6100 31116 6112
rect 31071 6072 31116 6100
rect 28353 6063 28411 6069
rect 31110 6060 31116 6072
rect 31168 6060 31174 6112
rect 33502 6100 33508 6112
rect 33463 6072 33508 6100
rect 33502 6060 33508 6072
rect 33560 6060 33566 6112
rect 39390 6100 39396 6112
rect 39351 6072 39396 6100
rect 39390 6060 39396 6072
rect 39448 6060 39454 6112
rect 39868 6100 39896 6199
rect 40218 6100 40224 6112
rect 39868 6072 40224 6100
rect 40218 6060 40224 6072
rect 40276 6100 40282 6112
rect 40586 6100 40592 6112
rect 40276 6072 40592 6100
rect 40276 6060 40282 6072
rect 40586 6060 40592 6072
rect 40644 6060 40650 6112
rect 43346 6060 43352 6112
rect 43404 6100 43410 6112
rect 45189 6103 45247 6109
rect 45189 6100 45201 6103
rect 43404 6072 45201 6100
rect 43404 6060 43410 6072
rect 45189 6069 45201 6072
rect 45235 6069 45247 6103
rect 45664 6100 45692 6199
rect 46860 6112 46888 6208
rect 52730 6196 52736 6248
rect 52788 6236 52794 6248
rect 53285 6239 53343 6245
rect 53285 6236 53297 6239
rect 52788 6208 53297 6236
rect 52788 6196 52794 6208
rect 53285 6205 53297 6208
rect 53331 6205 53343 6239
rect 53285 6199 53343 6205
rect 46842 6100 46848 6112
rect 45664 6072 46848 6100
rect 45189 6063 45247 6069
rect 46842 6060 46848 6072
rect 46900 6060 46906 6112
rect 47026 6100 47032 6112
rect 46987 6072 47032 6100
rect 47026 6060 47032 6072
rect 47084 6060 47090 6112
rect 51166 6100 51172 6112
rect 51127 6072 51172 6100
rect 51166 6060 51172 6072
rect 51224 6060 51230 6112
rect 1104 6010 59340 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 59340 6010
rect 1104 5936 59340 5958
rect 10226 5856 10232 5908
rect 10284 5896 10290 5908
rect 10321 5899 10379 5905
rect 10321 5896 10333 5899
rect 10284 5868 10333 5896
rect 10284 5856 10290 5868
rect 10321 5865 10333 5868
rect 10367 5865 10379 5899
rect 10321 5859 10379 5865
rect 16206 5856 16212 5908
rect 16264 5896 16270 5908
rect 17681 5899 17739 5905
rect 17681 5896 17693 5899
rect 16264 5868 17693 5896
rect 16264 5856 16270 5868
rect 17681 5865 17693 5868
rect 17727 5865 17739 5899
rect 20622 5896 20628 5908
rect 20583 5868 20628 5896
rect 17681 5859 17739 5865
rect 20622 5856 20628 5868
rect 20680 5856 20686 5908
rect 23198 5896 23204 5908
rect 23159 5868 23204 5896
rect 23198 5856 23204 5868
rect 23256 5856 23262 5908
rect 26970 5856 26976 5908
rect 27028 5896 27034 5908
rect 27028 5868 28580 5896
rect 27028 5856 27034 5868
rect 3970 5760 3976 5772
rect 3931 5732 3976 5760
rect 3970 5720 3976 5732
rect 4028 5720 4034 5772
rect 5810 5760 5816 5772
rect 5771 5732 5816 5760
rect 5810 5720 5816 5732
rect 5868 5720 5874 5772
rect 8938 5760 8944 5772
rect 8899 5732 8944 5760
rect 8938 5720 8944 5732
rect 8996 5720 9002 5772
rect 10686 5720 10692 5772
rect 10744 5760 10750 5772
rect 10781 5763 10839 5769
rect 10781 5760 10793 5763
rect 10744 5732 10793 5760
rect 10744 5720 10750 5732
rect 10781 5729 10793 5732
rect 10827 5729 10839 5763
rect 16298 5760 16304 5772
rect 16259 5732 16304 5760
rect 10781 5723 10839 5729
rect 16298 5720 16304 5732
rect 16356 5720 16362 5772
rect 27632 5769 27660 5868
rect 28552 5828 28580 5868
rect 28902 5856 28908 5908
rect 28960 5896 28966 5908
rect 28997 5899 29055 5905
rect 28997 5896 29009 5899
rect 28960 5868 29009 5896
rect 28960 5856 28966 5868
rect 28997 5865 29009 5868
rect 29043 5865 29055 5899
rect 29730 5896 29736 5908
rect 28997 5859 29055 5865
rect 29104 5868 29736 5896
rect 29104 5828 29132 5868
rect 29730 5856 29736 5868
rect 29788 5856 29794 5908
rect 30926 5896 30932 5908
rect 30887 5868 30932 5896
rect 30926 5856 30932 5868
rect 30984 5856 30990 5908
rect 35342 5856 35348 5908
rect 35400 5896 35406 5908
rect 35802 5896 35808 5908
rect 35400 5868 35808 5896
rect 35400 5856 35406 5868
rect 35802 5856 35808 5868
rect 35860 5896 35866 5908
rect 36357 5899 36415 5905
rect 36357 5896 36369 5899
rect 35860 5868 36369 5896
rect 35860 5856 35866 5868
rect 36357 5865 36369 5868
rect 36403 5865 36415 5899
rect 36357 5859 36415 5865
rect 39390 5856 39396 5908
rect 39448 5896 39454 5908
rect 41506 5896 41512 5908
rect 39448 5868 41512 5896
rect 39448 5856 39454 5868
rect 41506 5856 41512 5868
rect 41564 5856 41570 5908
rect 41690 5896 41696 5908
rect 41651 5868 41696 5896
rect 41690 5856 41696 5868
rect 41748 5856 41754 5908
rect 52730 5896 52736 5908
rect 52691 5868 52736 5896
rect 52730 5856 52736 5868
rect 52788 5856 52794 5908
rect 28552 5800 29132 5828
rect 27617 5763 27675 5769
rect 27617 5729 27629 5763
rect 27663 5729 27675 5763
rect 27617 5723 27675 5729
rect 29178 5720 29184 5772
rect 29236 5760 29242 5772
rect 29549 5763 29607 5769
rect 29549 5760 29561 5763
rect 29236 5732 29561 5760
rect 29236 5720 29242 5732
rect 29549 5729 29561 5732
rect 29595 5729 29607 5763
rect 29549 5723 29607 5729
rect 32122 5720 32128 5772
rect 32180 5760 32186 5772
rect 32677 5763 32735 5769
rect 32677 5760 32689 5763
rect 32180 5732 32689 5760
rect 32180 5720 32186 5732
rect 32677 5729 32689 5732
rect 32723 5729 32735 5763
rect 32677 5723 32735 5729
rect 40218 5720 40224 5772
rect 40276 5760 40282 5772
rect 40313 5763 40371 5769
rect 40313 5760 40325 5763
rect 40276 5732 40325 5760
rect 40276 5720 40282 5732
rect 40313 5729 40325 5732
rect 40359 5729 40371 5763
rect 40313 5723 40371 5729
rect 48038 5720 48044 5772
rect 48096 5760 48102 5772
rect 48096 5732 51488 5760
rect 48096 5720 48102 5732
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 4229 5695 4287 5701
rect 4229 5692 4241 5695
rect 4120 5664 4241 5692
rect 4120 5652 4126 5664
rect 4229 5661 4241 5664
rect 4275 5661 4287 5695
rect 4229 5655 4287 5661
rect 9208 5695 9266 5701
rect 9208 5661 9220 5695
rect 9254 5692 9266 5695
rect 9950 5692 9956 5704
rect 9254 5664 9956 5692
rect 9254 5661 9266 5664
rect 9208 5655 9266 5661
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 13722 5652 13728 5704
rect 13780 5692 13786 5704
rect 16574 5701 16580 5704
rect 14461 5695 14519 5701
rect 14461 5692 14473 5695
rect 13780 5664 14473 5692
rect 13780 5652 13786 5664
rect 14461 5661 14473 5664
rect 14507 5661 14519 5695
rect 14461 5655 14519 5661
rect 16568 5655 16580 5701
rect 16632 5692 16638 5704
rect 19245 5695 19303 5701
rect 16632 5664 16668 5692
rect 16574 5652 16580 5655
rect 16632 5652 16638 5664
rect 19245 5661 19257 5695
rect 19291 5692 19303 5695
rect 21821 5695 21879 5701
rect 21821 5692 21833 5695
rect 19291 5664 21833 5692
rect 19291 5661 19303 5664
rect 19245 5655 19303 5661
rect 21821 5661 21833 5664
rect 21867 5692 21879 5695
rect 21910 5692 21916 5704
rect 21867 5664 21916 5692
rect 21867 5661 21879 5664
rect 21821 5655 21879 5661
rect 21910 5652 21916 5664
rect 21968 5652 21974 5704
rect 24670 5652 24676 5704
rect 24728 5692 24734 5704
rect 26050 5701 26056 5704
rect 25777 5695 25835 5701
rect 25777 5692 25789 5695
rect 24728 5664 25789 5692
rect 24728 5652 24734 5664
rect 25777 5661 25789 5664
rect 25823 5661 25835 5695
rect 25777 5655 25835 5661
rect 26044 5655 26056 5701
rect 26108 5692 26114 5704
rect 27884 5695 27942 5701
rect 26108 5664 26144 5692
rect 26050 5652 26056 5655
rect 26108 5652 26114 5664
rect 27884 5661 27896 5695
rect 27930 5692 27942 5695
rect 28994 5692 29000 5704
rect 27930 5664 29000 5692
rect 27930 5661 27942 5664
rect 27884 5655 27942 5661
rect 28994 5652 29000 5664
rect 29052 5652 29058 5704
rect 32944 5695 33002 5701
rect 32944 5661 32956 5695
rect 32990 5692 33002 5695
rect 33502 5692 33508 5704
rect 32990 5664 33508 5692
rect 32990 5661 33002 5664
rect 32944 5655 33002 5661
rect 33502 5652 33508 5664
rect 33560 5652 33566 5704
rect 37734 5652 37740 5704
rect 37792 5692 37798 5704
rect 37921 5695 37979 5701
rect 37921 5692 37933 5695
rect 37792 5664 37933 5692
rect 37792 5652 37798 5664
rect 37921 5661 37933 5664
rect 37967 5661 37979 5695
rect 37921 5655 37979 5661
rect 38188 5695 38246 5701
rect 38188 5661 38200 5695
rect 38234 5692 38246 5695
rect 38234 5664 42748 5692
rect 38234 5661 38246 5664
rect 38188 5655 38246 5661
rect 6086 5633 6092 5636
rect 6080 5587 6092 5633
rect 6144 5624 6150 5636
rect 11054 5633 11060 5636
rect 6144 5596 6180 5624
rect 6086 5584 6092 5587
rect 6144 5584 6150 5596
rect 11048 5587 11060 5633
rect 11112 5624 11118 5636
rect 14728 5627 14786 5633
rect 11112 5596 11148 5624
rect 11054 5584 11060 5587
rect 11112 5584 11118 5596
rect 14728 5593 14740 5627
rect 14774 5624 14786 5627
rect 15470 5624 15476 5636
rect 14774 5596 15476 5624
rect 14774 5593 14786 5596
rect 14728 5587 14786 5593
rect 15470 5584 15476 5596
rect 15528 5584 15534 5636
rect 19512 5627 19570 5633
rect 19512 5593 19524 5627
rect 19558 5624 19570 5627
rect 22088 5627 22146 5633
rect 19558 5596 22048 5624
rect 19558 5593 19570 5596
rect 19512 5587 19570 5593
rect 5350 5556 5356 5568
rect 5311 5528 5356 5556
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 7190 5556 7196 5568
rect 7151 5528 7196 5556
rect 7190 5516 7196 5528
rect 7248 5516 7254 5568
rect 11146 5516 11152 5568
rect 11204 5556 11210 5568
rect 12161 5559 12219 5565
rect 12161 5556 12173 5559
rect 11204 5528 12173 5556
rect 11204 5516 11210 5528
rect 12161 5525 12173 5528
rect 12207 5525 12219 5559
rect 12161 5519 12219 5525
rect 15841 5559 15899 5565
rect 15841 5525 15853 5559
rect 15887 5556 15899 5559
rect 16758 5556 16764 5568
rect 15887 5528 16764 5556
rect 15887 5525 15899 5528
rect 15841 5519 15899 5525
rect 16758 5516 16764 5528
rect 16816 5516 16822 5568
rect 22020 5556 22048 5596
rect 22088 5593 22100 5627
rect 22134 5624 22146 5627
rect 23290 5624 23296 5636
rect 22134 5596 23296 5624
rect 22134 5593 22146 5596
rect 22088 5587 22146 5593
rect 23290 5584 23296 5596
rect 23348 5584 23354 5636
rect 29638 5624 29644 5636
rect 26206 5596 29644 5624
rect 26206 5556 26234 5596
rect 29638 5584 29644 5596
rect 29696 5584 29702 5636
rect 29816 5627 29874 5633
rect 29816 5593 29828 5627
rect 29862 5624 29874 5627
rect 35069 5627 35127 5633
rect 29862 5596 34192 5624
rect 29862 5593 29874 5596
rect 29816 5587 29874 5593
rect 22020 5528 26234 5556
rect 27157 5559 27215 5565
rect 27157 5525 27169 5559
rect 27203 5556 27215 5559
rect 27246 5556 27252 5568
rect 27203 5528 27252 5556
rect 27203 5525 27215 5528
rect 27157 5519 27215 5525
rect 27246 5516 27252 5528
rect 27304 5516 27310 5568
rect 34054 5556 34060 5568
rect 34015 5528 34060 5556
rect 34054 5516 34060 5528
rect 34112 5516 34118 5568
rect 34164 5556 34192 5596
rect 35069 5593 35081 5627
rect 35115 5624 35127 5627
rect 40580 5627 40638 5633
rect 35115 5596 38148 5624
rect 35115 5593 35127 5596
rect 35069 5587 35127 5593
rect 35986 5556 35992 5568
rect 34164 5528 35992 5556
rect 35986 5516 35992 5528
rect 36044 5516 36050 5568
rect 38120 5556 38148 5596
rect 40580 5593 40592 5627
rect 40626 5624 40638 5627
rect 41230 5624 41236 5636
rect 40626 5596 41236 5624
rect 40626 5593 40638 5596
rect 40580 5587 40638 5593
rect 41230 5584 41236 5596
rect 41288 5584 41294 5636
rect 42720 5624 42748 5664
rect 42794 5652 42800 5704
rect 42852 5692 42858 5704
rect 43346 5701 43352 5704
rect 43073 5695 43131 5701
rect 43073 5692 43085 5695
rect 42852 5664 43085 5692
rect 42852 5652 42858 5664
rect 43073 5661 43085 5664
rect 43119 5661 43131 5695
rect 43340 5692 43352 5701
rect 43307 5664 43352 5692
rect 43073 5655 43131 5661
rect 43340 5655 43352 5664
rect 43346 5652 43352 5655
rect 43404 5652 43410 5704
rect 43898 5652 43904 5704
rect 43956 5692 43962 5704
rect 45005 5695 45063 5701
rect 45005 5692 45017 5695
rect 43956 5664 45017 5692
rect 43956 5652 43962 5664
rect 45005 5661 45017 5664
rect 45051 5661 45063 5695
rect 45005 5655 45063 5661
rect 45272 5695 45330 5701
rect 45272 5661 45284 5695
rect 45318 5692 45330 5695
rect 49602 5692 49608 5704
rect 45318 5664 49608 5692
rect 45318 5661 45330 5664
rect 45272 5655 45330 5661
rect 43806 5624 43812 5636
rect 42720 5596 43812 5624
rect 43806 5584 43812 5596
rect 43864 5584 43870 5636
rect 45020 5624 45048 5655
rect 49602 5652 49608 5664
rect 49660 5652 49666 5704
rect 51460 5701 51488 5732
rect 51445 5695 51503 5701
rect 51445 5661 51457 5695
rect 51491 5692 51503 5695
rect 53834 5692 53840 5704
rect 51491 5664 53840 5692
rect 51491 5661 51503 5664
rect 51445 5655 51503 5661
rect 53834 5652 53840 5664
rect 53892 5652 53898 5704
rect 46845 5627 46903 5633
rect 45020 5596 46796 5624
rect 39206 5556 39212 5568
rect 38120 5528 39212 5556
rect 39206 5516 39212 5528
rect 39264 5516 39270 5568
rect 39301 5559 39359 5565
rect 39301 5525 39313 5559
rect 39347 5556 39359 5559
rect 42702 5556 42708 5568
rect 39347 5528 42708 5556
rect 39347 5525 39359 5528
rect 39301 5519 39359 5525
rect 42702 5516 42708 5528
rect 42760 5516 42766 5568
rect 44266 5516 44272 5568
rect 44324 5556 44330 5568
rect 44453 5559 44511 5565
rect 44453 5556 44465 5559
rect 44324 5528 44465 5556
rect 44324 5516 44330 5528
rect 44453 5525 44465 5528
rect 44499 5525 44511 5559
rect 46382 5556 46388 5568
rect 46343 5528 46388 5556
rect 44453 5519 44511 5525
rect 46382 5516 46388 5528
rect 46440 5516 46446 5568
rect 46768 5556 46796 5596
rect 46845 5593 46857 5627
rect 46891 5624 46903 5627
rect 48038 5624 48044 5636
rect 46891 5596 48044 5624
rect 46891 5593 46903 5596
rect 46845 5587 46903 5593
rect 48038 5584 48044 5596
rect 48096 5584 48102 5636
rect 48133 5559 48191 5565
rect 48133 5556 48145 5559
rect 46768 5528 48145 5556
rect 48133 5525 48145 5528
rect 48179 5556 48191 5559
rect 48222 5556 48228 5568
rect 48179 5528 48228 5556
rect 48179 5525 48191 5528
rect 48133 5519 48191 5525
rect 48222 5516 48228 5528
rect 48280 5516 48286 5568
rect 1104 5466 59340 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 59340 5466
rect 1104 5392 59340 5414
rect 3789 5355 3847 5361
rect 3789 5321 3801 5355
rect 3835 5321 3847 5355
rect 3789 5315 3847 5321
rect 10597 5355 10655 5361
rect 10597 5321 10609 5355
rect 10643 5352 10655 5355
rect 11054 5352 11060 5364
rect 10643 5324 11060 5352
rect 10643 5321 10655 5324
rect 10597 5315 10655 5321
rect 3804 5284 3832 5315
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 44450 5352 44456 5364
rect 35866 5324 44456 5352
rect 4494 5287 4552 5293
rect 4494 5284 4506 5287
rect 3804 5256 4506 5284
rect 4494 5253 4506 5256
rect 4540 5253 4552 5287
rect 4494 5247 4552 5253
rect 6632 5287 6690 5293
rect 6632 5253 6644 5287
rect 6678 5284 6690 5287
rect 7190 5284 7196 5296
rect 6678 5256 7196 5284
rect 6678 5253 6690 5256
rect 6632 5247 6690 5253
rect 7190 5244 7196 5256
rect 7248 5244 7254 5296
rect 9484 5287 9542 5293
rect 9484 5253 9496 5287
rect 9530 5284 9542 5287
rect 10318 5284 10324 5296
rect 9530 5256 10324 5284
rect 9530 5253 9542 5256
rect 9484 5247 9542 5253
rect 10318 5244 10324 5256
rect 10376 5244 10382 5296
rect 11977 5287 12035 5293
rect 11977 5253 11989 5287
rect 12023 5284 12035 5287
rect 12434 5284 12440 5296
rect 12023 5256 12440 5284
rect 12023 5253 12035 5256
rect 11977 5247 12035 5253
rect 12434 5244 12440 5256
rect 12492 5244 12498 5296
rect 20156 5287 20214 5293
rect 20156 5253 20168 5287
rect 20202 5284 20214 5287
rect 25774 5284 25780 5296
rect 20202 5256 25780 5284
rect 20202 5253 20214 5256
rect 20156 5247 20214 5253
rect 25774 5244 25780 5256
rect 25832 5244 25838 5296
rect 29730 5284 29736 5296
rect 29691 5256 29736 5284
rect 29730 5244 29736 5256
rect 29788 5244 29794 5296
rect 32760 5287 32818 5293
rect 32760 5253 32772 5287
rect 32806 5284 32818 5287
rect 34054 5284 34060 5296
rect 32806 5256 34060 5284
rect 32806 5253 32818 5256
rect 32760 5247 32818 5253
rect 34054 5244 34060 5256
rect 34112 5244 34118 5296
rect 35428 5287 35486 5293
rect 35428 5253 35440 5287
rect 35474 5284 35486 5287
rect 35866 5284 35894 5324
rect 44450 5312 44456 5324
rect 44508 5312 44514 5364
rect 45370 5352 45376 5364
rect 45331 5324 45376 5352
rect 45370 5312 45376 5324
rect 45428 5312 45434 5364
rect 51537 5355 51595 5361
rect 51537 5352 51549 5355
rect 48700 5324 51549 5352
rect 35474 5256 35894 5284
rect 35474 5253 35486 5256
rect 35428 5247 35486 5253
rect 39206 5244 39212 5296
rect 39264 5284 39270 5296
rect 39577 5287 39635 5293
rect 39577 5284 39589 5287
rect 39264 5256 39589 5284
rect 39264 5244 39270 5256
rect 39577 5253 39589 5256
rect 39623 5284 39635 5287
rect 39850 5284 39856 5296
rect 39623 5256 39856 5284
rect 39623 5253 39635 5256
rect 39577 5247 39635 5253
rect 39850 5244 39856 5256
rect 39908 5244 39914 5296
rect 44260 5287 44318 5293
rect 44260 5253 44272 5287
rect 44306 5284 44318 5287
rect 46382 5284 46388 5296
rect 44306 5256 46388 5284
rect 44306 5253 44318 5256
rect 44260 5247 44318 5253
rect 46382 5244 46388 5256
rect 46440 5244 46446 5296
rect 48584 5287 48642 5293
rect 48584 5253 48596 5287
rect 48630 5284 48642 5287
rect 48700 5284 48728 5324
rect 51537 5321 51549 5324
rect 51583 5321 51595 5355
rect 51537 5315 51595 5321
rect 54110 5312 54116 5364
rect 54168 5352 54174 5364
rect 54205 5355 54263 5361
rect 54205 5352 54217 5355
rect 54168 5324 54217 5352
rect 54168 5312 54174 5324
rect 54205 5321 54217 5324
rect 54251 5321 54263 5355
rect 54205 5315 54263 5321
rect 48630 5256 48728 5284
rect 50424 5287 50482 5293
rect 48630 5253 48642 5256
rect 48584 5247 48642 5253
rect 50424 5253 50436 5287
rect 50470 5284 50482 5287
rect 51166 5284 51172 5296
rect 50470 5256 51172 5284
rect 50470 5253 50482 5256
rect 50424 5247 50482 5253
rect 51166 5244 51172 5256
rect 51224 5244 51230 5296
rect 1946 5176 1952 5228
rect 2004 5216 2010 5228
rect 2409 5219 2467 5225
rect 2409 5216 2421 5219
rect 2004 5188 2421 5216
rect 2004 5176 2010 5188
rect 2409 5185 2421 5188
rect 2455 5185 2467 5219
rect 2409 5179 2467 5185
rect 2676 5219 2734 5225
rect 2676 5185 2688 5219
rect 2722 5216 2734 5219
rect 5350 5216 5356 5228
rect 2722 5188 5356 5216
rect 2722 5185 2734 5188
rect 2676 5179 2734 5185
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 5810 5176 5816 5228
rect 5868 5216 5874 5228
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 5868 5188 6377 5216
rect 5868 5176 5874 5188
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 8938 5176 8944 5228
rect 8996 5216 9002 5228
rect 9217 5219 9275 5225
rect 9217 5216 9229 5219
rect 8996 5188 9229 5216
rect 8996 5176 9002 5188
rect 9217 5185 9229 5188
rect 9263 5216 9275 5219
rect 9766 5216 9772 5228
rect 9263 5188 9772 5216
rect 9263 5185 9275 5188
rect 9217 5179 9275 5185
rect 9766 5176 9772 5188
rect 9824 5176 9830 5228
rect 14452 5219 14510 5225
rect 14452 5185 14464 5219
rect 14498 5216 14510 5219
rect 14734 5216 14740 5228
rect 14498 5188 14740 5216
rect 14498 5185 14510 5188
rect 14452 5179 14510 5185
rect 14734 5176 14740 5188
rect 14792 5176 14798 5228
rect 18598 5176 18604 5228
rect 18656 5216 18662 5228
rect 23385 5219 23443 5225
rect 23385 5216 23397 5219
rect 18656 5188 23397 5216
rect 18656 5176 18662 5188
rect 23385 5185 23397 5188
rect 23431 5216 23443 5219
rect 28169 5219 28227 5225
rect 28169 5216 28181 5219
rect 23431 5188 28181 5216
rect 23431 5185 23443 5188
rect 23385 5179 23443 5185
rect 28169 5185 28181 5188
rect 28215 5185 28227 5219
rect 28169 5179 28227 5185
rect 32493 5219 32551 5225
rect 32493 5185 32505 5219
rect 32539 5216 32551 5219
rect 32582 5216 32588 5228
rect 32539 5188 32588 5216
rect 32539 5185 32551 5188
rect 32493 5179 32551 5185
rect 32582 5176 32588 5188
rect 32640 5176 32646 5228
rect 38004 5219 38062 5225
rect 38004 5185 38016 5219
rect 38050 5216 38062 5219
rect 39482 5216 39488 5228
rect 38050 5188 39488 5216
rect 38050 5185 38062 5188
rect 38004 5179 38062 5185
rect 39482 5176 39488 5188
rect 39540 5176 39546 5228
rect 43898 5176 43904 5228
rect 43956 5216 43962 5228
rect 43993 5219 44051 5225
rect 43993 5216 44005 5219
rect 43956 5188 44005 5216
rect 43956 5176 43962 5188
rect 43993 5185 44005 5188
rect 44039 5185 44051 5219
rect 43993 5179 44051 5185
rect 48317 5219 48375 5225
rect 48317 5185 48329 5219
rect 48363 5216 48375 5219
rect 48363 5188 50200 5216
rect 48363 5185 48375 5188
rect 48317 5179 48375 5185
rect 50172 5160 50200 5188
rect 52638 5176 52644 5228
rect 52696 5216 52702 5228
rect 52825 5219 52883 5225
rect 52825 5216 52837 5219
rect 52696 5188 52837 5216
rect 52696 5176 52702 5188
rect 52825 5185 52837 5188
rect 52871 5185 52883 5219
rect 52825 5179 52883 5185
rect 53092 5219 53150 5225
rect 53092 5185 53104 5219
rect 53138 5216 53150 5219
rect 54018 5216 54024 5228
rect 53138 5188 54024 5216
rect 53138 5185 53150 5188
rect 53092 5179 53150 5185
rect 54018 5176 54024 5188
rect 54076 5176 54082 5228
rect 3970 5108 3976 5160
rect 4028 5148 4034 5160
rect 4249 5151 4307 5157
rect 4249 5148 4261 5151
rect 4028 5120 4261 5148
rect 4028 5108 4034 5120
rect 4249 5117 4261 5120
rect 4295 5117 4307 5151
rect 13722 5148 13728 5160
rect 4249 5111 4307 5117
rect 13280 5120 13728 5148
rect 4062 4972 4068 5024
rect 4120 5012 4126 5024
rect 5629 5015 5687 5021
rect 5629 5012 5641 5015
rect 4120 4984 5641 5012
rect 4120 4972 4126 4984
rect 5629 4981 5641 4984
rect 5675 4981 5687 5015
rect 5629 4975 5687 4981
rect 7374 4972 7380 5024
rect 7432 5012 7438 5024
rect 7745 5015 7803 5021
rect 7745 5012 7757 5015
rect 7432 4984 7757 5012
rect 7432 4972 7438 4984
rect 7745 4981 7757 4984
rect 7791 4981 7803 5015
rect 7745 4975 7803 4981
rect 10686 4972 10692 5024
rect 10744 5012 10750 5024
rect 13280 5021 13308 5120
rect 13722 5108 13728 5120
rect 13780 5148 13786 5160
rect 14185 5151 14243 5157
rect 14185 5148 14197 5151
rect 13780 5120 14197 5148
rect 13780 5108 13786 5120
rect 14185 5117 14197 5120
rect 14231 5117 14243 5151
rect 14185 5111 14243 5117
rect 19889 5151 19947 5157
rect 19889 5117 19901 5151
rect 19935 5117 19947 5151
rect 19889 5111 19947 5117
rect 13265 5015 13323 5021
rect 13265 5012 13277 5015
rect 10744 4984 13277 5012
rect 10744 4972 10750 4984
rect 13265 4981 13277 4984
rect 13311 4981 13323 5015
rect 13265 4975 13323 4981
rect 13814 4972 13820 5024
rect 13872 5012 13878 5024
rect 15565 5015 15623 5021
rect 15565 5012 15577 5015
rect 13872 4984 15577 5012
rect 13872 4972 13878 4984
rect 15565 4981 15577 4984
rect 15611 4981 15623 5015
rect 19904 5012 19932 5111
rect 34606 5108 34612 5160
rect 34664 5148 34670 5160
rect 35161 5151 35219 5157
rect 35161 5148 35173 5151
rect 34664 5120 35173 5148
rect 34664 5108 34670 5120
rect 35161 5117 35173 5120
rect 35207 5117 35219 5151
rect 37734 5148 37740 5160
rect 37695 5120 37740 5148
rect 35161 5111 35219 5117
rect 37734 5108 37740 5120
rect 37792 5108 37798 5160
rect 41325 5151 41383 5157
rect 41325 5117 41337 5151
rect 41371 5148 41383 5151
rect 41690 5148 41696 5160
rect 41371 5120 41696 5148
rect 41371 5117 41383 5120
rect 41325 5111 41383 5117
rect 41690 5108 41696 5120
rect 41748 5108 41754 5160
rect 50154 5148 50160 5160
rect 50115 5120 50160 5148
rect 50154 5108 50160 5120
rect 50212 5108 50218 5160
rect 22002 5080 22008 5092
rect 20824 5052 22008 5080
rect 20824 5012 20852 5052
rect 22002 5040 22008 5052
rect 22060 5040 22066 5092
rect 19904 4984 20852 5012
rect 21269 5015 21327 5021
rect 15565 4975 15623 4981
rect 21269 4981 21281 5015
rect 21315 5012 21327 5015
rect 22738 5012 22744 5024
rect 21315 4984 22744 5012
rect 21315 4981 21327 4984
rect 21269 4975 21327 4981
rect 22738 4972 22744 4984
rect 22796 4972 22802 5024
rect 24026 4972 24032 5024
rect 24084 5012 24090 5024
rect 24670 5012 24676 5024
rect 24084 4984 24676 5012
rect 24084 4972 24090 4984
rect 24670 4972 24676 4984
rect 24728 4972 24734 5024
rect 33870 5012 33876 5024
rect 33831 4984 33876 5012
rect 33870 4972 33876 4984
rect 33928 4972 33934 5024
rect 36538 5012 36544 5024
rect 36499 4984 36544 5012
rect 36538 4972 36544 4984
rect 36596 4972 36602 5024
rect 39117 5015 39175 5021
rect 39117 4981 39129 5015
rect 39163 5012 39175 5015
rect 39942 5012 39948 5024
rect 39163 4984 39948 5012
rect 39163 4981 39175 4984
rect 39117 4975 39175 4981
rect 39942 4972 39948 4984
rect 40000 4972 40006 5024
rect 49697 5015 49755 5021
rect 49697 4981 49709 5015
rect 49743 5012 49755 5015
rect 50430 5012 50436 5024
rect 49743 4984 50436 5012
rect 49743 4981 49755 4984
rect 49697 4975 49755 4981
rect 50430 4972 50436 4984
rect 50488 4972 50494 5024
rect 1104 4922 59340 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 59340 4922
rect 1104 4848 59340 4870
rect 15470 4808 15476 4820
rect 15431 4780 15476 4808
rect 15470 4768 15476 4780
rect 15528 4768 15534 4820
rect 16298 4808 16304 4820
rect 15948 4780 16304 4808
rect 9766 4672 9772 4684
rect 9727 4644 9772 4672
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 10778 4632 10784 4684
rect 10836 4672 10842 4684
rect 15948 4681 15976 4780
rect 16298 4768 16304 4780
rect 16356 4768 16362 4820
rect 21453 4811 21511 4817
rect 21453 4777 21465 4811
rect 21499 4808 21511 4811
rect 22094 4808 22100 4820
rect 21499 4780 22100 4808
rect 21499 4777 21511 4780
rect 21453 4771 21511 4777
rect 22094 4768 22100 4780
rect 22152 4768 22158 4820
rect 23290 4808 23296 4820
rect 23251 4780 23296 4808
rect 23290 4768 23296 4780
rect 23348 4768 23354 4820
rect 36722 4808 36728 4820
rect 36683 4780 36728 4808
rect 36722 4768 36728 4780
rect 36780 4768 36786 4820
rect 41230 4808 41236 4820
rect 41191 4780 41236 4808
rect 41230 4768 41236 4780
rect 41288 4768 41294 4820
rect 47394 4768 47400 4820
rect 47452 4808 47458 4820
rect 48961 4811 49019 4817
rect 48961 4808 48973 4811
rect 47452 4780 48973 4808
rect 47452 4768 47458 4780
rect 48961 4777 48973 4780
rect 49007 4777 49019 4811
rect 48961 4771 49019 4777
rect 11609 4675 11667 4681
rect 11609 4672 11621 4675
rect 10836 4644 11621 4672
rect 10836 4632 10842 4644
rect 11609 4641 11621 4644
rect 11655 4641 11667 4675
rect 11609 4635 11667 4641
rect 15933 4675 15991 4681
rect 15933 4641 15945 4675
rect 15979 4641 15991 4675
rect 26970 4672 26976 4684
rect 26931 4644 26976 4672
rect 15933 4635 15991 4641
rect 26970 4632 26976 4644
rect 27028 4632 27034 4684
rect 29178 4632 29184 4684
rect 29236 4672 29242 4684
rect 30009 4675 30067 4681
rect 30009 4672 30021 4675
rect 29236 4644 30021 4672
rect 29236 4632 29242 4644
rect 30009 4641 30021 4644
rect 30055 4641 30067 4675
rect 30009 4635 30067 4641
rect 4062 4613 4068 4616
rect 3789 4607 3847 4613
rect 3789 4573 3801 4607
rect 3835 4573 3847 4607
rect 4056 4604 4068 4613
rect 4023 4576 4068 4604
rect 3789 4567 3847 4573
rect 4056 4567 4068 4576
rect 3804 4536 3832 4567
rect 4062 4564 4068 4567
rect 4120 4564 4126 4616
rect 5629 4607 5687 4613
rect 5629 4604 5641 4607
rect 4172 4576 5641 4604
rect 4172 4536 4200 4576
rect 5629 4573 5641 4576
rect 5675 4604 5687 4607
rect 5718 4604 5724 4616
rect 5675 4576 5724 4604
rect 5675 4573 5687 4576
rect 5629 4567 5687 4573
rect 5718 4564 5724 4576
rect 5776 4564 5782 4616
rect 10036 4607 10094 4613
rect 10036 4573 10048 4607
rect 10082 4604 10094 4607
rect 11146 4604 11152 4616
rect 10082 4576 11152 4604
rect 10082 4573 10094 4576
rect 10036 4567 10094 4573
rect 11146 4564 11152 4576
rect 11204 4564 11210 4616
rect 13354 4564 13360 4616
rect 13412 4604 13418 4616
rect 14093 4607 14151 4613
rect 14093 4604 14105 4607
rect 13412 4576 14105 4604
rect 13412 4564 13418 4576
rect 14093 4573 14105 4576
rect 14139 4573 14151 4607
rect 14093 4567 14151 4573
rect 19426 4564 19432 4616
rect 19484 4604 19490 4616
rect 20073 4607 20131 4613
rect 20073 4604 20085 4607
rect 19484 4576 20085 4604
rect 19484 4564 19490 4576
rect 20073 4573 20085 4576
rect 20119 4604 20131 4607
rect 20622 4604 20628 4616
rect 20119 4576 20628 4604
rect 20119 4573 20131 4576
rect 20073 4567 20131 4573
rect 20622 4564 20628 4576
rect 20680 4564 20686 4616
rect 21913 4607 21971 4613
rect 21913 4573 21925 4607
rect 21959 4604 21971 4607
rect 22002 4604 22008 4616
rect 21959 4576 22008 4604
rect 21959 4573 21971 4576
rect 21913 4567 21971 4573
rect 22002 4564 22008 4576
rect 22060 4564 22066 4616
rect 25133 4607 25191 4613
rect 25133 4573 25145 4607
rect 25179 4604 25191 4607
rect 26988 4604 27016 4632
rect 27246 4613 27252 4616
rect 27240 4604 27252 4613
rect 25179 4576 27016 4604
rect 27207 4576 27252 4604
rect 25179 4573 25191 4576
rect 25133 4567 25191 4573
rect 27240 4567 27252 4576
rect 27246 4564 27252 4567
rect 27304 4564 27310 4616
rect 30276 4607 30334 4613
rect 30276 4573 30288 4607
rect 30322 4604 30334 4607
rect 31110 4604 31116 4616
rect 30322 4576 31116 4604
rect 30322 4573 30334 4576
rect 30276 4567 30334 4573
rect 31110 4564 31116 4576
rect 31168 4564 31174 4616
rect 32582 4564 32588 4616
rect 32640 4604 32646 4616
rect 32769 4607 32827 4613
rect 32769 4604 32781 4607
rect 32640 4576 32781 4604
rect 32640 4564 32646 4576
rect 32769 4573 32781 4576
rect 32815 4573 32827 4607
rect 32769 4567 32827 4573
rect 33036 4607 33094 4613
rect 33036 4573 33048 4607
rect 33082 4604 33094 4607
rect 33870 4604 33876 4616
rect 33082 4576 33876 4604
rect 33082 4573 33094 4576
rect 33036 4567 33094 4573
rect 33870 4564 33876 4576
rect 33928 4564 33934 4616
rect 34606 4564 34612 4616
rect 34664 4604 34670 4616
rect 35345 4607 35403 4613
rect 35345 4604 35357 4607
rect 34664 4576 35357 4604
rect 34664 4564 34670 4576
rect 35345 4573 35357 4576
rect 35391 4573 35403 4607
rect 35345 4567 35403 4573
rect 35612 4607 35670 4613
rect 35612 4573 35624 4607
rect 35658 4604 35670 4607
rect 36538 4604 36544 4616
rect 35658 4576 36544 4604
rect 35658 4573 35670 4576
rect 35612 4567 35670 4573
rect 3804 4508 4200 4536
rect 5534 4496 5540 4548
rect 5592 4536 5598 4548
rect 5874 4539 5932 4545
rect 5874 4536 5886 4539
rect 5592 4508 5886 4536
rect 5592 4496 5598 4508
rect 5874 4505 5886 4508
rect 5920 4505 5932 4539
rect 11854 4539 11912 4545
rect 11854 4536 11866 4539
rect 5874 4499 5932 4505
rect 11164 4508 11866 4536
rect 5166 4468 5172 4480
rect 5127 4440 5172 4468
rect 5166 4428 5172 4440
rect 5224 4428 5230 4480
rect 5994 4428 6000 4480
rect 6052 4468 6058 4480
rect 11164 4477 11192 4508
rect 11854 4505 11866 4508
rect 11900 4505 11912 4539
rect 11854 4499 11912 4505
rect 14360 4539 14418 4545
rect 14360 4505 14372 4539
rect 14406 4536 14418 4539
rect 15470 4536 15476 4548
rect 14406 4508 15476 4536
rect 14406 4505 14418 4508
rect 14360 4499 14418 4505
rect 15470 4496 15476 4508
rect 15528 4496 15534 4548
rect 16200 4539 16258 4545
rect 16200 4505 16212 4539
rect 16246 4536 16258 4539
rect 17126 4536 17132 4548
rect 16246 4508 17132 4536
rect 16246 4505 16258 4508
rect 16200 4499 16258 4505
rect 17126 4496 17132 4508
rect 17184 4496 17190 4548
rect 20340 4539 20398 4545
rect 20340 4505 20352 4539
rect 20386 4536 20398 4539
rect 21818 4536 21824 4548
rect 20386 4508 21824 4536
rect 20386 4505 20398 4508
rect 20340 4499 20398 4505
rect 21818 4496 21824 4508
rect 21876 4496 21882 4548
rect 22180 4539 22238 4545
rect 22180 4505 22192 4539
rect 22226 4536 22238 4539
rect 23198 4536 23204 4548
rect 22226 4508 23204 4536
rect 22226 4505 22238 4508
rect 22180 4499 22238 4505
rect 23198 4496 23204 4508
rect 23256 4496 23262 4548
rect 25400 4539 25458 4545
rect 25400 4505 25412 4539
rect 25446 4536 25458 4539
rect 35360 4536 35388 4567
rect 36538 4564 36544 4576
rect 36596 4564 36602 4616
rect 37185 4607 37243 4613
rect 37185 4573 37197 4607
rect 37231 4573 37243 4607
rect 39850 4604 39856 4616
rect 39763 4576 39856 4604
rect 37185 4567 37243 4573
rect 35802 4536 35808 4548
rect 25446 4508 28396 4536
rect 35360 4508 35808 4536
rect 25446 4505 25458 4508
rect 25400 4499 25458 4505
rect 7009 4471 7067 4477
rect 7009 4468 7021 4471
rect 6052 4440 7021 4468
rect 6052 4428 6058 4440
rect 7009 4437 7021 4440
rect 7055 4437 7067 4471
rect 7009 4431 7067 4437
rect 11149 4471 11207 4477
rect 11149 4437 11161 4471
rect 11195 4437 11207 4471
rect 11149 4431 11207 4437
rect 11238 4428 11244 4480
rect 11296 4468 11302 4480
rect 12989 4471 13047 4477
rect 12989 4468 13001 4471
rect 11296 4440 13001 4468
rect 11296 4428 11302 4440
rect 12989 4437 13001 4440
rect 13035 4437 13047 4471
rect 17310 4468 17316 4480
rect 17271 4440 17316 4468
rect 12989 4431 13047 4437
rect 17310 4428 17316 4440
rect 17368 4428 17374 4480
rect 26510 4468 26516 4480
rect 26471 4440 26516 4468
rect 26510 4428 26516 4440
rect 26568 4428 26574 4480
rect 28368 4477 28396 4508
rect 35802 4496 35808 4508
rect 35860 4536 35866 4548
rect 37200 4536 37228 4567
rect 35860 4508 37228 4536
rect 37452 4539 37510 4545
rect 35860 4496 35866 4508
rect 37452 4505 37464 4539
rect 37498 4536 37510 4539
rect 38838 4536 38844 4548
rect 37498 4508 38844 4536
rect 37498 4505 37510 4508
rect 37452 4499 37510 4505
rect 38838 4496 38844 4508
rect 38896 4496 38902 4548
rect 39776 4536 39804 4576
rect 39850 4564 39856 4576
rect 39908 4564 39914 4616
rect 39942 4564 39948 4616
rect 40000 4604 40006 4616
rect 40109 4607 40167 4613
rect 40109 4604 40121 4607
rect 40000 4576 40121 4604
rect 40000 4564 40006 4576
rect 40109 4573 40121 4576
rect 40155 4573 40167 4607
rect 41690 4604 41696 4616
rect 40109 4567 40167 4573
rect 40236 4576 41696 4604
rect 40236 4536 40264 4576
rect 41690 4564 41696 4576
rect 41748 4604 41754 4616
rect 42426 4604 42432 4616
rect 41748 4576 42432 4604
rect 41748 4564 41754 4576
rect 42426 4564 42432 4576
rect 42484 4564 42490 4616
rect 47581 4607 47639 4613
rect 47581 4573 47593 4607
rect 47627 4573 47639 4607
rect 47581 4567 47639 4573
rect 39776 4508 40264 4536
rect 41506 4496 41512 4548
rect 41564 4536 41570 4548
rect 41938 4539 41996 4545
rect 41938 4536 41950 4539
rect 41564 4508 41950 4536
rect 41564 4496 41570 4508
rect 41938 4505 41950 4508
rect 41984 4505 41996 4539
rect 47596 4536 47624 4567
rect 47670 4564 47676 4616
rect 47728 4604 47734 4616
rect 47837 4607 47895 4613
rect 47837 4604 47849 4607
rect 47728 4576 47849 4604
rect 47728 4564 47734 4576
rect 47837 4573 47849 4576
rect 47883 4573 47895 4607
rect 50154 4604 50160 4616
rect 50115 4576 50160 4604
rect 47837 4567 47895 4573
rect 50154 4564 50160 4576
rect 50212 4564 50218 4616
rect 50430 4613 50436 4616
rect 50424 4604 50436 4613
rect 50391 4576 50436 4604
rect 50424 4567 50436 4576
rect 50430 4564 50436 4567
rect 50488 4564 50494 4616
rect 51997 4607 52055 4613
rect 51997 4573 52009 4607
rect 52043 4604 52055 4607
rect 52730 4604 52736 4616
rect 52043 4576 52736 4604
rect 52043 4573 52055 4576
rect 51997 4567 52055 4573
rect 52730 4564 52736 4576
rect 52788 4564 52794 4616
rect 48222 4536 48228 4548
rect 47596 4508 48228 4536
rect 41938 4499 41996 4505
rect 48222 4496 48228 4508
rect 48280 4496 48286 4548
rect 52264 4539 52322 4545
rect 52264 4505 52276 4539
rect 52310 4536 52322 4539
rect 53558 4536 53564 4548
rect 52310 4508 53564 4536
rect 52310 4505 52322 4508
rect 52264 4499 52322 4505
rect 53558 4496 53564 4508
rect 53616 4496 53622 4548
rect 28353 4471 28411 4477
rect 28353 4437 28365 4471
rect 28399 4437 28411 4471
rect 31386 4468 31392 4480
rect 31347 4440 31392 4468
rect 28353 4431 28411 4437
rect 31386 4428 31392 4440
rect 31444 4428 31450 4480
rect 34146 4468 34152 4480
rect 34107 4440 34152 4468
rect 34146 4428 34152 4440
rect 34204 4428 34210 4480
rect 38562 4468 38568 4480
rect 38523 4440 38568 4468
rect 38562 4428 38568 4440
rect 38620 4428 38626 4480
rect 43070 4468 43076 4480
rect 43031 4440 43076 4468
rect 43070 4428 43076 4440
rect 43128 4428 43134 4480
rect 51534 4468 51540 4480
rect 51495 4440 51540 4468
rect 51534 4428 51540 4440
rect 51592 4428 51598 4480
rect 53374 4468 53380 4480
rect 53335 4440 53380 4468
rect 53374 4428 53380 4440
rect 53432 4428 53438 4480
rect 1104 4378 59340 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 59340 4378
rect 1104 4304 59340 4326
rect 3970 4224 3976 4276
rect 4028 4224 4034 4276
rect 14734 4264 14740 4276
rect 14695 4236 14740 4264
rect 14734 4224 14740 4236
rect 14792 4224 14798 4276
rect 23198 4264 23204 4276
rect 23159 4236 23204 4264
rect 23198 4224 23204 4236
rect 23256 4224 23262 4276
rect 3988 4196 4016 4224
rect 18598 4196 18604 4208
rect 3712 4168 4016 4196
rect 18559 4168 18604 4196
rect 3712 4137 3740 4168
rect 18598 4156 18604 4168
rect 18656 4156 18662 4208
rect 22002 4196 22008 4208
rect 21836 4168 22008 4196
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4097 3755 4131
rect 3697 4091 3755 4097
rect 3964 4131 4022 4137
rect 3964 4097 3976 4131
rect 4010 4128 4022 4131
rect 5166 4128 5172 4140
rect 4010 4100 5172 4128
rect 4010 4097 4022 4100
rect 3964 4091 4022 4097
rect 5166 4088 5172 4100
rect 5224 4088 5230 4140
rect 5718 4088 5724 4140
rect 5776 4128 5782 4140
rect 6365 4131 6423 4137
rect 6365 4128 6377 4131
rect 5776 4100 6377 4128
rect 5776 4088 5782 4100
rect 6365 4097 6377 4100
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 6632 4131 6690 4137
rect 6632 4097 6644 4131
rect 6678 4128 6690 4131
rect 7374 4128 7380 4140
rect 6678 4100 7380 4128
rect 6678 4097 6690 4100
rect 6632 4091 6690 4097
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 10778 4088 10784 4140
rect 10836 4128 10842 4140
rect 11790 4137 11796 4140
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 10836 4100 11529 4128
rect 10836 4088 10842 4100
rect 11517 4097 11529 4100
rect 11563 4097 11575 4131
rect 11517 4091 11575 4097
rect 11784 4091 11796 4137
rect 11848 4128 11854 4140
rect 11848 4100 11884 4128
rect 11790 4088 11796 4091
rect 11848 4088 11854 4100
rect 13078 4088 13084 4140
rect 13136 4128 13142 4140
rect 13613 4131 13671 4137
rect 13613 4128 13625 4131
rect 13136 4100 13625 4128
rect 13136 4088 13142 4100
rect 13613 4097 13625 4100
rect 13659 4097 13671 4131
rect 13613 4091 13671 4097
rect 16298 4088 16304 4140
rect 16356 4128 16362 4140
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 16356 4100 16681 4128
rect 16356 4088 16362 4100
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 16758 4088 16764 4140
rect 16816 4128 16822 4140
rect 21836 4137 21864 4168
rect 22002 4156 22008 4168
rect 22060 4156 22066 4208
rect 26510 4156 26516 4208
rect 26568 4196 26574 4208
rect 27218 4199 27276 4205
rect 27218 4196 27230 4199
rect 26568 4168 27230 4196
rect 26568 4156 26574 4168
rect 27218 4165 27230 4168
rect 27264 4165 27276 4199
rect 37734 4196 37740 4208
rect 27218 4159 27276 4165
rect 37292 4168 37740 4196
rect 37292 4140 37320 4168
rect 37734 4156 37740 4168
rect 37792 4196 37798 4208
rect 39850 4196 39856 4208
rect 37792 4168 39856 4196
rect 37792 4156 37798 4168
rect 22094 4137 22100 4140
rect 16925 4131 16983 4137
rect 16925 4128 16937 4131
rect 16816 4100 16937 4128
rect 16816 4088 16822 4100
rect 16925 4097 16937 4100
rect 16971 4097 16983 4131
rect 16925 4091 16983 4097
rect 21821 4131 21879 4137
rect 21821 4097 21833 4131
rect 21867 4097 21879 4131
rect 22088 4128 22100 4137
rect 22055 4100 22100 4128
rect 21821 4091 21879 4097
rect 22088 4091 22100 4100
rect 22094 4088 22100 4091
rect 22152 4088 22158 4140
rect 24296 4131 24354 4137
rect 24296 4097 24308 4131
rect 24342 4128 24354 4131
rect 25682 4128 25688 4140
rect 24342 4100 25688 4128
rect 24342 4097 24354 4100
rect 24296 4091 24354 4097
rect 25682 4088 25688 4100
rect 25740 4088 25746 4140
rect 26970 4128 26976 4140
rect 26931 4100 26976 4128
rect 26970 4088 26976 4100
rect 27028 4088 27034 4140
rect 30000 4131 30058 4137
rect 30000 4097 30012 4131
rect 30046 4128 30058 4131
rect 31386 4128 31392 4140
rect 30046 4100 31392 4128
rect 30046 4097 30058 4100
rect 30000 4091 30058 4097
rect 31386 4088 31392 4100
rect 31444 4088 31450 4140
rect 33036 4131 33094 4137
rect 33036 4097 33048 4131
rect 33082 4128 33094 4131
rect 34146 4128 34152 4140
rect 33082 4100 34152 4128
rect 33082 4097 33094 4100
rect 33036 4091 33094 4097
rect 34146 4088 34152 4100
rect 34204 4088 34210 4140
rect 34865 4131 34923 4137
rect 34865 4128 34877 4131
rect 34532 4100 34877 4128
rect 13354 4060 13360 4072
rect 13315 4032 13360 4060
rect 13354 4020 13360 4032
rect 13412 4020 13418 4072
rect 20349 4063 20407 4069
rect 20349 4029 20361 4063
rect 20395 4060 20407 4063
rect 20622 4060 20628 4072
rect 20395 4032 20628 4060
rect 20395 4029 20407 4032
rect 20349 4023 20407 4029
rect 20622 4020 20628 4032
rect 20680 4020 20686 4072
rect 24026 4060 24032 4072
rect 23987 4032 24032 4060
rect 24026 4020 24032 4032
rect 24084 4020 24090 4072
rect 29733 4063 29791 4069
rect 29733 4029 29745 4063
rect 29779 4029 29791 4063
rect 32582 4060 32588 4072
rect 29733 4023 29791 4029
rect 30944 4032 32588 4060
rect 5077 3995 5135 4001
rect 5077 3961 5089 3995
rect 5123 3992 5135 3995
rect 5534 3992 5540 4004
rect 5123 3964 5540 3992
rect 5123 3961 5135 3964
rect 5077 3955 5135 3961
rect 5534 3952 5540 3964
rect 5592 3952 5598 4004
rect 7742 3992 7748 4004
rect 7703 3964 7748 3992
rect 7742 3952 7748 3964
rect 7800 3952 7806 4004
rect 12894 3924 12900 3936
rect 12855 3896 12900 3924
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 18046 3924 18052 3936
rect 18007 3896 18052 3924
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 25406 3924 25412 3936
rect 25367 3896 25412 3924
rect 25406 3884 25412 3896
rect 25464 3884 25470 3936
rect 28350 3924 28356 3936
rect 28311 3896 28356 3924
rect 28350 3884 28356 3896
rect 28408 3884 28414 3936
rect 29748 3924 29776 4023
rect 30944 3924 30972 4032
rect 32582 4020 32588 4032
rect 32640 4060 32646 4072
rect 32769 4063 32827 4069
rect 32769 4060 32781 4063
rect 32640 4032 32781 4060
rect 32640 4020 32646 4032
rect 32769 4029 32781 4032
rect 32815 4029 32827 4063
rect 34532 4060 34560 4100
rect 34865 4097 34877 4100
rect 34911 4097 34923 4131
rect 37274 4128 37280 4140
rect 37187 4100 37280 4128
rect 34865 4091 34923 4097
rect 37274 4088 37280 4100
rect 37332 4088 37338 4140
rect 37544 4131 37602 4137
rect 37544 4097 37556 4131
rect 37590 4128 37602 4131
rect 38746 4128 38752 4140
rect 37590 4100 38752 4128
rect 37590 4097 37602 4100
rect 37544 4091 37602 4097
rect 38746 4088 38752 4100
rect 38804 4088 38810 4140
rect 39132 4137 39160 4168
rect 39850 4156 39856 4168
rect 39908 4156 39914 4208
rect 53000 4199 53058 4205
rect 53000 4165 53012 4199
rect 53046 4196 53058 4199
rect 53374 4196 53380 4208
rect 53046 4168 53380 4196
rect 53046 4165 53058 4168
rect 53000 4159 53058 4165
rect 53374 4156 53380 4168
rect 53432 4156 53438 4208
rect 39117 4131 39175 4137
rect 39117 4097 39129 4131
rect 39163 4097 39175 4131
rect 39117 4091 39175 4097
rect 39384 4131 39442 4137
rect 39384 4097 39396 4131
rect 39430 4128 39442 4131
rect 40402 4128 40408 4140
rect 39430 4100 40408 4128
rect 39430 4097 39442 4100
rect 39384 4091 39442 4097
rect 40402 4088 40408 4100
rect 40460 4088 40466 4140
rect 44266 4137 44272 4140
rect 44260 4128 44272 4137
rect 44227 4100 44272 4128
rect 44260 4091 44272 4100
rect 44266 4088 44272 4091
rect 44324 4088 44330 4140
rect 47026 4088 47032 4140
rect 47084 4128 47090 4140
rect 47837 4131 47895 4137
rect 47837 4128 47849 4131
rect 47084 4100 47849 4128
rect 47084 4088 47090 4100
rect 47837 4097 47849 4100
rect 47883 4097 47895 4131
rect 47837 4091 47895 4097
rect 49881 4131 49939 4137
rect 49881 4097 49893 4131
rect 49927 4128 49939 4131
rect 49970 4128 49976 4140
rect 49927 4100 49976 4128
rect 49927 4097 49939 4100
rect 49881 4091 49939 4097
rect 49970 4088 49976 4100
rect 50028 4088 50034 4140
rect 50148 4131 50206 4137
rect 50148 4097 50160 4131
rect 50194 4128 50206 4131
rect 51534 4128 51540 4140
rect 50194 4100 51540 4128
rect 50194 4097 50206 4100
rect 50148 4091 50206 4097
rect 51534 4088 51540 4100
rect 51592 4088 51598 4140
rect 52730 4128 52736 4140
rect 52691 4100 52736 4128
rect 52730 4088 52736 4100
rect 52788 4088 52794 4140
rect 32769 4023 32827 4029
rect 34164 4032 34560 4060
rect 34164 4001 34192 4032
rect 34606 4020 34612 4072
rect 34664 4060 34670 4072
rect 34664 4032 34709 4060
rect 34664 4020 34670 4032
rect 42426 4020 42432 4072
rect 42484 4060 42490 4072
rect 43993 4063 44051 4069
rect 43993 4060 44005 4063
rect 42484 4032 44005 4060
rect 42484 4020 42490 4032
rect 43993 4029 44005 4032
rect 44039 4029 44051 4063
rect 43993 4023 44051 4029
rect 46934 4020 46940 4072
rect 46992 4060 46998 4072
rect 47581 4063 47639 4069
rect 47581 4060 47593 4063
rect 46992 4032 47593 4060
rect 46992 4020 46998 4032
rect 47581 4029 47593 4032
rect 47627 4029 47639 4063
rect 47581 4023 47639 4029
rect 34149 3995 34207 4001
rect 34149 3961 34161 3995
rect 34195 3961 34207 3995
rect 35986 3992 35992 4004
rect 35947 3964 35992 3992
rect 34149 3955 34207 3961
rect 35986 3952 35992 3964
rect 36044 3952 36050 4004
rect 45278 3952 45284 4004
rect 45336 3992 45342 4004
rect 45373 3995 45431 4001
rect 45373 3992 45385 3995
rect 45336 3964 45385 3992
rect 45336 3952 45342 3964
rect 45373 3961 45385 3964
rect 45419 3961 45431 3995
rect 45373 3955 45431 3961
rect 31110 3924 31116 3936
rect 29748 3896 30972 3924
rect 31071 3896 31116 3924
rect 31110 3884 31116 3896
rect 31168 3884 31174 3936
rect 38654 3924 38660 3936
rect 38615 3896 38660 3924
rect 38654 3884 38660 3896
rect 38712 3884 38718 3936
rect 40494 3924 40500 3936
rect 40455 3896 40500 3924
rect 40494 3884 40500 3896
rect 40552 3884 40558 3936
rect 48958 3924 48964 3936
rect 48919 3896 48964 3924
rect 48958 3884 48964 3896
rect 49016 3884 49022 3936
rect 50614 3884 50620 3936
rect 50672 3924 50678 3936
rect 51261 3927 51319 3933
rect 51261 3924 51273 3927
rect 50672 3896 51273 3924
rect 50672 3884 50678 3896
rect 51261 3893 51273 3896
rect 51307 3893 51319 3927
rect 54110 3924 54116 3936
rect 54071 3896 54116 3924
rect 51261 3887 51319 3893
rect 54110 3884 54116 3896
rect 54168 3884 54174 3936
rect 1104 3834 59340 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 59340 3834
rect 1104 3760 59340 3782
rect 5718 3720 5724 3732
rect 4632 3692 5724 3720
rect 4632 3593 4660 3692
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 5997 3723 6055 3729
rect 5997 3689 6009 3723
rect 6043 3720 6055 3723
rect 6086 3720 6092 3732
rect 6043 3692 6092 3720
rect 6043 3689 6055 3692
rect 5997 3683 6055 3689
rect 6086 3680 6092 3692
rect 6144 3680 6150 3732
rect 10778 3720 10784 3732
rect 10428 3692 10784 3720
rect 10428 3593 10456 3692
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 11790 3720 11796 3732
rect 11751 3692 11796 3720
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 15470 3720 15476 3732
rect 15431 3692 15476 3720
rect 15470 3680 15476 3692
rect 15528 3680 15534 3732
rect 16298 3720 16304 3732
rect 15948 3692 16304 3720
rect 4617 3587 4675 3593
rect 4617 3553 4629 3587
rect 4663 3553 4675 3587
rect 4617 3547 4675 3553
rect 10413 3587 10471 3593
rect 10413 3553 10425 3587
rect 10459 3553 10471 3587
rect 10413 3547 10471 3553
rect 13354 3544 13360 3596
rect 13412 3584 13418 3596
rect 15948 3593 15976 3692
rect 16298 3680 16304 3692
rect 16356 3680 16362 3732
rect 17126 3680 17132 3732
rect 17184 3720 17190 3732
rect 17313 3723 17371 3729
rect 17313 3720 17325 3723
rect 17184 3692 17325 3720
rect 17184 3680 17190 3692
rect 17313 3689 17325 3692
rect 17359 3689 17371 3723
rect 17313 3683 17371 3689
rect 21818 3680 21824 3732
rect 21876 3720 21882 3732
rect 22465 3723 22523 3729
rect 22465 3720 22477 3723
rect 21876 3692 22477 3720
rect 21876 3680 21882 3692
rect 22465 3689 22477 3692
rect 22511 3689 22523 3723
rect 26970 3720 26976 3732
rect 22465 3683 22523 3689
rect 26712 3692 26976 3720
rect 26712 3593 26740 3692
rect 26970 3680 26976 3692
rect 27028 3680 27034 3732
rect 31018 3720 31024 3732
rect 30979 3692 31024 3720
rect 31018 3680 31024 3692
rect 31076 3680 31082 3732
rect 39482 3680 39488 3732
rect 39540 3720 39546 3732
rect 41233 3723 41291 3729
rect 41233 3720 41245 3723
rect 39540 3692 41245 3720
rect 39540 3680 39546 3692
rect 41233 3689 41245 3692
rect 41279 3689 41291 3723
rect 42794 3720 42800 3732
rect 41233 3683 41291 3689
rect 42444 3692 42800 3720
rect 14093 3587 14151 3593
rect 14093 3584 14105 3587
rect 13412 3556 14105 3584
rect 13412 3544 13418 3556
rect 14093 3553 14105 3556
rect 14139 3553 14151 3587
rect 14093 3547 14151 3553
rect 15933 3587 15991 3593
rect 15933 3553 15945 3587
rect 15979 3553 15991 3587
rect 15933 3547 15991 3553
rect 26697 3587 26755 3593
rect 26697 3553 26709 3587
rect 26743 3553 26755 3587
rect 32582 3584 32588 3596
rect 32543 3556 32588 3584
rect 26697 3547 26755 3553
rect 4884 3519 4942 3525
rect 4884 3485 4896 3519
rect 4930 3516 4942 3519
rect 5994 3516 6000 3528
rect 4930 3488 6000 3516
rect 4930 3485 4942 3488
rect 4884 3479 4942 3485
rect 5994 3476 6000 3488
rect 6052 3476 6058 3528
rect 10680 3519 10738 3525
rect 10680 3485 10692 3519
rect 10726 3516 10738 3519
rect 11238 3516 11244 3528
rect 10726 3488 11244 3516
rect 10726 3485 10738 3488
rect 10680 3479 10738 3485
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 16200 3519 16258 3525
rect 16200 3485 16212 3519
rect 16246 3516 16258 3519
rect 18046 3516 18052 3528
rect 16246 3488 18052 3516
rect 16246 3485 16258 3488
rect 16200 3479 16258 3485
rect 18046 3476 18052 3488
rect 18104 3476 18110 3528
rect 19245 3519 19303 3525
rect 19245 3485 19257 3519
rect 19291 3516 19303 3519
rect 19334 3516 19340 3528
rect 19291 3488 19340 3516
rect 19291 3485 19303 3488
rect 19245 3479 19303 3485
rect 19334 3476 19340 3488
rect 19392 3516 19398 3528
rect 20622 3516 20628 3528
rect 19392 3488 20628 3516
rect 19392 3476 19398 3488
rect 20622 3476 20628 3488
rect 20680 3516 20686 3528
rect 21085 3519 21143 3525
rect 21085 3516 21097 3519
rect 20680 3488 21097 3516
rect 20680 3476 20686 3488
rect 21085 3485 21097 3488
rect 21131 3485 21143 3519
rect 21085 3479 21143 3485
rect 24857 3519 24915 3525
rect 24857 3485 24869 3519
rect 24903 3516 24915 3519
rect 26712 3516 26740 3547
rect 32582 3544 32588 3556
rect 32640 3544 32646 3596
rect 34606 3544 34612 3596
rect 34664 3584 34670 3596
rect 34701 3587 34759 3593
rect 34701 3584 34713 3587
rect 34664 3556 34713 3584
rect 34664 3544 34670 3556
rect 34701 3553 34713 3556
rect 34747 3553 34759 3587
rect 39850 3584 39856 3596
rect 39811 3556 39856 3584
rect 34701 3547 34759 3553
rect 24903 3488 26740 3516
rect 26964 3519 27022 3525
rect 24903 3485 24915 3488
rect 24857 3479 24915 3485
rect 26964 3485 26976 3519
rect 27010 3516 27022 3519
rect 28350 3516 28356 3528
rect 27010 3488 28356 3516
rect 27010 3485 27022 3488
rect 26964 3479 27022 3485
rect 28350 3476 28356 3488
rect 28408 3476 28414 3528
rect 29641 3519 29699 3525
rect 29641 3485 29653 3519
rect 29687 3516 29699 3519
rect 29730 3516 29736 3528
rect 29687 3488 29736 3516
rect 29687 3485 29699 3488
rect 29641 3479 29699 3485
rect 29730 3476 29736 3488
rect 29788 3476 29794 3528
rect 29908 3519 29966 3525
rect 29908 3485 29920 3519
rect 29954 3516 29966 3519
rect 31110 3516 31116 3528
rect 29954 3488 31116 3516
rect 29954 3485 29966 3488
rect 29908 3479 29966 3485
rect 31110 3476 31116 3488
rect 31168 3476 31174 3528
rect 34716 3516 34744 3547
rect 39850 3544 39856 3556
rect 39908 3544 39914 3596
rect 42444 3593 42472 3692
rect 42794 3680 42800 3692
rect 42852 3680 42858 3732
rect 43806 3720 43812 3732
rect 43767 3692 43812 3720
rect 43806 3680 43812 3692
rect 43864 3680 43870 3732
rect 49602 3720 49608 3732
rect 49563 3692 49608 3720
rect 49602 3680 49608 3692
rect 49660 3680 49666 3732
rect 53558 3720 53564 3732
rect 53519 3692 53564 3720
rect 53558 3680 53564 3692
rect 53616 3680 53622 3732
rect 42429 3587 42487 3593
rect 42429 3553 42441 3587
rect 42475 3553 42487 3587
rect 42429 3547 42487 3553
rect 36541 3519 36599 3525
rect 36541 3516 36553 3519
rect 34716 3488 36553 3516
rect 36541 3485 36553 3488
rect 36587 3485 36599 3519
rect 36541 3479 36599 3485
rect 40120 3519 40178 3525
rect 40120 3485 40132 3519
rect 40166 3516 40178 3519
rect 40494 3516 40500 3528
rect 40166 3488 40500 3516
rect 40166 3485 40178 3488
rect 40120 3479 40178 3485
rect 40494 3476 40500 3488
rect 40552 3476 40558 3528
rect 42696 3519 42754 3525
rect 42696 3485 42708 3519
rect 42742 3516 42754 3519
rect 43070 3516 43076 3528
rect 42742 3488 43076 3516
rect 42742 3485 42754 3488
rect 42696 3479 42754 3485
rect 43070 3476 43076 3488
rect 43128 3476 43134 3528
rect 48222 3516 48228 3528
rect 48183 3488 48228 3516
rect 48222 3476 48228 3488
rect 48280 3476 48286 3528
rect 48492 3519 48550 3525
rect 48492 3485 48504 3519
rect 48538 3516 48550 3519
rect 48958 3516 48964 3528
rect 48538 3488 48964 3516
rect 48538 3485 48550 3488
rect 48492 3479 48550 3485
rect 48958 3476 48964 3488
rect 49016 3476 49022 3528
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50614 3525 50620 3528
rect 50341 3519 50399 3525
rect 50341 3516 50353 3519
rect 50212 3488 50353 3516
rect 50212 3476 50218 3488
rect 50341 3485 50353 3488
rect 50387 3485 50399 3519
rect 50608 3516 50620 3525
rect 50575 3488 50620 3516
rect 50341 3479 50399 3485
rect 50608 3479 50620 3488
rect 14360 3451 14418 3457
rect 14360 3417 14372 3451
rect 14406 3448 14418 3451
rect 14734 3448 14740 3460
rect 14406 3420 14740 3448
rect 14406 3417 14418 3420
rect 14360 3411 14418 3417
rect 14734 3408 14740 3420
rect 14792 3408 14798 3460
rect 18138 3408 18144 3460
rect 18196 3448 18202 3460
rect 19490 3451 19548 3457
rect 19490 3448 19502 3451
rect 18196 3420 19502 3448
rect 18196 3408 18202 3420
rect 19490 3417 19502 3420
rect 19536 3417 19548 3451
rect 19490 3411 19548 3417
rect 21352 3451 21410 3457
rect 21352 3417 21364 3451
rect 21398 3448 21410 3451
rect 23198 3448 23204 3460
rect 21398 3420 23204 3448
rect 21398 3417 21410 3420
rect 21352 3411 21410 3417
rect 23198 3408 23204 3420
rect 23256 3408 23262 3460
rect 25124 3451 25182 3457
rect 25124 3417 25136 3451
rect 25170 3448 25182 3451
rect 27338 3448 27344 3460
rect 25170 3420 27344 3448
rect 25170 3417 25182 3420
rect 25124 3411 25182 3417
rect 27338 3408 27344 3420
rect 27396 3408 27402 3460
rect 32852 3451 32910 3457
rect 32852 3417 32864 3451
rect 32898 3448 32910 3451
rect 33502 3448 33508 3460
rect 32898 3420 33508 3448
rect 32898 3417 32910 3420
rect 32852 3411 32910 3417
rect 33502 3408 33508 3420
rect 33560 3408 33566 3460
rect 34054 3408 34060 3460
rect 34112 3448 34118 3460
rect 34946 3451 35004 3457
rect 34946 3448 34958 3451
rect 34112 3420 34958 3448
rect 34112 3408 34118 3420
rect 34946 3417 34958 3420
rect 34992 3417 35004 3451
rect 34946 3411 35004 3417
rect 35894 3408 35900 3460
rect 35952 3448 35958 3460
rect 36786 3451 36844 3457
rect 36786 3448 36798 3451
rect 35952 3420 36798 3448
rect 35952 3408 35958 3420
rect 36786 3417 36798 3420
rect 36832 3417 36844 3451
rect 50356 3448 50384 3479
rect 50614 3476 50620 3479
rect 50672 3476 50678 3528
rect 52181 3519 52239 3525
rect 52181 3485 52193 3519
rect 52227 3516 52239 3519
rect 52730 3516 52736 3528
rect 52227 3488 52736 3516
rect 52227 3485 52239 3488
rect 52181 3479 52239 3485
rect 52196 3448 52224 3479
rect 52730 3476 52736 3488
rect 52788 3476 52794 3528
rect 50356 3420 52224 3448
rect 36786 3411 36844 3417
rect 52270 3408 52276 3460
rect 52328 3448 52334 3460
rect 52426 3451 52484 3457
rect 52426 3448 52438 3451
rect 52328 3420 52438 3448
rect 52328 3408 52334 3420
rect 52426 3417 52438 3420
rect 52472 3417 52484 3451
rect 52426 3411 52484 3417
rect 18046 3340 18052 3392
rect 18104 3380 18110 3392
rect 20625 3383 20683 3389
rect 20625 3380 20637 3383
rect 18104 3352 20637 3380
rect 18104 3340 18110 3352
rect 20625 3349 20637 3352
rect 20671 3349 20683 3383
rect 20625 3343 20683 3349
rect 26234 3340 26240 3392
rect 26292 3380 26298 3392
rect 28074 3380 28080 3392
rect 26292 3352 26337 3380
rect 28035 3352 28080 3380
rect 26292 3340 26298 3352
rect 28074 3340 28080 3352
rect 28132 3340 28138 3392
rect 33962 3380 33968 3392
rect 33923 3352 33968 3380
rect 33962 3340 33968 3352
rect 34020 3340 34026 3392
rect 36078 3380 36084 3392
rect 36039 3352 36084 3380
rect 36078 3340 36084 3352
rect 36136 3340 36142 3392
rect 36446 3340 36452 3392
rect 36504 3380 36510 3392
rect 37921 3383 37979 3389
rect 37921 3380 37933 3383
rect 36504 3352 37933 3380
rect 36504 3340 36510 3352
rect 37921 3349 37933 3352
rect 37967 3349 37979 3383
rect 51718 3380 51724 3392
rect 51679 3352 51724 3380
rect 37921 3343 37979 3349
rect 51718 3340 51724 3352
rect 51776 3340 51782 3392
rect 1104 3290 59340 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 59340 3290
rect 1104 3216 59340 3238
rect 14734 3176 14740 3188
rect 14695 3148 14740 3176
rect 14734 3136 14740 3148
rect 14792 3136 14798 3188
rect 18049 3179 18107 3185
rect 18049 3145 18061 3179
rect 18095 3176 18107 3179
rect 18138 3176 18144 3188
rect 18095 3148 18144 3176
rect 18095 3145 18107 3148
rect 18049 3139 18107 3145
rect 18138 3136 18144 3148
rect 18196 3136 18202 3188
rect 23845 3179 23903 3185
rect 23845 3145 23857 3179
rect 23891 3145 23903 3179
rect 25682 3176 25688 3188
rect 25643 3148 25688 3176
rect 23845 3139 23903 3145
rect 11784 3111 11842 3117
rect 11784 3077 11796 3111
rect 11830 3108 11842 3111
rect 12894 3108 12900 3120
rect 11830 3080 12900 3108
rect 11830 3077 11842 3080
rect 11784 3071 11842 3077
rect 12894 3068 12900 3080
rect 12952 3068 12958 3120
rect 13624 3111 13682 3117
rect 13624 3077 13636 3111
rect 13670 3108 13682 3111
rect 13814 3108 13820 3120
rect 13670 3080 13820 3108
rect 13670 3077 13682 3080
rect 13624 3071 13682 3077
rect 13814 3068 13820 3080
rect 13872 3068 13878 3120
rect 16936 3111 16994 3117
rect 16936 3077 16948 3111
rect 16982 3108 16994 3111
rect 17310 3108 17316 3120
rect 16982 3080 17316 3108
rect 16982 3077 16994 3080
rect 16936 3071 16994 3077
rect 17310 3068 17316 3080
rect 17368 3068 17374 3120
rect 19334 3108 19340 3120
rect 18524 3080 19340 3108
rect 10778 3000 10784 3052
rect 10836 3040 10842 3052
rect 11514 3040 11520 3052
rect 10836 3012 11520 3040
rect 10836 3000 10842 3012
rect 11514 3000 11520 3012
rect 11572 3040 11578 3052
rect 13354 3040 13360 3052
rect 11572 3012 13360 3040
rect 11572 3000 11578 3012
rect 13354 3000 13360 3012
rect 13412 3000 13418 3052
rect 16298 3000 16304 3052
rect 16356 3040 16362 3052
rect 16669 3043 16727 3049
rect 16669 3040 16681 3043
rect 16356 3012 16681 3040
rect 16356 3000 16362 3012
rect 16669 3009 16681 3012
rect 16715 3040 16727 3043
rect 17218 3040 17224 3052
rect 16715 3012 17224 3040
rect 16715 3009 16727 3012
rect 16669 3003 16727 3009
rect 17218 3000 17224 3012
rect 17276 3040 17282 3052
rect 18524 3049 18552 3080
rect 19334 3068 19340 3080
rect 19392 3068 19398 3120
rect 22738 3117 22744 3120
rect 22732 3108 22744 3117
rect 22699 3080 22744 3108
rect 22732 3071 22744 3080
rect 22738 3068 22744 3071
rect 22796 3068 22802 3120
rect 18509 3043 18567 3049
rect 18509 3040 18521 3043
rect 17276 3012 18521 3040
rect 17276 3000 17282 3012
rect 18509 3009 18521 3012
rect 18555 3009 18567 3043
rect 18509 3003 18567 3009
rect 18598 3000 18604 3052
rect 18656 3040 18662 3052
rect 18765 3043 18823 3049
rect 18765 3040 18777 3043
rect 18656 3012 18777 3040
rect 18656 3000 18662 3012
rect 18765 3009 18777 3012
rect 18811 3009 18823 3043
rect 18765 3003 18823 3009
rect 22465 3043 22523 3049
rect 22465 3009 22477 3043
rect 22511 3040 22523 3043
rect 23860 3040 23888 3139
rect 25682 3136 25688 3148
rect 25740 3136 25746 3188
rect 29638 3136 29644 3188
rect 29696 3176 29702 3188
rect 30193 3179 30251 3185
rect 30193 3176 30205 3179
rect 29696 3148 30205 3176
rect 29696 3136 29702 3148
rect 30193 3145 30205 3148
rect 30239 3145 30251 3179
rect 34054 3176 34060 3188
rect 34015 3148 34060 3176
rect 30193 3139 30251 3145
rect 34054 3136 34060 3148
rect 34112 3136 34118 3188
rect 35894 3136 35900 3188
rect 35952 3176 35958 3188
rect 35952 3148 35997 3176
rect 35952 3136 35958 3148
rect 40402 3136 40408 3188
rect 40460 3176 40466 3188
rect 40497 3179 40555 3185
rect 40497 3176 40509 3179
rect 40460 3148 40509 3176
rect 40460 3136 40466 3148
rect 40497 3145 40509 3148
rect 40543 3145 40555 3179
rect 40497 3139 40555 3145
rect 43530 3136 43536 3188
rect 43588 3176 43594 3188
rect 43809 3179 43867 3185
rect 43809 3176 43821 3179
rect 43588 3148 43821 3176
rect 43588 3136 43594 3148
rect 43809 3145 43821 3148
rect 43855 3145 43867 3179
rect 43809 3139 43867 3145
rect 52181 3179 52239 3185
rect 52181 3145 52193 3179
rect 52227 3176 52239 3179
rect 52270 3176 52276 3188
rect 52227 3148 52276 3176
rect 52227 3145 52239 3148
rect 52181 3139 52239 3145
rect 52270 3136 52276 3148
rect 52328 3136 52334 3188
rect 24572 3111 24630 3117
rect 24572 3077 24584 3111
rect 24618 3108 24630 3111
rect 26234 3108 26240 3120
rect 24618 3080 26240 3108
rect 24618 3077 24630 3080
rect 24572 3071 24630 3077
rect 26234 3068 26240 3080
rect 26292 3068 26298 3120
rect 27240 3111 27298 3117
rect 27240 3077 27252 3111
rect 27286 3108 27298 3111
rect 28074 3108 28080 3120
rect 27286 3080 28080 3108
rect 27286 3077 27298 3080
rect 27240 3071 27298 3077
rect 28074 3068 28080 3080
rect 28132 3068 28138 3120
rect 32944 3111 33002 3117
rect 32944 3077 32956 3111
rect 32990 3108 33002 3111
rect 33962 3108 33968 3120
rect 32990 3080 33968 3108
rect 32990 3077 33002 3080
rect 32944 3071 33002 3077
rect 33962 3068 33968 3080
rect 34020 3068 34026 3120
rect 34784 3111 34842 3117
rect 34784 3077 34796 3111
rect 34830 3108 34842 3111
rect 36078 3108 36084 3120
rect 34830 3080 36084 3108
rect 34830 3077 34842 3080
rect 34784 3071 34842 3077
rect 36078 3068 36084 3080
rect 36136 3068 36142 3120
rect 38654 3068 38660 3120
rect 38712 3108 38718 3120
rect 42702 3117 42708 3120
rect 39362 3111 39420 3117
rect 39362 3108 39374 3111
rect 38712 3080 39374 3108
rect 38712 3068 38718 3080
rect 39362 3077 39374 3080
rect 39408 3077 39420 3111
rect 42696 3108 42708 3117
rect 42663 3080 42708 3108
rect 39362 3071 39420 3077
rect 42696 3071 42708 3080
rect 42702 3068 42708 3071
rect 42760 3068 42766 3120
rect 51068 3111 51126 3117
rect 51068 3077 51080 3111
rect 51114 3108 51126 3111
rect 51718 3108 51724 3120
rect 51114 3080 51724 3108
rect 51114 3077 51126 3080
rect 51068 3071 51126 3077
rect 51718 3068 51724 3080
rect 51776 3068 51782 3120
rect 53000 3111 53058 3117
rect 53000 3077 53012 3111
rect 53046 3108 53058 3111
rect 54110 3108 54116 3120
rect 53046 3080 54116 3108
rect 53046 3077 53058 3080
rect 53000 3071 53058 3077
rect 54110 3068 54116 3080
rect 54168 3068 54174 3120
rect 29069 3043 29127 3049
rect 29069 3040 29081 3043
rect 22511 3012 23520 3040
rect 23860 3012 29081 3040
rect 22511 3009 22523 3012
rect 22465 3003 22523 3009
rect 23492 2972 23520 3012
rect 29069 3009 29081 3012
rect 29115 3009 29127 3043
rect 29069 3003 29127 3009
rect 32582 3000 32588 3052
rect 32640 3040 32646 3052
rect 32677 3043 32735 3049
rect 32677 3040 32689 3043
rect 32640 3012 32689 3040
rect 32640 3000 32646 3012
rect 32677 3009 32689 3012
rect 32723 3040 32735 3043
rect 34517 3043 34575 3049
rect 34517 3040 34529 3043
rect 32723 3012 34529 3040
rect 32723 3009 32735 3012
rect 32677 3003 32735 3009
rect 34517 3009 34529 3012
rect 34563 3040 34575 3043
rect 34606 3040 34612 3052
rect 34563 3012 34612 3040
rect 34563 3009 34575 3012
rect 34517 3003 34575 3009
rect 34606 3000 34612 3012
rect 34664 3000 34670 3052
rect 37274 3040 37280 3052
rect 37235 3012 37280 3040
rect 37274 3000 37280 3012
rect 37332 3000 37338 3052
rect 37550 3049 37556 3052
rect 37544 3003 37556 3049
rect 37608 3040 37614 3052
rect 39117 3043 39175 3049
rect 37608 3012 37644 3040
rect 37550 3000 37556 3003
rect 37608 3000 37614 3012
rect 39117 3009 39129 3043
rect 39163 3040 39175 3043
rect 39850 3040 39856 3052
rect 39163 3012 39856 3040
rect 39163 3009 39175 3012
rect 39117 3003 39175 3009
rect 39850 3000 39856 3012
rect 39908 3000 39914 3052
rect 42426 3040 42432 3052
rect 42387 3012 42432 3040
rect 42426 3000 42432 3012
rect 42484 3000 42490 3052
rect 48222 3000 48228 3052
rect 48280 3040 48286 3052
rect 50801 3043 50859 3049
rect 50801 3040 50813 3043
rect 48280 3012 50813 3040
rect 48280 3000 48286 3012
rect 50801 3009 50813 3012
rect 50847 3009 50859 3043
rect 52730 3040 52736 3052
rect 52691 3012 52736 3040
rect 50801 3003 50859 3009
rect 52730 3000 52736 3012
rect 52788 3000 52794 3052
rect 24026 2972 24032 2984
rect 23492 2944 24032 2972
rect 24026 2932 24032 2944
rect 24084 2972 24090 2984
rect 24305 2975 24363 2981
rect 24305 2972 24317 2975
rect 24084 2944 24317 2972
rect 24084 2932 24090 2944
rect 24305 2941 24317 2944
rect 24351 2941 24363 2975
rect 26970 2972 26976 2984
rect 26931 2944 26976 2972
rect 24305 2935 24363 2941
rect 24320 2848 24348 2935
rect 26970 2932 26976 2944
rect 27028 2932 27034 2984
rect 28813 2975 28871 2981
rect 28813 2941 28825 2975
rect 28859 2941 28871 2975
rect 28813 2935 28871 2941
rect 28828 2904 28856 2935
rect 27908 2876 28856 2904
rect 38657 2907 38715 2913
rect 12894 2836 12900 2848
rect 12855 2808 12900 2836
rect 12894 2796 12900 2808
rect 12952 2796 12958 2848
rect 19889 2839 19947 2845
rect 19889 2805 19901 2839
rect 19935 2836 19947 2839
rect 19978 2836 19984 2848
rect 19935 2808 19984 2836
rect 19935 2805 19947 2808
rect 19889 2799 19947 2805
rect 19978 2796 19984 2808
rect 20036 2796 20042 2848
rect 24302 2836 24308 2848
rect 24215 2808 24308 2836
rect 24302 2796 24308 2808
rect 24360 2836 24366 2848
rect 27908 2836 27936 2876
rect 38657 2873 38669 2907
rect 38703 2904 38715 2907
rect 38838 2904 38844 2916
rect 38703 2876 38844 2904
rect 38703 2873 38715 2876
rect 38657 2867 38715 2873
rect 38838 2864 38844 2876
rect 38896 2864 38902 2916
rect 54018 2864 54024 2916
rect 54076 2904 54082 2916
rect 54113 2907 54171 2913
rect 54113 2904 54125 2907
rect 54076 2876 54125 2904
rect 54076 2864 54082 2876
rect 54113 2873 54125 2876
rect 54159 2873 54171 2907
rect 54113 2867 54171 2873
rect 28350 2836 28356 2848
rect 24360 2808 27936 2836
rect 28311 2808 28356 2836
rect 24360 2796 24366 2808
rect 28350 2796 28356 2808
rect 28408 2796 28414 2848
rect 1104 2746 59340 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 59340 2746
rect 1104 2672 59340 2694
rect 18598 2632 18604 2644
rect 6886 2604 18460 2632
rect 18559 2604 18604 2632
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2428 1731 2431
rect 1949 2431 2007 2437
rect 1949 2428 1961 2431
rect 1719 2400 1961 2428
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 1949 2397 1961 2400
rect 1995 2428 2007 2431
rect 6886 2428 6914 2604
rect 13078 2564 13084 2576
rect 13039 2536 13084 2564
rect 13078 2524 13084 2536
rect 13136 2524 13142 2576
rect 18432 2564 18460 2604
rect 18598 2592 18604 2604
rect 18656 2592 18662 2644
rect 23198 2632 23204 2644
rect 18708 2604 22876 2632
rect 23159 2604 23204 2632
rect 18708 2564 18736 2604
rect 18432 2536 18736 2564
rect 11514 2456 11520 2508
rect 11572 2496 11578 2508
rect 11701 2499 11759 2505
rect 11701 2496 11713 2499
rect 11572 2468 11713 2496
rect 11572 2456 11578 2468
rect 11701 2465 11713 2468
rect 11747 2465 11759 2499
rect 17218 2496 17224 2508
rect 17179 2468 17224 2496
rect 11701 2459 11759 2465
rect 17218 2456 17224 2468
rect 17276 2456 17282 2508
rect 1995 2400 6914 2428
rect 11968 2431 12026 2437
rect 1995 2397 2007 2400
rect 1949 2391 2007 2397
rect 11968 2397 11980 2431
rect 12014 2428 12026 2431
rect 12894 2428 12900 2440
rect 12014 2400 12900 2428
rect 12014 2397 12026 2400
rect 11968 2391 12026 2397
rect 12894 2388 12900 2400
rect 12952 2388 12958 2440
rect 17488 2431 17546 2437
rect 17488 2397 17500 2431
rect 17534 2428 17546 2431
rect 18046 2428 18052 2440
rect 17534 2400 18052 2428
rect 17534 2397 17546 2400
rect 17488 2391 17546 2397
rect 18046 2388 18052 2400
rect 18104 2388 18110 2440
rect 19889 2431 19947 2437
rect 19889 2397 19901 2431
rect 19935 2397 19947 2431
rect 19889 2391 19947 2397
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1765 2363 1823 2369
rect 1765 2360 1777 2363
rect 72 2332 1777 2360
rect 72 2320 78 2332
rect 1765 2329 1777 2332
rect 1811 2329 1823 2363
rect 19904 2360 19932 2391
rect 19978 2388 19984 2440
rect 20036 2428 20042 2440
rect 20145 2431 20203 2437
rect 20145 2428 20157 2431
rect 20036 2400 20157 2428
rect 20036 2388 20042 2400
rect 20145 2397 20157 2400
rect 20191 2397 20203 2431
rect 20145 2391 20203 2397
rect 20622 2388 20628 2440
rect 20680 2428 20686 2440
rect 21821 2431 21879 2437
rect 21821 2428 21833 2431
rect 20680 2400 21833 2428
rect 20680 2388 20686 2400
rect 21821 2397 21833 2400
rect 21867 2397 21879 2431
rect 21821 2391 21879 2397
rect 20640 2360 20668 2388
rect 22066 2363 22124 2369
rect 22066 2360 22078 2363
rect 19904 2332 20668 2360
rect 21284 2332 22078 2360
rect 1765 2323 1823 2329
rect 21284 2301 21312 2332
rect 22066 2329 22078 2332
rect 22112 2329 22124 2363
rect 22848 2360 22876 2604
rect 23198 2592 23204 2604
rect 23256 2592 23262 2644
rect 25774 2632 25780 2644
rect 25735 2604 25780 2632
rect 25774 2592 25780 2604
rect 25832 2592 25838 2644
rect 27338 2592 27344 2644
rect 27396 2632 27402 2644
rect 28353 2635 28411 2641
rect 28353 2632 28365 2635
rect 27396 2604 28365 2632
rect 27396 2592 27402 2604
rect 28353 2601 28365 2604
rect 28399 2601 28411 2635
rect 28353 2595 28411 2601
rect 33502 2592 33508 2644
rect 33560 2632 33566 2644
rect 33965 2635 34023 2641
rect 33965 2632 33977 2635
rect 33560 2604 33977 2632
rect 33560 2592 33566 2604
rect 33965 2601 33977 2604
rect 34011 2601 34023 2635
rect 33965 2595 34023 2601
rect 36081 2635 36139 2641
rect 36081 2601 36093 2635
rect 36127 2632 36139 2635
rect 37550 2632 37556 2644
rect 36127 2604 37556 2632
rect 36127 2601 36139 2604
rect 36081 2595 36139 2601
rect 37550 2592 37556 2604
rect 37608 2592 37614 2644
rect 38657 2635 38715 2641
rect 38657 2601 38669 2635
rect 38703 2632 38715 2635
rect 38746 2632 38752 2644
rect 38703 2604 38752 2632
rect 38703 2601 38715 2604
rect 38657 2595 38715 2601
rect 38746 2592 38752 2604
rect 38804 2592 38810 2644
rect 24302 2456 24308 2508
rect 24360 2496 24366 2508
rect 24397 2499 24455 2505
rect 24397 2496 24409 2499
rect 24360 2468 24409 2496
rect 24360 2456 24366 2468
rect 24397 2465 24409 2468
rect 24443 2465 24455 2499
rect 26970 2496 26976 2508
rect 26931 2468 26976 2496
rect 24397 2459 24455 2465
rect 26970 2456 26976 2468
rect 27028 2456 27034 2508
rect 34606 2456 34612 2508
rect 34664 2496 34670 2508
rect 34701 2499 34759 2505
rect 34701 2496 34713 2499
rect 34664 2468 34713 2496
rect 34664 2456 34670 2468
rect 34701 2465 34713 2468
rect 34747 2465 34759 2499
rect 37274 2496 37280 2508
rect 37235 2468 37280 2496
rect 34701 2459 34759 2465
rect 37274 2456 37280 2468
rect 37332 2456 37338 2508
rect 24664 2431 24722 2437
rect 24664 2397 24676 2431
rect 24710 2428 24722 2431
rect 25406 2428 25412 2440
rect 24710 2400 25412 2428
rect 24710 2397 24722 2400
rect 24664 2391 24722 2397
rect 25406 2388 25412 2400
rect 25464 2388 25470 2440
rect 27240 2431 27298 2437
rect 27240 2397 27252 2431
rect 27286 2428 27298 2431
rect 28350 2428 28356 2440
rect 27286 2400 28356 2428
rect 27286 2397 27298 2400
rect 27240 2391 27298 2397
rect 28350 2388 28356 2400
rect 28408 2388 28414 2440
rect 34149 2431 34207 2437
rect 34149 2397 34161 2431
rect 34195 2428 34207 2431
rect 34238 2428 34244 2440
rect 34195 2400 34244 2428
rect 34195 2397 34207 2400
rect 34149 2391 34207 2397
rect 34238 2388 34244 2400
rect 34296 2388 34302 2440
rect 34968 2431 35026 2437
rect 34968 2397 34980 2431
rect 35014 2428 35026 2431
rect 36446 2428 36452 2440
rect 35014 2400 36452 2428
rect 35014 2397 35026 2400
rect 34968 2391 35026 2397
rect 36446 2388 36452 2400
rect 36504 2388 36510 2440
rect 37544 2431 37602 2437
rect 37544 2397 37556 2431
rect 37590 2428 37602 2431
rect 38562 2428 38568 2440
rect 37590 2400 38568 2428
rect 37590 2397 37602 2400
rect 37544 2391 37602 2397
rect 38562 2388 38568 2400
rect 38620 2388 38626 2440
rect 28534 2360 28540 2372
rect 22848 2332 28540 2360
rect 22066 2323 22124 2329
rect 28534 2320 28540 2332
rect 28592 2320 28598 2372
rect 21269 2295 21327 2301
rect 21269 2261 21281 2295
rect 21315 2261 21327 2295
rect 21269 2255 21327 2261
rect 1104 2202 59340 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 59340 2202
rect 1104 2128 59340 2150
<< via1 >>
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 34934 60358 34986 60410
rect 34998 60358 35050 60410
rect 35062 60358 35114 60410
rect 35126 60358 35178 60410
rect 35190 60358 35242 60410
rect 26240 60188 26292 60240
rect 60372 60188 60424 60240
rect 11520 60052 11572 60104
rect 29920 60095 29972 60104
rect 29920 60061 29929 60095
rect 29929 60061 29963 60095
rect 29963 60061 29972 60095
rect 29920 60052 29972 60061
rect 32128 60095 32180 60104
rect 7748 59984 7800 60036
rect 12900 59984 12952 60036
rect 28448 59984 28500 60036
rect 32128 60061 32137 60095
rect 32137 60061 32171 60095
rect 32171 60061 32180 60095
rect 32128 60052 32180 60061
rect 34060 60052 34112 60104
rect 37556 60052 37608 60104
rect 40408 60052 40460 60104
rect 43628 60052 43680 60104
rect 45560 60052 45612 60104
rect 48964 60052 49016 60104
rect 50804 60052 50856 60104
rect 54116 60052 54168 60104
rect 6920 59916 6972 59968
rect 8484 59916 8536 59968
rect 13084 59959 13136 59968
rect 13084 59925 13093 59959
rect 13093 59925 13127 59959
rect 13127 59925 13136 59959
rect 13084 59916 13136 59925
rect 29368 59916 29420 59968
rect 31576 59984 31628 60036
rect 36728 59959 36780 59968
rect 36728 59925 36737 59959
rect 36737 59925 36771 59959
rect 36771 59925 36780 59959
rect 36728 59916 36780 59925
rect 38752 59984 38804 60036
rect 46940 59984 46992 60036
rect 49332 59984 49384 60036
rect 50620 59984 50672 60036
rect 54944 59984 54996 60036
rect 58440 60027 58492 60036
rect 58440 59993 58449 60027
rect 58449 59993 58483 60027
rect 58483 59993 58492 60027
rect 58440 59984 58492 59993
rect 44180 59916 44232 59968
rect 48780 59916 48832 59968
rect 51540 59959 51592 59968
rect 51540 59925 51549 59959
rect 51549 59925 51583 59959
rect 51583 59925 51592 59959
rect 51540 59916 51592 59925
rect 53196 59916 53248 59968
rect 19574 59814 19626 59866
rect 19638 59814 19690 59866
rect 19702 59814 19754 59866
rect 19766 59814 19818 59866
rect 19830 59814 19882 59866
rect 50294 59814 50346 59866
rect 50358 59814 50410 59866
rect 50422 59814 50474 59866
rect 50486 59814 50538 59866
rect 50550 59814 50602 59866
rect 7748 59755 7800 59764
rect 7748 59721 7757 59755
rect 7757 59721 7791 59755
rect 7791 59721 7800 59755
rect 7748 59712 7800 59721
rect 12900 59755 12952 59764
rect 12900 59721 12909 59755
rect 12909 59721 12943 59755
rect 12943 59721 12952 59755
rect 12900 59712 12952 59721
rect 31576 59755 31628 59764
rect 31576 59721 31585 59755
rect 31585 59721 31619 59755
rect 31619 59721 31628 59755
rect 31576 59712 31628 59721
rect 6920 59644 6972 59696
rect 8116 59576 8168 59628
rect 9496 59576 9548 59628
rect 12256 59576 12308 59628
rect 14648 59576 14700 59628
rect 19984 59576 20036 59628
rect 21180 59576 21232 59628
rect 23848 59576 23900 59628
rect 25964 59576 26016 59628
rect 27528 59644 27580 59696
rect 38752 59712 38804 59764
rect 46940 59755 46992 59764
rect 46940 59721 46949 59755
rect 46949 59721 46983 59755
rect 46983 59721 46992 59755
rect 46940 59712 46992 59721
rect 54944 59755 54996 59764
rect 54944 59721 54953 59755
rect 54953 59721 54987 59755
rect 54987 59721 54996 59755
rect 54944 59712 54996 59721
rect 34060 59644 34112 59696
rect 55404 59644 55456 59696
rect 28540 59576 28592 59628
rect 29920 59576 29972 59628
rect 30288 59576 30340 59628
rect 31760 59576 31812 59628
rect 35440 59576 35492 59628
rect 37556 59619 37608 59628
rect 37556 59585 37565 59619
rect 37565 59585 37599 59619
rect 37599 59585 37608 59619
rect 37556 59576 37608 59585
rect 39028 59576 39080 59628
rect 41880 59576 41932 59628
rect 44456 59576 44508 59628
rect 45560 59619 45612 59628
rect 45560 59585 45569 59619
rect 45569 59585 45603 59619
rect 45603 59585 45612 59619
rect 45560 59576 45612 59585
rect 47032 59576 47084 59628
rect 48964 59576 49016 59628
rect 49516 59576 49568 59628
rect 51908 59576 51960 59628
rect 54760 59576 54812 59628
rect 54852 59576 54904 59628
rect 11520 59551 11572 59560
rect 11520 59517 11529 59551
rect 11529 59517 11563 59551
rect 11563 59517 11572 59551
rect 11520 59508 11572 59517
rect 22468 59551 22520 59560
rect 22468 59517 22477 59551
rect 22477 59517 22511 59551
rect 22511 59517 22520 59551
rect 22468 59508 22520 59517
rect 32128 59508 32180 59560
rect 34428 59551 34480 59560
rect 9588 59415 9640 59424
rect 9588 59381 9597 59415
rect 9597 59381 9631 59415
rect 9631 59381 9640 59415
rect 9588 59372 9640 59381
rect 14740 59415 14792 59424
rect 14740 59381 14749 59415
rect 14749 59381 14783 59415
rect 14783 59381 14792 59415
rect 14740 59372 14792 59381
rect 20168 59372 20220 59424
rect 23480 59372 23532 59424
rect 23940 59372 23992 59424
rect 27252 59372 27304 59424
rect 34428 59517 34437 59551
rect 34437 59517 34471 59551
rect 34471 59517 34480 59551
rect 34428 59508 34480 59517
rect 40408 59551 40460 59560
rect 40408 59517 40417 59551
rect 40417 59517 40451 59551
rect 40451 59517 40460 59551
rect 40408 59508 40460 59517
rect 43628 59551 43680 59560
rect 43628 59517 43637 59551
rect 43637 59517 43671 59551
rect 43671 59517 43680 59551
rect 43628 59508 43680 59517
rect 50804 59551 50856 59560
rect 50804 59517 50813 59551
rect 50813 59517 50847 59551
rect 50847 59517 50856 59551
rect 50804 59508 50856 59517
rect 53380 59508 53432 59560
rect 55864 59508 55916 59560
rect 32864 59372 32916 59424
rect 34612 59372 34664 59424
rect 40684 59372 40736 59424
rect 43352 59372 43404 59424
rect 48504 59372 48556 59424
rect 51080 59372 51132 59424
rect 55956 59372 56008 59424
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 34934 59270 34986 59322
rect 34998 59270 35050 59322
rect 35062 59270 35114 59322
rect 35126 59270 35178 59322
rect 35190 59270 35242 59322
rect 8116 59211 8168 59220
rect 8116 59177 8125 59211
rect 8125 59177 8159 59211
rect 8159 59177 8168 59211
rect 8116 59168 8168 59177
rect 23848 59211 23900 59220
rect 23848 59177 23857 59211
rect 23857 59177 23891 59211
rect 23891 59177 23900 59211
rect 23848 59168 23900 59177
rect 27528 59168 27580 59220
rect 39028 59211 39080 59220
rect 39028 59177 39037 59211
rect 39037 59177 39071 59211
rect 39071 59177 39080 59211
rect 39028 59168 39080 59177
rect 44456 59211 44508 59220
rect 44456 59177 44465 59211
rect 44465 59177 44499 59211
rect 44499 59177 44508 59211
rect 44456 59168 44508 59177
rect 54760 59211 54812 59220
rect 54760 59177 54769 59211
rect 54769 59177 54803 59211
rect 54803 59177 54812 59211
rect 54760 59168 54812 59177
rect 57520 59168 57572 59220
rect 58440 59168 58492 59220
rect 37556 59032 37608 59084
rect 6184 58964 6236 59016
rect 6828 58964 6880 59016
rect 8208 58964 8260 59016
rect 9588 58964 9640 59016
rect 11520 58964 11572 59016
rect 14096 59007 14148 59016
rect 14096 58973 14105 59007
rect 14105 58973 14139 59007
rect 14139 58973 14148 59007
rect 14096 58964 14148 58973
rect 14740 58964 14792 59016
rect 15936 59007 15988 59016
rect 15936 58973 15945 59007
rect 15945 58973 15979 59007
rect 15979 58973 15988 59007
rect 15936 58964 15988 58973
rect 19984 58964 20036 59016
rect 27252 58964 27304 59016
rect 27528 58964 27580 59016
rect 29368 58964 29420 59016
rect 30288 59007 30340 59016
rect 30288 58973 30297 59007
rect 30297 58973 30331 59007
rect 30331 58973 30340 59007
rect 30288 58964 30340 58973
rect 32864 58964 32916 59016
rect 34520 58964 34572 59016
rect 35348 58964 35400 59016
rect 36728 58964 36780 59016
rect 42800 58964 42852 59016
rect 48964 58964 49016 59016
rect 50804 58964 50856 59016
rect 53196 58964 53248 59016
rect 53380 59007 53432 59016
rect 53380 58973 53389 59007
rect 53389 58973 53423 59007
rect 53423 58973 53432 59007
rect 53380 58964 53432 58973
rect 55404 58964 55456 59016
rect 57060 58964 57112 59016
rect 6000 58896 6052 58948
rect 7748 58896 7800 58948
rect 12808 58896 12860 58948
rect 15844 58896 15896 58948
rect 21272 58896 21324 58948
rect 23848 58896 23900 58948
rect 6276 58871 6328 58880
rect 6276 58837 6285 58871
rect 6285 58837 6319 58871
rect 6319 58837 6328 58871
rect 6276 58828 6328 58837
rect 10324 58871 10376 58880
rect 10324 58837 10333 58871
rect 10333 58837 10367 58871
rect 10367 58837 10376 58871
rect 10324 58828 10376 58837
rect 12164 58871 12216 58880
rect 12164 58837 12173 58871
rect 12173 58837 12207 58871
rect 12207 58837 12216 58871
rect 12164 58828 12216 58837
rect 15476 58871 15528 58880
rect 15476 58837 15485 58871
rect 15485 58837 15519 58871
rect 15519 58837 15528 58871
rect 15476 58828 15528 58837
rect 17316 58871 17368 58880
rect 17316 58837 17325 58871
rect 17325 58837 17359 58871
rect 17359 58837 17368 58871
rect 17316 58828 17368 58837
rect 21916 58871 21968 58880
rect 21916 58837 21925 58871
rect 21925 58837 21959 58871
rect 21959 58837 21968 58871
rect 21916 58828 21968 58837
rect 27160 58871 27212 58880
rect 27160 58837 27169 58871
rect 27169 58837 27203 58871
rect 27203 58837 27212 58871
rect 27160 58828 27212 58837
rect 29000 58871 29052 58880
rect 29000 58837 29009 58871
rect 29009 58837 29043 58871
rect 29043 58837 29052 58871
rect 29000 58828 29052 58837
rect 31668 58871 31720 58880
rect 31668 58837 31677 58871
rect 31677 58837 31711 58871
rect 31711 58837 31720 58871
rect 31668 58828 31720 58837
rect 31852 58896 31904 58948
rect 38844 58896 38896 58948
rect 43168 58896 43220 58948
rect 45192 58896 45244 58948
rect 47308 58896 47360 58948
rect 49424 58896 49476 58948
rect 54760 58896 54812 58948
rect 56784 58896 56836 58948
rect 37004 58871 37056 58880
rect 37004 58837 37013 58871
rect 37013 58837 37047 58871
rect 37047 58837 37056 58871
rect 37004 58828 37056 58837
rect 42616 58871 42668 58880
rect 42616 58837 42625 58871
rect 42625 58837 42659 58871
rect 42659 58837 42668 58871
rect 42616 58828 42668 58837
rect 47768 58871 47820 58880
rect 47768 58837 47777 58871
rect 47777 58837 47811 58871
rect 47811 58837 47820 58871
rect 47768 58828 47820 58837
rect 48320 58828 48372 58880
rect 52552 58828 52604 58880
rect 58624 58871 58676 58880
rect 58624 58837 58633 58871
rect 58633 58837 58667 58871
rect 58667 58837 58676 58871
rect 58624 58828 58676 58837
rect 19574 58726 19626 58778
rect 19638 58726 19690 58778
rect 19702 58726 19754 58778
rect 19766 58726 19818 58778
rect 19830 58726 19882 58778
rect 50294 58726 50346 58778
rect 50358 58726 50410 58778
rect 50422 58726 50474 58778
rect 50486 58726 50538 58778
rect 50550 58726 50602 58778
rect 7748 58667 7800 58676
rect 7748 58633 7757 58667
rect 7757 58633 7791 58667
rect 7791 58633 7800 58667
rect 7748 58624 7800 58633
rect 9496 58624 9548 58676
rect 14648 58624 14700 58676
rect 21180 58624 21232 58676
rect 25964 58667 26016 58676
rect 25964 58633 25973 58667
rect 25973 58633 26007 58667
rect 26007 58633 26016 58667
rect 25964 58624 26016 58633
rect 31760 58624 31812 58676
rect 38844 58667 38896 58676
rect 38844 58633 38853 58667
rect 38853 58633 38887 58667
rect 38887 58633 38896 58667
rect 38844 58624 38896 58633
rect 41880 58667 41932 58676
rect 41880 58633 41889 58667
rect 41889 58633 41923 58667
rect 41923 58633 41932 58667
rect 41880 58624 41932 58633
rect 45192 58667 45244 58676
rect 45192 58633 45201 58667
rect 45201 58633 45235 58667
rect 45235 58633 45244 58667
rect 45192 58624 45244 58633
rect 47032 58667 47084 58676
rect 47032 58633 47041 58667
rect 47041 58633 47075 58667
rect 47075 58633 47084 58667
rect 47032 58624 47084 58633
rect 6184 58556 6236 58608
rect 6276 58556 6328 58608
rect 8484 58599 8536 58608
rect 8484 58565 8518 58599
rect 8518 58565 8536 58599
rect 8484 58556 8536 58565
rect 12164 58556 12216 58608
rect 13084 58556 13136 58608
rect 21916 58556 21968 58608
rect 23940 58556 23992 58608
rect 29000 58556 29052 58608
rect 31668 58556 31720 58608
rect 39028 58556 39080 58608
rect 42616 58556 42668 58608
rect 44180 58556 44232 58608
rect 47768 58556 47820 58608
rect 5172 58488 5224 58540
rect 6920 58488 6972 58540
rect 8208 58531 8260 58540
rect 8208 58497 8217 58531
rect 8217 58497 8251 58531
rect 8251 58497 8260 58531
rect 8208 58488 8260 58497
rect 14096 58488 14148 58540
rect 19156 58488 19208 58540
rect 19984 58488 20036 58540
rect 22468 58488 22520 58540
rect 26424 58488 26476 58540
rect 30288 58488 30340 58540
rect 37280 58488 37332 58540
rect 37556 58488 37608 58540
rect 38568 58488 38620 58540
rect 43628 58488 43680 58540
rect 45560 58488 45612 58540
rect 47124 58488 47176 58540
rect 53104 58556 53156 58608
rect 55956 58556 56008 58608
rect 58624 58556 58676 58608
rect 52920 58488 52972 58540
rect 54116 58531 54168 58540
rect 54116 58497 54125 58531
rect 54125 58497 54159 58531
rect 54159 58497 54168 58531
rect 54116 58488 54168 58497
rect 55220 58488 55272 58540
rect 55864 58488 55916 58540
rect 6276 58420 6328 58472
rect 11520 58463 11572 58472
rect 11520 58429 11529 58463
rect 11529 58429 11563 58463
rect 11563 58429 11572 58463
rect 11520 58420 11572 58429
rect 18052 58463 18104 58472
rect 18052 58429 18061 58463
rect 18061 58429 18095 58463
rect 18095 58429 18104 58463
rect 18052 58420 18104 58429
rect 27528 58420 27580 58472
rect 40408 58420 40460 58472
rect 50804 58463 50856 58472
rect 50804 58429 50813 58463
rect 50813 58429 50847 58463
rect 50847 58429 50856 58463
rect 50804 58420 50856 58429
rect 57060 58488 57112 58540
rect 5540 58327 5592 58336
rect 5540 58293 5549 58327
rect 5549 58293 5583 58327
rect 5583 58293 5592 58327
rect 5540 58284 5592 58293
rect 12900 58327 12952 58336
rect 12900 58293 12909 58327
rect 12909 58293 12943 58327
rect 12943 58293 12952 58327
rect 12900 58284 12952 58293
rect 19340 58284 19392 58336
rect 24124 58327 24176 58336
rect 24124 58293 24133 58327
rect 24133 58293 24167 58327
rect 24167 58293 24176 58327
rect 24124 58284 24176 58293
rect 29276 58327 29328 58336
rect 29276 58293 29285 58327
rect 29285 58293 29319 58327
rect 29319 58293 29328 58327
rect 29276 58284 29328 58293
rect 35348 58327 35400 58336
rect 35348 58293 35357 58327
rect 35357 58293 35391 58327
rect 35391 58293 35400 58327
rect 35348 58284 35400 58293
rect 48964 58284 49016 58336
rect 52184 58327 52236 58336
rect 52184 58293 52193 58327
rect 52193 58293 52227 58327
rect 52227 58293 52236 58327
rect 52184 58284 52236 58293
rect 54392 58284 54444 58336
rect 56876 58284 56928 58336
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 34934 58182 34986 58234
rect 34998 58182 35050 58234
rect 35062 58182 35114 58234
rect 35126 58182 35178 58234
rect 35190 58182 35242 58234
rect 5172 58123 5224 58132
rect 5172 58089 5181 58123
rect 5181 58089 5215 58123
rect 5215 58089 5224 58123
rect 5172 58080 5224 58089
rect 38568 58123 38620 58132
rect 38568 58089 38577 58123
rect 38577 58089 38611 58123
rect 38611 58089 38620 58123
rect 38568 58080 38620 58089
rect 47308 58080 47360 58132
rect 19984 58012 20036 58064
rect 3884 57876 3936 57928
rect 6920 57876 6972 57928
rect 4988 57808 5040 57860
rect 5540 57808 5592 57860
rect 10324 57876 10376 57928
rect 15936 57944 15988 57996
rect 40408 57987 40460 57996
rect 10784 57919 10836 57928
rect 10784 57885 10793 57919
rect 10793 57885 10827 57919
rect 10827 57885 10836 57919
rect 10784 57876 10836 57885
rect 40408 57953 40417 57987
rect 40417 57953 40451 57987
rect 40451 57953 40460 57987
rect 40408 57944 40460 57953
rect 48964 58080 49016 58132
rect 52920 58123 52972 58132
rect 52920 58089 52929 58123
rect 52929 58089 52963 58123
rect 52963 58089 52972 58123
rect 52920 58080 52972 58089
rect 54760 58123 54812 58132
rect 54760 58089 54769 58123
rect 54769 58089 54803 58123
rect 54803 58089 54812 58123
rect 54760 58080 54812 58089
rect 18052 57876 18104 57928
rect 25044 57876 25096 57928
rect 27528 57876 27580 57928
rect 29276 57876 29328 57928
rect 30288 57876 30340 57928
rect 32864 57876 32916 57928
rect 34612 57876 34664 57928
rect 34704 57876 34756 57928
rect 35348 57919 35400 57928
rect 35348 57885 35357 57919
rect 35357 57885 35391 57919
rect 35391 57885 35400 57919
rect 35348 57876 35400 57885
rect 37004 57876 37056 57928
rect 37280 57876 37332 57928
rect 40684 57919 40736 57928
rect 40684 57885 40718 57919
rect 40718 57885 40736 57919
rect 40684 57876 40736 57885
rect 43352 57919 43404 57928
rect 43352 57885 43386 57919
rect 43386 57885 43404 57919
rect 13820 57808 13872 57860
rect 18604 57808 18656 57860
rect 20444 57851 20496 57860
rect 20444 57817 20453 57851
rect 20453 57817 20487 57851
rect 20487 57817 20496 57851
rect 20444 57808 20496 57817
rect 28908 57808 28960 57860
rect 32220 57808 32272 57860
rect 38660 57808 38712 57860
rect 43352 57876 43404 57885
rect 44272 57808 44324 57860
rect 48780 57876 48832 57928
rect 50804 57876 50856 57928
rect 53380 57919 53432 57928
rect 53380 57885 53389 57919
rect 53389 57885 53423 57919
rect 53423 57885 53432 57919
rect 53380 57876 53432 57885
rect 54392 57876 54444 57928
rect 55220 57876 55272 57928
rect 57060 57876 57112 57928
rect 51080 57808 51132 57860
rect 52828 57808 52880 57860
rect 6000 57740 6052 57792
rect 8944 57740 8996 57792
rect 10784 57740 10836 57792
rect 12164 57783 12216 57792
rect 12164 57749 12173 57783
rect 12173 57749 12207 57783
rect 12207 57749 12216 57783
rect 12164 57740 12216 57749
rect 14096 57740 14148 57792
rect 18696 57783 18748 57792
rect 18696 57749 18705 57783
rect 18705 57749 18739 57783
rect 18739 57749 18748 57783
rect 18696 57740 18748 57749
rect 27252 57740 27304 57792
rect 29000 57783 29052 57792
rect 29000 57749 29009 57783
rect 29009 57749 29043 57783
rect 29043 57749 29052 57783
rect 29000 57740 29052 57749
rect 32312 57783 32364 57792
rect 32312 57749 32321 57783
rect 32321 57749 32355 57783
rect 32355 57749 32364 57783
rect 32312 57740 32364 57749
rect 34152 57783 34204 57792
rect 34152 57749 34161 57783
rect 34161 57749 34195 57783
rect 34195 57749 34204 57783
rect 34152 57740 34204 57749
rect 35440 57740 35492 57792
rect 41144 57740 41196 57792
rect 43168 57740 43220 57792
rect 49608 57783 49660 57792
rect 49608 57749 49617 57783
rect 49617 57749 49651 57783
rect 49651 57749 49660 57783
rect 49608 57740 49660 57749
rect 56600 57740 56652 57792
rect 58440 57808 58492 57860
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 4988 57579 5040 57588
rect 4988 57545 4997 57579
rect 4997 57545 5031 57579
rect 5031 57545 5040 57579
rect 4988 57536 5040 57545
rect 12808 57536 12860 57588
rect 21272 57579 21324 57588
rect 21272 57545 21281 57579
rect 21281 57545 21315 57579
rect 21315 57545 21324 57579
rect 21272 57536 21324 57545
rect 26424 57579 26476 57588
rect 26424 57545 26433 57579
rect 26433 57545 26467 57579
rect 26467 57545 26476 57579
rect 26424 57536 26476 57545
rect 31852 57536 31904 57588
rect 40408 57536 40460 57588
rect 49516 57536 49568 57588
rect 53380 57536 53432 57588
rect 12164 57468 12216 57520
rect 15476 57468 15528 57520
rect 20628 57468 20680 57520
rect 24124 57468 24176 57520
rect 27160 57468 27212 57520
rect 29000 57468 29052 57520
rect 32312 57468 32364 57520
rect 34152 57468 34204 57520
rect 39028 57511 39080 57520
rect 39028 57477 39037 57511
rect 39037 57477 39071 57511
rect 39071 57477 39080 57511
rect 39028 57468 39080 57477
rect 41788 57468 41840 57520
rect 5172 57400 5224 57452
rect 8300 57400 8352 57452
rect 8760 57443 8812 57452
rect 8760 57409 8769 57443
rect 8769 57409 8803 57443
rect 8803 57409 8812 57443
rect 8760 57400 8812 57409
rect 13820 57400 13872 57452
rect 14096 57443 14148 57452
rect 14096 57409 14105 57443
rect 14105 57409 14139 57443
rect 14139 57409 14148 57443
rect 14096 57400 14148 57409
rect 18052 57443 18104 57452
rect 18052 57409 18061 57443
rect 18061 57409 18095 57443
rect 18095 57409 18104 57443
rect 19892 57443 19944 57452
rect 18052 57400 18104 57409
rect 19892 57409 19901 57443
rect 19901 57409 19935 57443
rect 19935 57409 19944 57443
rect 19892 57400 19944 57409
rect 23756 57400 23808 57452
rect 30288 57400 30340 57452
rect 34060 57400 34112 57452
rect 42800 57468 42852 57520
rect 52184 57468 52236 57520
rect 53104 57511 53156 57520
rect 53104 57477 53113 57511
rect 53113 57477 53147 57511
rect 53147 57477 53156 57511
rect 53104 57468 53156 57477
rect 56140 57468 56192 57520
rect 43812 57400 43864 57452
rect 44272 57443 44324 57452
rect 44272 57409 44281 57443
rect 44281 57409 44315 57443
rect 44315 57409 44324 57443
rect 44272 57400 44324 57409
rect 45652 57400 45704 57452
rect 51540 57400 51592 57452
rect 55220 57400 55272 57452
rect 56692 57400 56744 57452
rect 6920 57375 6972 57384
rect 6920 57341 6929 57375
rect 6929 57341 6963 57375
rect 6963 57341 6972 57375
rect 6920 57332 6972 57341
rect 10784 57332 10836 57384
rect 22468 57332 22520 57384
rect 25044 57375 25096 57384
rect 3884 57196 3936 57248
rect 8392 57196 8444 57248
rect 15476 57239 15528 57248
rect 15476 57205 15485 57239
rect 15485 57205 15519 57239
rect 15519 57205 15528 57239
rect 15476 57196 15528 57205
rect 19432 57239 19484 57248
rect 19432 57205 19441 57239
rect 19441 57205 19475 57239
rect 19475 57205 19484 57239
rect 19432 57196 19484 57205
rect 25044 57341 25053 57375
rect 25053 57341 25087 57375
rect 25087 57341 25096 57375
rect 25044 57332 25096 57341
rect 27528 57332 27580 57384
rect 32772 57332 32824 57384
rect 34704 57375 34756 57384
rect 34704 57341 34713 57375
rect 34713 57341 34747 57375
rect 34747 57341 34756 57375
rect 34704 57332 34756 57341
rect 48964 57375 49016 57384
rect 48964 57341 48973 57375
rect 48973 57341 49007 57375
rect 49007 57341 49016 57375
rect 48964 57332 49016 57341
rect 50160 57332 50212 57384
rect 50804 57375 50856 57384
rect 50804 57341 50813 57375
rect 50813 57341 50847 57375
rect 50847 57341 50856 57375
rect 50804 57332 50856 57341
rect 24584 57239 24636 57248
rect 24584 57205 24593 57239
rect 24593 57205 24627 57239
rect 24627 57205 24636 57239
rect 24584 57196 24636 57205
rect 29000 57239 29052 57248
rect 29000 57205 29009 57239
rect 29009 57205 29043 57239
rect 29043 57205 29052 57239
rect 29000 57196 29052 57205
rect 31208 57196 31260 57248
rect 36084 57239 36136 57248
rect 36084 57205 36093 57239
rect 36093 57205 36127 57239
rect 36127 57205 36136 57239
rect 36084 57196 36136 57205
rect 44548 57196 44600 57248
rect 45560 57196 45612 57248
rect 52184 57239 52236 57248
rect 52184 57205 52193 57239
rect 52193 57205 52227 57239
rect 52227 57205 52236 57239
rect 52184 57196 52236 57205
rect 57244 57196 57296 57248
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 5172 57035 5224 57044
rect 5172 57001 5181 57035
rect 5181 57001 5215 57035
rect 5215 57001 5224 57035
rect 5172 56992 5224 57001
rect 8300 57035 8352 57044
rect 8300 57001 8309 57035
rect 8309 57001 8343 57035
rect 8343 57001 8352 57035
rect 8300 56992 8352 57001
rect 12256 56992 12308 57044
rect 15844 57035 15896 57044
rect 15844 57001 15853 57035
rect 15853 57001 15887 57035
rect 15887 57001 15896 57035
rect 15844 56992 15896 57001
rect 18604 56992 18656 57044
rect 23848 57035 23900 57044
rect 23848 57001 23857 57035
rect 23857 57001 23891 57035
rect 23891 57001 23900 57035
rect 23848 56992 23900 57001
rect 25044 56992 25096 57044
rect 28908 57035 28960 57044
rect 28908 57001 28917 57035
rect 28917 57001 28951 57035
rect 28951 57001 28960 57035
rect 28908 56992 28960 57001
rect 32220 56992 32272 57044
rect 34060 56992 34112 57044
rect 38660 57035 38712 57044
rect 38660 57001 38669 57035
rect 38669 57001 38703 57035
rect 38703 57001 38712 57035
rect 38660 56992 38712 57001
rect 49424 56992 49476 57044
rect 52828 56992 52880 57044
rect 54852 56992 54904 57044
rect 56692 57035 56744 57044
rect 56692 57001 56701 57035
rect 56701 57001 56735 57035
rect 56735 57001 56744 57035
rect 56692 56992 56744 57001
rect 58440 56992 58492 57044
rect 8944 56899 8996 56908
rect 8944 56865 8953 56899
rect 8953 56865 8987 56899
rect 8987 56865 8996 56899
rect 8944 56856 8996 56865
rect 14096 56856 14148 56908
rect 19892 56899 19944 56908
rect 19892 56865 19901 56899
rect 19901 56865 19935 56899
rect 19935 56865 19944 56899
rect 19892 56856 19944 56865
rect 22468 56899 22520 56908
rect 22468 56865 22477 56899
rect 22477 56865 22511 56899
rect 22511 56865 22520 56899
rect 22468 56856 22520 56865
rect 32772 56899 32824 56908
rect 32772 56865 32781 56899
rect 32781 56865 32815 56899
rect 32815 56865 32824 56899
rect 32772 56856 32824 56865
rect 37280 56899 37332 56908
rect 37280 56865 37289 56899
rect 37289 56865 37323 56899
rect 37323 56865 37332 56899
rect 37280 56856 37332 56865
rect 40408 56856 40460 56908
rect 42708 56899 42760 56908
rect 42708 56865 42717 56899
rect 42717 56865 42751 56899
rect 42751 56865 42760 56899
rect 42708 56856 42760 56865
rect 44272 56856 44324 56908
rect 45008 56899 45060 56908
rect 45008 56865 45017 56899
rect 45017 56865 45051 56899
rect 45051 56865 45060 56899
rect 45008 56856 45060 56865
rect 50160 56856 50212 56908
rect 3884 56788 3936 56840
rect 6920 56831 6972 56840
rect 6920 56797 6929 56831
rect 6929 56797 6963 56831
rect 6963 56797 6972 56831
rect 6920 56788 6972 56797
rect 8300 56788 8352 56840
rect 11520 56831 11572 56840
rect 11520 56797 11529 56831
rect 11529 56797 11563 56831
rect 11563 56797 11572 56831
rect 11520 56788 11572 56797
rect 12900 56788 12952 56840
rect 15476 56788 15528 56840
rect 17868 56788 17920 56840
rect 20168 56831 20220 56840
rect 20168 56797 20202 56831
rect 20202 56797 20220 56831
rect 20168 56788 20220 56797
rect 24584 56788 24636 56840
rect 26976 56788 27028 56840
rect 27528 56831 27580 56840
rect 27528 56797 27537 56831
rect 27537 56797 27571 56831
rect 27571 56797 27580 56831
rect 27528 56788 27580 56797
rect 29000 56788 29052 56840
rect 31208 56831 31260 56840
rect 31208 56797 31242 56831
rect 31242 56797 31260 56831
rect 4988 56720 5040 56772
rect 10324 56695 10376 56704
rect 10324 56661 10333 56695
rect 10333 56661 10367 56695
rect 10367 56661 10376 56695
rect 10324 56652 10376 56661
rect 19248 56720 19300 56772
rect 27620 56720 27672 56772
rect 31208 56788 31260 56797
rect 32864 56788 32916 56840
rect 34704 56831 34756 56840
rect 34704 56797 34713 56831
rect 34713 56797 34747 56831
rect 34747 56797 34756 56831
rect 34704 56788 34756 56797
rect 36084 56788 36136 56840
rect 41144 56831 41196 56840
rect 41144 56797 41178 56831
rect 41178 56797 41196 56831
rect 41144 56788 41196 56797
rect 48504 56831 48556 56840
rect 48504 56797 48538 56831
rect 48538 56797 48556 56831
rect 32772 56720 32824 56772
rect 34244 56720 34296 56772
rect 39028 56720 39080 56772
rect 42800 56720 42852 56772
rect 46296 56720 46348 56772
rect 48504 56788 48556 56797
rect 48964 56720 49016 56772
rect 55220 56856 55272 56908
rect 52552 56788 52604 56840
rect 53380 56831 53432 56840
rect 53380 56797 53389 56831
rect 53389 56797 53423 56831
rect 53423 56797 53432 56831
rect 53380 56788 53432 56797
rect 52644 56720 52696 56772
rect 56876 56788 56928 56840
rect 57060 56788 57112 56840
rect 57244 56788 57296 56840
rect 55680 56720 55732 56772
rect 20996 56652 21048 56704
rect 21272 56695 21324 56704
rect 21272 56661 21281 56695
rect 21281 56661 21315 56695
rect 21315 56661 21324 56695
rect 21272 56652 21324 56661
rect 36084 56695 36136 56704
rect 36084 56661 36093 56695
rect 36093 56661 36127 56695
rect 36127 56661 36136 56695
rect 36084 56652 36136 56661
rect 42248 56695 42300 56704
rect 42248 56661 42257 56695
rect 42257 56661 42291 56695
rect 42291 56661 42300 56695
rect 42248 56652 42300 56661
rect 42340 56652 42392 56704
rect 46388 56695 46440 56704
rect 46388 56661 46397 56695
rect 46397 56661 46431 56695
rect 46431 56661 46440 56695
rect 46388 56652 46440 56661
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 4988 56491 5040 56500
rect 4988 56457 4997 56491
rect 4997 56457 5031 56491
rect 5031 56457 5040 56491
rect 4988 56448 5040 56457
rect 8300 56491 8352 56500
rect 8300 56457 8309 56491
rect 8309 56457 8343 56491
rect 8343 56457 8352 56491
rect 8300 56448 8352 56457
rect 8944 56448 8996 56500
rect 15936 56448 15988 56500
rect 23756 56491 23808 56500
rect 23756 56457 23765 56491
rect 23765 56457 23799 56491
rect 23799 56457 23808 56491
rect 23756 56448 23808 56457
rect 34244 56491 34296 56500
rect 34244 56457 34253 56491
rect 34253 56457 34287 56491
rect 34287 56457 34296 56491
rect 34244 56448 34296 56457
rect 39028 56491 39080 56500
rect 39028 56457 39037 56491
rect 39037 56457 39071 56491
rect 39071 56457 39080 56491
rect 39028 56448 39080 56457
rect 42800 56448 42852 56500
rect 43812 56491 43864 56500
rect 43812 56457 43821 56491
rect 43821 56457 43855 56491
rect 43855 56457 43864 56491
rect 43812 56448 43864 56457
rect 45652 56491 45704 56500
rect 45652 56457 45661 56491
rect 45661 56457 45695 56491
rect 45695 56457 45704 56491
rect 45652 56448 45704 56457
rect 50620 56448 50672 56500
rect 55680 56491 55732 56500
rect 55680 56457 55689 56491
rect 55689 56457 55723 56491
rect 55723 56457 55732 56491
rect 55680 56448 55732 56457
rect 5172 56312 5224 56364
rect 8208 56312 8260 56364
rect 10324 56380 10376 56432
rect 11520 56380 11572 56432
rect 14096 56380 14148 56432
rect 17316 56380 17368 56432
rect 19432 56380 19484 56432
rect 21272 56380 21324 56432
rect 23480 56380 23532 56432
rect 27620 56380 27672 56432
rect 36084 56380 36136 56432
rect 42248 56380 42300 56432
rect 44548 56423 44600 56432
rect 44548 56389 44582 56423
rect 44582 56389 44600 56423
rect 44548 56380 44600 56389
rect 49608 56380 49660 56432
rect 52184 56380 52236 56432
rect 15568 56312 15620 56364
rect 19984 56312 20036 56364
rect 22468 56312 22520 56364
rect 25044 56312 25096 56364
rect 28356 56312 28408 56364
rect 32864 56355 32916 56364
rect 32864 56321 32873 56355
rect 32873 56321 32907 56355
rect 32907 56321 32916 56355
rect 32864 56312 32916 56321
rect 6920 56287 6972 56296
rect 6920 56253 6929 56287
rect 6929 56253 6963 56287
rect 6963 56253 6972 56287
rect 6920 56244 6972 56253
rect 17868 56244 17920 56296
rect 19248 56176 19300 56228
rect 3884 56108 3936 56160
rect 10140 56151 10192 56160
rect 10140 56117 10149 56151
rect 10149 56117 10183 56151
rect 10183 56117 10192 56151
rect 10140 56108 10192 56117
rect 14188 56151 14240 56160
rect 14188 56117 14197 56151
rect 14197 56117 14231 56151
rect 14231 56117 14240 56151
rect 14188 56108 14240 56117
rect 16120 56151 16172 56160
rect 16120 56117 16129 56151
rect 16129 56117 16163 56151
rect 16163 56117 16172 56151
rect 16120 56108 16172 56117
rect 21272 56151 21324 56160
rect 21272 56117 21281 56151
rect 21281 56117 21315 56151
rect 21315 56117 21324 56151
rect 21272 56108 21324 56117
rect 21732 56108 21784 56160
rect 28264 56244 28316 56296
rect 34704 56287 34756 56296
rect 34704 56253 34713 56287
rect 34713 56253 34747 56287
rect 34747 56253 34756 56287
rect 34704 56244 34756 56253
rect 25596 56151 25648 56160
rect 25596 56117 25605 56151
rect 25605 56117 25639 56151
rect 25639 56117 25648 56151
rect 25596 56108 25648 56117
rect 29184 56108 29236 56160
rect 30380 56108 30432 56160
rect 37280 56312 37332 56364
rect 37648 56355 37700 56364
rect 37648 56321 37657 56355
rect 37657 56321 37691 56355
rect 37691 56321 37700 56355
rect 37648 56312 37700 56321
rect 39028 56312 39080 56364
rect 40408 56355 40460 56364
rect 40408 56321 40417 56355
rect 40417 56321 40451 56355
rect 40451 56321 40460 56355
rect 40408 56312 40460 56321
rect 41880 56312 41932 56364
rect 48964 56355 49016 56364
rect 48964 56321 48973 56355
rect 48973 56321 49007 56355
rect 49007 56321 49016 56355
rect 48964 56312 49016 56321
rect 35348 56108 35400 56160
rect 42800 56108 42852 56160
rect 53380 56244 53432 56296
rect 55128 56380 55180 56432
rect 55956 56312 56008 56364
rect 51908 56176 51960 56228
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 20628 55904 20680 55956
rect 28540 55947 28592 55956
rect 28540 55913 28549 55947
rect 28549 55913 28583 55947
rect 28583 55913 28592 55947
rect 28540 55904 28592 55913
rect 39028 55947 39080 55956
rect 39028 55913 39037 55947
rect 39037 55913 39071 55947
rect 39071 55913 39080 55947
rect 39028 55904 39080 55913
rect 42800 55904 42852 55956
rect 43076 55904 43128 55956
rect 46296 55904 46348 55956
rect 49332 55904 49384 55956
rect 56784 55904 56836 55956
rect 8944 55811 8996 55820
rect 8944 55777 8953 55811
rect 8953 55777 8987 55811
rect 8987 55777 8996 55811
rect 8944 55768 8996 55777
rect 14096 55768 14148 55820
rect 37648 55811 37700 55820
rect 37648 55777 37657 55811
rect 37657 55777 37691 55811
rect 37691 55777 37700 55811
rect 37648 55768 37700 55777
rect 45008 55811 45060 55820
rect 45008 55777 45017 55811
rect 45017 55777 45051 55811
rect 45051 55777 45060 55811
rect 45008 55768 45060 55777
rect 5540 55632 5592 55684
rect 8760 55632 8812 55684
rect 10140 55700 10192 55752
rect 11704 55700 11756 55752
rect 16120 55700 16172 55752
rect 9312 55632 9364 55684
rect 13728 55632 13780 55684
rect 18696 55700 18748 55752
rect 19984 55700 20036 55752
rect 21272 55700 21324 55752
rect 21732 55743 21784 55752
rect 21732 55709 21741 55743
rect 21741 55709 21775 55743
rect 21775 55709 21784 55743
rect 21732 55700 21784 55709
rect 21824 55700 21876 55752
rect 22468 55700 22520 55752
rect 23664 55700 23716 55752
rect 24400 55743 24452 55752
rect 24400 55709 24409 55743
rect 24409 55709 24443 55743
rect 24443 55709 24452 55743
rect 24400 55700 24452 55709
rect 26976 55700 27028 55752
rect 27252 55700 27304 55752
rect 32128 55743 32180 55752
rect 32128 55709 32137 55743
rect 32137 55709 32171 55743
rect 32171 55709 32180 55743
rect 32128 55700 32180 55709
rect 32772 55700 32824 55752
rect 35348 55700 35400 55752
rect 40132 55700 40184 55752
rect 42340 55700 42392 55752
rect 17868 55632 17920 55684
rect 23204 55632 23256 55684
rect 25412 55632 25464 55684
rect 33140 55632 33192 55684
rect 36728 55632 36780 55684
rect 6276 55607 6328 55616
rect 6276 55573 6285 55607
rect 6285 55573 6319 55607
rect 6319 55573 6328 55607
rect 6276 55564 6328 55573
rect 10324 55607 10376 55616
rect 10324 55573 10333 55607
rect 10333 55573 10367 55607
rect 10367 55573 10376 55607
rect 10324 55564 10376 55573
rect 14372 55564 14424 55616
rect 16028 55607 16080 55616
rect 16028 55573 16037 55607
rect 16037 55573 16071 55607
rect 16071 55573 16080 55607
rect 16028 55564 16080 55573
rect 18696 55607 18748 55616
rect 18696 55573 18705 55607
rect 18705 55573 18739 55607
rect 18739 55573 18748 55607
rect 18696 55564 18748 55573
rect 23848 55564 23900 55616
rect 28356 55564 28408 55616
rect 33508 55607 33560 55616
rect 33508 55573 33517 55607
rect 33517 55573 33551 55607
rect 33551 55573 33560 55607
rect 33508 55564 33560 55573
rect 41788 55632 41840 55684
rect 45560 55700 45612 55752
rect 48320 55743 48372 55752
rect 48320 55709 48354 55743
rect 48354 55709 48372 55743
rect 48320 55700 48372 55709
rect 50160 55743 50212 55752
rect 50160 55709 50169 55743
rect 50169 55709 50203 55743
rect 50203 55709 50212 55743
rect 50160 55700 50212 55709
rect 52736 55700 52788 55752
rect 53380 55743 53432 55752
rect 53380 55709 53389 55743
rect 53389 55709 53423 55743
rect 53423 55709 53432 55743
rect 53380 55700 53432 55709
rect 56600 55700 56652 55752
rect 51172 55632 51224 55684
rect 56140 55675 56192 55684
rect 56140 55641 56149 55675
rect 56149 55641 56183 55675
rect 56183 55641 56192 55675
rect 56140 55632 56192 55641
rect 41420 55607 41472 55616
rect 41420 55573 41429 55607
rect 41429 55573 41463 55607
rect 41463 55573 41472 55607
rect 41420 55564 41472 55573
rect 51540 55607 51592 55616
rect 51540 55573 51549 55607
rect 51549 55573 51583 55607
rect 51583 55573 51592 55607
rect 51540 55564 51592 55573
rect 57060 55564 57112 55616
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 5172 55403 5224 55412
rect 5172 55369 5181 55403
rect 5181 55369 5215 55403
rect 5215 55369 5224 55403
rect 5172 55360 5224 55369
rect 8208 55403 8260 55412
rect 8208 55369 8217 55403
rect 8217 55369 8251 55403
rect 8251 55369 8260 55403
rect 8208 55360 8260 55369
rect 13728 55403 13780 55412
rect 13728 55369 13737 55403
rect 13737 55369 13771 55403
rect 13771 55369 13780 55403
rect 13728 55360 13780 55369
rect 15568 55403 15620 55412
rect 15568 55369 15577 55403
rect 15577 55369 15611 55403
rect 15611 55369 15620 55403
rect 15568 55360 15620 55369
rect 19156 55403 19208 55412
rect 19156 55369 19165 55403
rect 19165 55369 19199 55403
rect 19199 55369 19208 55403
rect 19156 55360 19208 55369
rect 20996 55403 21048 55412
rect 20996 55369 21005 55403
rect 21005 55369 21039 55403
rect 21039 55369 21048 55403
rect 20996 55360 21048 55369
rect 23204 55403 23256 55412
rect 23204 55369 23213 55403
rect 23213 55369 23247 55403
rect 23247 55369 23256 55403
rect 23204 55360 23256 55369
rect 25044 55403 25096 55412
rect 25044 55369 25053 55403
rect 25053 55369 25087 55403
rect 25087 55369 25096 55403
rect 25044 55360 25096 55369
rect 29828 55360 29880 55412
rect 32404 55360 32456 55412
rect 36728 55403 36780 55412
rect 36728 55369 36737 55403
rect 36737 55369 36771 55403
rect 36771 55369 36780 55403
rect 36728 55360 36780 55369
rect 38936 55360 38988 55412
rect 41880 55403 41932 55412
rect 41880 55369 41889 55403
rect 41889 55369 41923 55403
rect 41923 55369 41932 55403
rect 41880 55360 41932 55369
rect 49700 55360 49752 55412
rect 52552 55360 52604 55412
rect 55956 55403 56008 55412
rect 55956 55369 55965 55403
rect 55965 55369 55999 55403
rect 55999 55369 56008 55403
rect 55956 55360 56008 55369
rect 8392 55292 8444 55344
rect 10324 55292 10376 55344
rect 14188 55292 14240 55344
rect 16028 55292 16080 55344
rect 18696 55292 18748 55344
rect 19340 55292 19392 55344
rect 19984 55292 20036 55344
rect 24400 55292 24452 55344
rect 28264 55292 28316 55344
rect 3884 55224 3936 55276
rect 6920 55224 6972 55276
rect 7932 55224 7984 55276
rect 17868 55224 17920 55276
rect 23112 55224 23164 55276
rect 23664 55267 23716 55276
rect 23664 55233 23673 55267
rect 23673 55233 23707 55267
rect 23707 55233 23716 55267
rect 23664 55224 23716 55233
rect 25044 55224 25096 55276
rect 28172 55224 28224 55276
rect 9312 55199 9364 55208
rect 9312 55165 9321 55199
rect 9321 55165 9355 55199
rect 9355 55165 9364 55199
rect 9312 55156 9364 55165
rect 14096 55156 14148 55208
rect 21824 55199 21876 55208
rect 21824 55165 21833 55199
rect 21833 55165 21867 55199
rect 21867 55165 21876 55199
rect 21824 55156 21876 55165
rect 7012 55020 7064 55072
rect 10692 55063 10744 55072
rect 10692 55029 10701 55063
rect 10701 55029 10735 55063
rect 10735 55029 10744 55063
rect 10692 55020 10744 55029
rect 26976 55020 27028 55072
rect 29276 55224 29328 55276
rect 30196 55224 30248 55276
rect 33416 55224 33468 55276
rect 35348 55267 35400 55276
rect 35348 55233 35357 55267
rect 35357 55233 35391 55267
rect 35391 55233 35400 55267
rect 35348 55224 35400 55233
rect 36636 55224 36688 55276
rect 40132 55292 40184 55344
rect 40500 55292 40552 55344
rect 41420 55292 41472 55344
rect 46388 55292 46440 55344
rect 41328 55224 41380 55276
rect 45192 55224 45244 55276
rect 29184 55199 29236 55208
rect 29184 55165 29193 55199
rect 29193 55165 29227 55199
rect 29227 55165 29236 55199
rect 29184 55156 29236 55165
rect 32128 55199 32180 55208
rect 32128 55165 32137 55199
rect 32137 55165 32171 55199
rect 32171 55165 32180 55199
rect 32128 55156 32180 55165
rect 40500 55199 40552 55208
rect 40500 55165 40509 55199
rect 40509 55165 40543 55199
rect 40543 55165 40552 55199
rect 40500 55156 40552 55165
rect 47584 55156 47636 55208
rect 49056 55224 49108 55276
rect 51540 55292 51592 55344
rect 50896 55224 50948 55276
rect 52644 55224 52696 55276
rect 29460 55020 29512 55072
rect 46480 55063 46532 55072
rect 46480 55029 46489 55063
rect 46489 55029 46523 55063
rect 46523 55029 46532 55063
rect 46480 55020 46532 55029
rect 51264 55063 51316 55072
rect 51264 55029 51273 55063
rect 51273 55029 51307 55063
rect 51307 55029 51316 55063
rect 51264 55020 51316 55029
rect 56140 55224 56192 55276
rect 55496 55020 55548 55072
rect 57060 55020 57112 55072
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 23112 54859 23164 54868
rect 23112 54825 23121 54859
rect 23121 54825 23155 54859
rect 23155 54825 23164 54859
rect 23112 54816 23164 54825
rect 25412 54816 25464 54868
rect 28172 54816 28224 54868
rect 36636 54859 36688 54868
rect 36636 54825 36645 54859
rect 36645 54825 36679 54859
rect 36679 54825 36688 54859
rect 36636 54816 36688 54825
rect 41328 54816 41380 54868
rect 49056 54859 49108 54868
rect 49056 54825 49065 54859
rect 49065 54825 49099 54859
rect 49099 54825 49108 54859
rect 49056 54816 49108 54825
rect 51172 54816 51224 54868
rect 6920 54723 6972 54732
rect 6920 54689 6929 54723
rect 6929 54689 6963 54723
rect 6963 54689 6972 54723
rect 14096 54723 14148 54732
rect 6920 54680 6972 54689
rect 14096 54689 14105 54723
rect 14105 54689 14139 54723
rect 14139 54689 14148 54723
rect 14096 54680 14148 54689
rect 21732 54723 21784 54732
rect 21732 54689 21741 54723
rect 21741 54689 21775 54723
rect 21775 54689 21784 54723
rect 21732 54680 21784 54689
rect 57060 54723 57112 54732
rect 57060 54689 57069 54723
rect 57069 54689 57103 54723
rect 57103 54689 57112 54723
rect 57060 54680 57112 54689
rect 3884 54612 3936 54664
rect 5632 54612 5684 54664
rect 6276 54612 6328 54664
rect 9496 54655 9548 54664
rect 9496 54621 9505 54655
rect 9505 54621 9539 54655
rect 9539 54621 9548 54655
rect 9496 54612 9548 54621
rect 10692 54612 10744 54664
rect 14372 54655 14424 54664
rect 14372 54621 14406 54655
rect 14406 54621 14424 54655
rect 14372 54612 14424 54621
rect 16580 54612 16632 54664
rect 20720 54612 20772 54664
rect 23664 54612 23716 54664
rect 24400 54655 24452 54664
rect 24400 54621 24409 54655
rect 24409 54621 24443 54655
rect 24443 54621 24452 54655
rect 24400 54612 24452 54621
rect 25596 54612 25648 54664
rect 26976 54612 27028 54664
rect 29460 54612 29512 54664
rect 37648 54612 37700 54664
rect 40592 54612 40644 54664
rect 45284 54612 45336 54664
rect 46480 54612 46532 54664
rect 47584 54612 47636 54664
rect 50160 54655 50212 54664
rect 50160 54621 50169 54655
rect 50169 54621 50203 54655
rect 50203 54621 50212 54655
rect 50160 54612 50212 54621
rect 51264 54612 51316 54664
rect 5816 54544 5868 54596
rect 7748 54544 7800 54596
rect 16212 54587 16264 54596
rect 16212 54553 16246 54587
rect 16246 54553 16264 54587
rect 16212 54544 16264 54553
rect 21088 54544 21140 54596
rect 23204 54544 23256 54596
rect 28356 54544 28408 54596
rect 29276 54544 29328 54596
rect 32496 54544 32548 54596
rect 33968 54587 34020 54596
rect 33968 54553 33977 54587
rect 33977 54553 34011 54587
rect 34011 54553 34020 54587
rect 33968 54544 34020 54553
rect 6460 54519 6512 54528
rect 6460 54485 6469 54519
rect 6469 54485 6503 54519
rect 6503 54485 6512 54519
rect 6460 54476 6512 54485
rect 7564 54476 7616 54528
rect 10876 54519 10928 54528
rect 10876 54485 10885 54519
rect 10885 54485 10919 54519
rect 10919 54485 10928 54519
rect 10876 54476 10928 54485
rect 15476 54519 15528 54528
rect 15476 54485 15485 54519
rect 15485 54485 15519 54519
rect 15519 54485 15528 54519
rect 15476 54476 15528 54485
rect 16672 54476 16724 54528
rect 21272 54519 21324 54528
rect 21272 54485 21281 54519
rect 21281 54485 21315 54519
rect 21315 54485 21324 54519
rect 21272 54476 21324 54485
rect 30932 54519 30984 54528
rect 30932 54485 30941 54519
rect 30941 54485 30975 54519
rect 30975 54485 30984 54519
rect 30932 54476 30984 54485
rect 39304 54544 39356 54596
rect 41788 54544 41840 54596
rect 44548 54544 44600 54596
rect 48964 54544 49016 54596
rect 52552 54612 52604 54664
rect 52736 54544 52788 54596
rect 57336 54587 57388 54596
rect 57336 54553 57370 54587
rect 57370 54553 57388 54587
rect 57336 54544 57388 54553
rect 44180 54476 44232 54528
rect 47216 54519 47268 54528
rect 47216 54485 47225 54519
rect 47225 54485 47259 54519
rect 47259 54485 47268 54519
rect 47216 54476 47268 54485
rect 52552 54476 52604 54528
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 7748 54315 7800 54324
rect 7748 54281 7757 54315
rect 7757 54281 7791 54315
rect 7791 54281 7800 54315
rect 7748 54272 7800 54281
rect 23204 54315 23256 54324
rect 23204 54281 23213 54315
rect 23213 54281 23247 54315
rect 23247 54281 23256 54315
rect 23204 54272 23256 54281
rect 25044 54315 25096 54324
rect 25044 54281 25053 54315
rect 25053 54281 25087 54315
rect 25087 54281 25096 54315
rect 25044 54272 25096 54281
rect 28356 54315 28408 54324
rect 28356 54281 28365 54315
rect 28365 54281 28399 54315
rect 28399 54281 28408 54315
rect 28356 54272 28408 54281
rect 30196 54315 30248 54324
rect 30196 54281 30205 54315
rect 30205 54281 30239 54315
rect 30239 54281 30248 54315
rect 30196 54272 30248 54281
rect 33416 54272 33468 54324
rect 48964 54315 49016 54324
rect 48964 54281 48973 54315
rect 48973 54281 49007 54315
rect 49007 54281 49016 54315
rect 48964 54272 49016 54281
rect 49700 54272 49752 54324
rect 50896 54315 50948 54324
rect 6460 54204 6512 54256
rect 10876 54204 10928 54256
rect 15476 54204 15528 54256
rect 16580 54204 16632 54256
rect 5356 54136 5408 54188
rect 6276 54136 6328 54188
rect 9312 54136 9364 54188
rect 11244 54136 11296 54188
rect 17868 54204 17920 54256
rect 20076 54204 20128 54256
rect 20444 54204 20496 54256
rect 21272 54204 21324 54256
rect 23940 54247 23992 54256
rect 23940 54213 23974 54247
rect 23974 54213 23992 54247
rect 23940 54204 23992 54213
rect 30932 54204 30984 54256
rect 17776 54136 17828 54188
rect 23664 54179 23716 54188
rect 23664 54145 23673 54179
rect 23673 54145 23707 54179
rect 23707 54145 23716 54179
rect 23664 54136 23716 54145
rect 26976 54179 27028 54188
rect 26976 54145 26985 54179
rect 26985 54145 27019 54179
rect 27019 54145 27028 54179
rect 26976 54136 27028 54145
rect 27252 54179 27304 54188
rect 27252 54145 27286 54179
rect 27286 54145 27304 54179
rect 27252 54136 27304 54145
rect 29552 54136 29604 54188
rect 32128 54179 32180 54188
rect 32128 54145 32137 54179
rect 32137 54145 32171 54179
rect 32171 54145 32180 54179
rect 33968 54204 34020 54256
rect 32128 54136 32180 54145
rect 32772 54136 32824 54188
rect 33508 54136 33560 54188
rect 40500 54204 40552 54256
rect 40040 54136 40092 54188
rect 42616 54136 42668 54188
rect 45284 54204 45336 54256
rect 47216 54204 47268 54256
rect 50896 54281 50905 54315
rect 50905 54281 50939 54315
rect 50939 54281 50948 54315
rect 50896 54272 50948 54281
rect 56140 54272 56192 54324
rect 44824 54136 44876 54188
rect 48964 54136 49016 54188
rect 50160 54136 50212 54188
rect 52460 54136 52512 54188
rect 55404 54136 55456 54188
rect 2872 54111 2924 54120
rect 2872 54077 2881 54111
rect 2881 54077 2915 54111
rect 2915 54077 2924 54111
rect 2872 54068 2924 54077
rect 4620 53932 4672 53984
rect 10968 53975 11020 53984
rect 10968 53941 10977 53975
rect 10977 53941 11011 53975
rect 11011 53941 11020 53975
rect 10968 53932 11020 53941
rect 20812 54068 20864 54120
rect 21824 54111 21876 54120
rect 21824 54077 21833 54111
rect 21833 54077 21867 54111
rect 21867 54077 21876 54111
rect 21824 54068 21876 54077
rect 33968 54111 34020 54120
rect 33968 54077 33977 54111
rect 33977 54077 34011 54111
rect 34011 54077 34020 54111
rect 33968 54068 34020 54077
rect 40500 54111 40552 54120
rect 40500 54077 40509 54111
rect 40509 54077 40543 54111
rect 40543 54077 40552 54111
rect 40500 54068 40552 54077
rect 45284 54068 45336 54120
rect 47584 54111 47636 54120
rect 47584 54077 47593 54111
rect 47593 54077 47627 54111
rect 47627 54077 47636 54111
rect 47584 54068 47636 54077
rect 52736 54111 52788 54120
rect 52736 54077 52745 54111
rect 52745 54077 52779 54111
rect 52779 54077 52788 54111
rect 52736 54068 52788 54077
rect 55496 54111 55548 54120
rect 55496 54077 55505 54111
rect 55505 54077 55539 54111
rect 55539 54077 55548 54111
rect 55496 54068 55548 54077
rect 11704 53932 11756 53984
rect 12900 53975 12952 53984
rect 12900 53941 12909 53975
rect 12909 53941 12943 53975
rect 12943 53941 12952 53975
rect 12900 53932 12952 53941
rect 16028 53975 16080 53984
rect 16028 53941 16037 53975
rect 16037 53941 16071 53975
rect 16071 53941 16080 53975
rect 16028 53932 16080 53941
rect 18052 53975 18104 53984
rect 18052 53941 18061 53975
rect 18061 53941 18095 53975
rect 18095 53941 18104 53975
rect 18052 53932 18104 53941
rect 33232 53932 33284 53984
rect 38660 53932 38712 53984
rect 41420 53932 41472 53984
rect 45192 53975 45244 53984
rect 45192 53941 45201 53975
rect 45201 53941 45235 53975
rect 45235 53941 45244 53975
rect 45192 53932 45244 53941
rect 47032 53975 47084 53984
rect 47032 53941 47041 53975
rect 47041 53941 47075 53975
rect 47075 53941 47084 53975
rect 47032 53932 47084 53941
rect 52920 53932 52972 53984
rect 54116 53975 54168 53984
rect 54116 53941 54125 53975
rect 54125 53941 54159 53975
rect 54159 53941 54168 53975
rect 54116 53932 54168 53941
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 11244 53771 11296 53780
rect 11244 53737 11253 53771
rect 11253 53737 11287 53771
rect 11287 53737 11296 53771
rect 11244 53728 11296 53737
rect 16212 53728 16264 53780
rect 17776 53771 17828 53780
rect 17776 53737 17785 53771
rect 17785 53737 17819 53771
rect 17819 53737 17828 53771
rect 17776 53728 17828 53737
rect 21088 53728 21140 53780
rect 27252 53728 27304 53780
rect 32772 53771 32824 53780
rect 32772 53737 32781 53771
rect 32781 53737 32815 53771
rect 32815 53737 32824 53771
rect 32772 53728 32824 53737
rect 39304 53771 39356 53780
rect 39304 53737 39313 53771
rect 39313 53737 39347 53771
rect 39347 53737 39356 53771
rect 39304 53728 39356 53737
rect 42616 53771 42668 53780
rect 42616 53737 42625 53771
rect 42625 53737 42659 53771
rect 42659 53737 42668 53771
rect 42616 53728 42668 53737
rect 52460 53771 52512 53780
rect 52460 53737 52469 53771
rect 52469 53737 52503 53771
rect 52503 53737 52512 53771
rect 52460 53728 52512 53737
rect 2872 53592 2924 53644
rect 3792 53635 3844 53644
rect 3792 53601 3801 53635
rect 3801 53601 3835 53635
rect 3835 53601 3844 53635
rect 3792 53592 3844 53601
rect 5632 53635 5684 53644
rect 5632 53601 5641 53635
rect 5641 53601 5675 53635
rect 5675 53601 5684 53635
rect 5632 53592 5684 53601
rect 43076 53635 43128 53644
rect 4620 53524 4672 53576
rect 9496 53524 9548 53576
rect 10968 53524 11020 53576
rect 11704 53567 11756 53576
rect 11704 53533 11713 53567
rect 11713 53533 11747 53567
rect 11747 53533 11756 53567
rect 11704 53524 11756 53533
rect 12900 53524 12952 53576
rect 43076 53601 43085 53635
rect 43085 53601 43119 53635
rect 43119 53601 43128 53635
rect 43076 53592 43128 53601
rect 50160 53592 50212 53644
rect 16028 53524 16080 53576
rect 16672 53567 16724 53576
rect 16672 53533 16706 53567
rect 16706 53533 16724 53567
rect 14648 53456 14700 53508
rect 16672 53524 16724 53533
rect 17868 53524 17920 53576
rect 18512 53524 18564 53576
rect 20812 53524 20864 53576
rect 21824 53524 21876 53576
rect 25044 53524 25096 53576
rect 26976 53524 27028 53576
rect 29552 53567 29604 53576
rect 29552 53533 29561 53567
rect 29561 53533 29595 53567
rect 29595 53533 29604 53567
rect 29552 53524 29604 53533
rect 29828 53567 29880 53576
rect 29828 53533 29862 53567
rect 29862 53533 29880 53567
rect 29828 53524 29880 53533
rect 19984 53456 20036 53508
rect 20720 53456 20772 53508
rect 26424 53456 26476 53508
rect 32128 53524 32180 53576
rect 34704 53567 34756 53576
rect 34704 53533 34713 53567
rect 34713 53533 34747 53567
rect 34747 53533 34756 53567
rect 34704 53524 34756 53533
rect 37924 53567 37976 53576
rect 37924 53533 37933 53567
rect 37933 53533 37967 53567
rect 37967 53533 37976 53567
rect 37924 53524 37976 53533
rect 38660 53524 38712 53576
rect 40500 53524 40552 53576
rect 45284 53567 45336 53576
rect 45284 53533 45293 53567
rect 45293 53533 45327 53567
rect 45327 53533 45336 53567
rect 45284 53524 45336 53533
rect 47032 53524 47084 53576
rect 47124 53567 47176 53576
rect 47124 53533 47133 53567
rect 47133 53533 47167 53567
rect 47167 53533 47176 53567
rect 47124 53524 47176 53533
rect 52552 53524 52604 53576
rect 52920 53567 52972 53576
rect 52920 53533 52929 53567
rect 52929 53533 52963 53567
rect 52963 53533 52972 53567
rect 52920 53524 52972 53533
rect 54116 53524 54168 53576
rect 55956 53524 56008 53576
rect 30840 53456 30892 53508
rect 34060 53456 34112 53508
rect 41880 53456 41932 53508
rect 44364 53456 44416 53508
rect 57704 53456 57756 53508
rect 7012 53431 7064 53440
rect 7012 53397 7021 53431
rect 7021 53397 7055 53431
rect 7055 53397 7064 53431
rect 7012 53388 7064 53397
rect 13084 53431 13136 53440
rect 13084 53397 13093 53431
rect 13093 53397 13127 53431
rect 13127 53397 13136 53431
rect 13084 53388 13136 53397
rect 20628 53431 20680 53440
rect 20628 53397 20637 53431
rect 20637 53397 20671 53431
rect 20671 53397 20680 53431
rect 20628 53388 20680 53397
rect 30932 53431 30984 53440
rect 30932 53397 30941 53431
rect 30941 53397 30975 53431
rect 30975 53397 30984 53431
rect 30932 53388 30984 53397
rect 36084 53431 36136 53440
rect 36084 53397 36093 53431
rect 36093 53397 36127 53431
rect 36127 53397 36136 53431
rect 36084 53388 36136 53397
rect 44456 53431 44508 53440
rect 44456 53397 44465 53431
rect 44465 53397 44499 53431
rect 44499 53397 44508 53431
rect 44456 53388 44508 53397
rect 46664 53431 46716 53440
rect 46664 53397 46673 53431
rect 46673 53397 46707 53431
rect 46707 53397 46716 53431
rect 46664 53388 46716 53397
rect 47584 53388 47636 53440
rect 51356 53388 51408 53440
rect 58164 53431 58216 53440
rect 58164 53397 58173 53431
rect 58173 53397 58207 53431
rect 58207 53397 58216 53431
rect 58164 53388 58216 53397
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 5356 53227 5408 53236
rect 2872 53116 2924 53168
rect 5356 53193 5365 53227
rect 5365 53193 5399 53227
rect 5399 53193 5408 53227
rect 5356 53184 5408 53193
rect 7932 53227 7984 53236
rect 7932 53193 7941 53227
rect 7941 53193 7975 53227
rect 7975 53193 7984 53227
rect 7932 53184 7984 53193
rect 19984 53184 20036 53236
rect 26424 53227 26476 53236
rect 26424 53193 26433 53227
rect 26433 53193 26467 53227
rect 26467 53193 26476 53227
rect 26424 53184 26476 53193
rect 3240 53048 3292 53100
rect 7564 53116 7616 53168
rect 13360 53116 13412 53168
rect 13820 53116 13872 53168
rect 14648 53159 14700 53168
rect 14648 53125 14657 53159
rect 14657 53125 14691 53159
rect 14691 53125 14700 53159
rect 14648 53116 14700 53125
rect 18052 53116 18104 53168
rect 30380 53184 30432 53236
rect 30840 53227 30892 53236
rect 30840 53193 30849 53227
rect 30849 53193 30883 53227
rect 30883 53193 30892 53227
rect 30840 53184 30892 53193
rect 33140 53184 33192 53236
rect 40040 53227 40092 53236
rect 40040 53193 40049 53227
rect 40049 53193 40083 53227
rect 40083 53193 40092 53227
rect 40040 53184 40092 53193
rect 41880 53227 41932 53236
rect 41880 53193 41889 53227
rect 41889 53193 41923 53227
rect 41923 53193 41932 53227
rect 41880 53184 41932 53193
rect 44824 53227 44876 53236
rect 44824 53193 44833 53227
rect 44833 53193 44867 53227
rect 44867 53193 44876 53227
rect 44824 53184 44876 53193
rect 48964 53227 49016 53236
rect 48964 53193 48973 53227
rect 48973 53193 49007 53227
rect 49007 53193 49016 53227
rect 48964 53184 49016 53193
rect 55404 53184 55456 53236
rect 57336 53227 57388 53236
rect 57336 53193 57345 53227
rect 57345 53193 57379 53227
rect 57379 53193 57388 53227
rect 57336 53184 57388 53193
rect 30932 53116 30984 53168
rect 32404 53159 32456 53168
rect 32404 53125 32438 53159
rect 32438 53125 32456 53159
rect 32404 53116 32456 53125
rect 36084 53116 36136 53168
rect 38936 53159 38988 53168
rect 38936 53125 38970 53159
rect 38970 53125 38988 53159
rect 38936 53116 38988 53125
rect 44180 53116 44232 53168
rect 46664 53116 46716 53168
rect 58164 53116 58216 53168
rect 6276 53048 6328 53100
rect 18512 53091 18564 53100
rect 18512 53057 18521 53091
rect 18521 53057 18555 53091
rect 18555 53057 18564 53091
rect 18512 53048 18564 53057
rect 18604 53048 18656 53100
rect 24860 53048 24912 53100
rect 25044 53091 25096 53100
rect 25044 53057 25053 53091
rect 25053 53057 25087 53091
rect 25087 53057 25096 53091
rect 25044 53048 25096 53057
rect 26240 53048 26292 53100
rect 29460 53091 29512 53100
rect 29460 53057 29469 53091
rect 29469 53057 29503 53091
rect 29503 53057 29512 53091
rect 29460 53048 29512 53057
rect 33968 53091 34020 53100
rect 33968 53057 33977 53091
rect 33977 53057 34011 53091
rect 34011 53057 34020 53091
rect 33968 53048 34020 53057
rect 34704 53048 34756 53100
rect 37924 53048 37976 53100
rect 40500 53091 40552 53100
rect 40500 53057 40509 53091
rect 40509 53057 40543 53091
rect 40543 53057 40552 53091
rect 40500 53048 40552 53057
rect 45284 53023 45336 53032
rect 17408 52844 17460 52896
rect 26792 52844 26844 52896
rect 35348 52887 35400 52896
rect 35348 52853 35357 52887
rect 35357 52853 35391 52887
rect 35391 52853 35400 52887
rect 35348 52844 35400 52853
rect 43076 52844 43128 52896
rect 45284 52989 45293 53023
rect 45293 52989 45327 53023
rect 45327 52989 45336 53023
rect 45284 52980 45336 52989
rect 48320 53048 48372 53100
rect 52920 53048 52972 53100
rect 54760 53048 54812 53100
rect 55956 53091 56008 53100
rect 55956 53057 55965 53091
rect 55965 53057 55999 53091
rect 55999 53057 56008 53091
rect 55956 53048 56008 53057
rect 47584 53023 47636 53032
rect 47584 52989 47593 53023
rect 47593 52989 47627 53023
rect 47627 52989 47636 53023
rect 47584 52980 47636 52989
rect 45468 52844 45520 52896
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 3240 52683 3292 52692
rect 3240 52649 3249 52683
rect 3249 52649 3283 52683
rect 3283 52649 3292 52683
rect 3240 52640 3292 52649
rect 5816 52683 5868 52692
rect 5816 52649 5825 52683
rect 5825 52649 5859 52683
rect 5859 52649 5868 52683
rect 5816 52640 5868 52649
rect 9496 52640 9548 52692
rect 18604 52640 18656 52692
rect 26240 52683 26292 52692
rect 26240 52649 26249 52683
rect 26249 52649 26283 52683
rect 26283 52649 26292 52683
rect 34060 52683 34112 52692
rect 26240 52640 26292 52649
rect 34060 52649 34069 52683
rect 34069 52649 34103 52683
rect 34103 52649 34112 52683
rect 34060 52640 34112 52649
rect 41788 52683 41840 52692
rect 41788 52649 41797 52683
rect 41797 52649 41831 52683
rect 41831 52649 41840 52683
rect 41788 52640 41840 52649
rect 44364 52640 44416 52692
rect 48320 52683 48372 52692
rect 48320 52649 48329 52683
rect 48329 52649 48363 52683
rect 48363 52649 48372 52683
rect 48320 52640 48372 52649
rect 54760 52683 54812 52692
rect 54760 52649 54769 52683
rect 54769 52649 54803 52683
rect 54803 52649 54812 52683
rect 54760 52640 54812 52649
rect 57704 52683 57756 52692
rect 57704 52649 57713 52683
rect 57713 52649 57747 52683
rect 57747 52649 57756 52683
rect 57704 52640 57756 52649
rect 10140 52572 10192 52624
rect 23020 52572 23072 52624
rect 24860 52547 24912 52556
rect 24860 52513 24869 52547
rect 24869 52513 24903 52547
rect 24903 52513 24912 52547
rect 24860 52504 24912 52513
rect 43076 52547 43128 52556
rect 43076 52513 43085 52547
rect 43085 52513 43119 52547
rect 43119 52513 43128 52547
rect 43076 52504 43128 52513
rect 55956 52504 56008 52556
rect 1584 52436 1636 52488
rect 3424 52436 3476 52488
rect 7012 52436 7064 52488
rect 10968 52436 11020 52488
rect 11612 52436 11664 52488
rect 13084 52436 13136 52488
rect 14096 52479 14148 52488
rect 14096 52445 14105 52479
rect 14105 52445 14139 52479
rect 14139 52445 14148 52479
rect 14096 52436 14148 52445
rect 14648 52436 14700 52488
rect 16672 52436 16724 52488
rect 17408 52479 17460 52488
rect 17408 52445 17442 52479
rect 17442 52445 17460 52479
rect 17408 52436 17460 52445
rect 4620 52368 4672 52420
rect 13820 52368 13872 52420
rect 20628 52436 20680 52488
rect 21732 52436 21784 52488
rect 23756 52436 23808 52488
rect 25688 52436 25740 52488
rect 20812 52368 20864 52420
rect 24860 52368 24912 52420
rect 26792 52436 26844 52488
rect 33232 52436 33284 52488
rect 39856 52436 39908 52488
rect 41420 52436 41472 52488
rect 45192 52436 45244 52488
rect 45468 52436 45520 52488
rect 48964 52436 49016 52488
rect 51356 52479 51408 52488
rect 47584 52368 47636 52420
rect 51356 52445 51390 52479
rect 51390 52445 51408 52479
rect 51356 52436 51408 52445
rect 53104 52436 53156 52488
rect 54484 52436 54536 52488
rect 57336 52368 57388 52420
rect 12900 52343 12952 52352
rect 12900 52309 12909 52343
rect 12909 52309 12943 52343
rect 12943 52309 12952 52343
rect 12900 52300 12952 52309
rect 15200 52300 15252 52352
rect 21364 52343 21416 52352
rect 21364 52309 21373 52343
rect 21373 52309 21407 52343
rect 21407 52309 21416 52343
rect 21364 52300 21416 52309
rect 26976 52300 27028 52352
rect 28080 52343 28132 52352
rect 28080 52309 28089 52343
rect 28089 52309 28123 52343
rect 28123 52309 28132 52343
rect 28080 52300 28132 52309
rect 33232 52300 33284 52352
rect 52460 52343 52512 52352
rect 52460 52309 52469 52343
rect 52469 52309 52503 52343
rect 52503 52309 52512 52343
rect 52460 52300 52512 52309
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 3424 52139 3476 52148
rect 3424 52105 3433 52139
rect 3433 52105 3467 52139
rect 3467 52105 3476 52139
rect 3424 52096 3476 52105
rect 10968 52139 11020 52148
rect 10968 52105 10977 52139
rect 10977 52105 11011 52139
rect 11011 52105 11020 52139
rect 10968 52096 11020 52105
rect 13360 52139 13412 52148
rect 13360 52105 13369 52139
rect 13369 52105 13403 52139
rect 13403 52105 13412 52139
rect 13360 52096 13412 52105
rect 20720 52096 20772 52148
rect 40316 52139 40368 52148
rect 40316 52105 40325 52139
rect 40325 52105 40359 52139
rect 40359 52105 40368 52139
rect 40316 52096 40368 52105
rect 41696 52096 41748 52148
rect 43076 52096 43128 52148
rect 44548 52139 44600 52148
rect 44548 52105 44557 52139
rect 44557 52105 44591 52139
rect 44591 52105 44600 52139
rect 44548 52096 44600 52105
rect 47124 52096 47176 52148
rect 48964 52139 49016 52148
rect 48964 52105 48973 52139
rect 48973 52105 49007 52139
rect 49007 52105 49016 52139
rect 48964 52096 49016 52105
rect 54484 52139 54536 52148
rect 54484 52105 54493 52139
rect 54493 52105 54527 52139
rect 54527 52105 54536 52139
rect 54484 52096 54536 52105
rect 57336 52139 57388 52148
rect 57336 52105 57345 52139
rect 57345 52105 57379 52139
rect 57379 52105 57388 52139
rect 57336 52096 57388 52105
rect 3240 51960 3292 52012
rect 7012 52028 7064 52080
rect 8392 51960 8444 52012
rect 10968 51960 11020 52012
rect 12900 52028 12952 52080
rect 21364 52028 21416 52080
rect 28080 52028 28132 52080
rect 35348 52028 35400 52080
rect 44456 52028 44508 52080
rect 52460 52028 52512 52080
rect 11612 51960 11664 52012
rect 1584 51892 1636 51944
rect 13636 51960 13688 52012
rect 16672 52003 16724 52012
rect 16672 51969 16681 52003
rect 16681 51969 16715 52003
rect 16715 51969 16724 52003
rect 16672 51960 16724 51969
rect 18052 51960 18104 52012
rect 23204 51960 23256 52012
rect 24492 51960 24544 52012
rect 28908 51960 28960 52012
rect 29920 51960 29972 52012
rect 33232 51960 33284 52012
rect 34704 51960 34756 52012
rect 35992 51960 36044 52012
rect 39948 51960 40000 52012
rect 40960 51960 41012 52012
rect 49056 51960 49108 52012
rect 53104 52003 53156 52012
rect 53104 51969 53113 52003
rect 53113 51969 53147 52003
rect 53147 51969 53156 52003
rect 53104 51960 53156 51969
rect 54300 51960 54352 52012
rect 55956 52003 56008 52012
rect 55956 51969 55965 52003
rect 55965 51969 55999 52003
rect 55999 51969 56008 52003
rect 55956 51960 56008 51969
rect 57152 51960 57204 52012
rect 14004 51892 14056 51944
rect 14096 51935 14148 51944
rect 14096 51901 14105 51935
rect 14105 51901 14139 51935
rect 14139 51901 14148 51935
rect 19248 51935 19300 51944
rect 14096 51892 14148 51901
rect 19248 51901 19257 51935
rect 19257 51901 19291 51935
rect 19291 51901 19300 51935
rect 19248 51892 19300 51901
rect 21824 51935 21876 51944
rect 21824 51901 21833 51935
rect 21833 51901 21867 51935
rect 21867 51901 21876 51935
rect 21824 51892 21876 51901
rect 23664 51935 23716 51944
rect 23664 51901 23673 51935
rect 23673 51901 23707 51935
rect 23707 51901 23716 51935
rect 23664 51892 23716 51901
rect 26976 51935 27028 51944
rect 26976 51901 26985 51935
rect 26985 51901 27019 51935
rect 27019 51901 27028 51935
rect 26976 51892 27028 51901
rect 37188 51892 37240 51944
rect 43168 51935 43220 51944
rect 43168 51901 43177 51935
rect 43177 51901 43211 51935
rect 43211 51901 43220 51935
rect 43168 51892 43220 51901
rect 47584 51935 47636 51944
rect 47584 51901 47593 51935
rect 47593 51901 47627 51935
rect 47627 51901 47636 51935
rect 47584 51892 47636 51901
rect 48780 51892 48832 51944
rect 13820 51824 13872 51876
rect 7932 51799 7984 51808
rect 7932 51765 7941 51799
rect 7941 51765 7975 51799
rect 7975 51765 7984 51799
rect 7932 51756 7984 51765
rect 15476 51799 15528 51808
rect 15476 51765 15485 51799
rect 15485 51765 15519 51799
rect 15519 51765 15528 51799
rect 15476 51756 15528 51765
rect 17776 51756 17828 51808
rect 23940 51756 23992 51808
rect 24952 51756 25004 51808
rect 28356 51799 28408 51808
rect 28356 51765 28365 51799
rect 28365 51765 28399 51799
rect 28399 51765 28408 51799
rect 28356 51756 28408 51765
rect 30196 51799 30248 51808
rect 30196 51765 30205 51799
rect 30205 51765 30239 51799
rect 30239 51765 30248 51799
rect 30196 51756 30248 51765
rect 33048 51756 33100 51808
rect 36636 51756 36688 51808
rect 40132 51756 40184 51808
rect 52184 51799 52236 51808
rect 52184 51765 52193 51799
rect 52193 51765 52227 51799
rect 52227 51765 52236 51799
rect 52184 51756 52236 51765
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 3240 51595 3292 51604
rect 3240 51561 3249 51595
rect 3249 51561 3283 51595
rect 3283 51561 3292 51595
rect 3240 51552 3292 51561
rect 8392 51595 8444 51604
rect 8392 51561 8401 51595
rect 8401 51561 8435 51595
rect 8435 51561 8444 51595
rect 8392 51552 8444 51561
rect 13636 51552 13688 51604
rect 14004 51552 14056 51604
rect 19340 51484 19392 51536
rect 20076 51484 20128 51536
rect 14096 51459 14148 51468
rect 1584 51348 1636 51400
rect 4436 51348 4488 51400
rect 5172 51391 5224 51400
rect 5172 51357 5181 51391
rect 5181 51357 5215 51391
rect 5215 51357 5224 51391
rect 5172 51348 5224 51357
rect 7012 51391 7064 51400
rect 7012 51357 7021 51391
rect 7021 51357 7055 51391
rect 7055 51357 7064 51391
rect 7012 51348 7064 51357
rect 11704 51348 11756 51400
rect 14096 51425 14105 51459
rect 14105 51425 14139 51459
rect 14139 51425 14148 51459
rect 14096 51416 14148 51425
rect 15476 51348 15528 51400
rect 16672 51348 16724 51400
rect 20720 51484 20772 51536
rect 24768 51552 24820 51604
rect 49056 51595 49108 51604
rect 49056 51561 49065 51595
rect 49065 51561 49099 51595
rect 49099 51561 49108 51595
rect 49056 51552 49108 51561
rect 54300 51595 54352 51604
rect 54300 51561 54309 51595
rect 54309 51561 54343 51595
rect 54343 51561 54352 51595
rect 54300 51552 54352 51561
rect 55956 51552 56008 51604
rect 39856 51459 39908 51468
rect 39856 51425 39865 51459
rect 39865 51425 39899 51459
rect 39899 51425 39908 51459
rect 39856 51416 39908 51425
rect 45560 51416 45612 51468
rect 20812 51348 20864 51400
rect 21824 51348 21876 51400
rect 25780 51348 25832 51400
rect 27620 51348 27672 51400
rect 30104 51348 30156 51400
rect 33048 51391 33100 51400
rect 33048 51357 33082 51391
rect 33082 51357 33100 51391
rect 3424 51280 3476 51332
rect 6184 51280 6236 51332
rect 9128 51280 9180 51332
rect 12164 51280 12216 51332
rect 15200 51280 15252 51332
rect 15568 51280 15620 51332
rect 21272 51280 21324 51332
rect 25044 51280 25096 51332
rect 30472 51280 30524 51332
rect 33048 51348 33100 51357
rect 33232 51280 33284 51332
rect 36544 51391 36596 51400
rect 36544 51357 36553 51391
rect 36553 51357 36587 51391
rect 36587 51357 36596 51391
rect 36544 51348 36596 51357
rect 37188 51348 37240 51400
rect 47584 51348 47636 51400
rect 50620 51348 50672 51400
rect 52184 51348 52236 51400
rect 53012 51348 53064 51400
rect 58532 51348 58584 51400
rect 34612 51280 34664 51332
rect 37832 51280 37884 51332
rect 41144 51280 41196 51332
rect 47768 51280 47820 51332
rect 48964 51280 49016 51332
rect 56048 51280 56100 51332
rect 6552 51255 6604 51264
rect 6552 51221 6561 51255
rect 6561 51221 6595 51255
rect 6595 51221 6604 51255
rect 6552 51212 6604 51221
rect 11612 51255 11664 51264
rect 11612 51221 11621 51255
rect 11621 51221 11655 51255
rect 11655 51221 11664 51255
rect 11612 51212 11664 51221
rect 15476 51255 15528 51264
rect 15476 51221 15485 51255
rect 15485 51221 15519 51255
rect 15519 51221 15528 51255
rect 15476 51212 15528 51221
rect 17316 51255 17368 51264
rect 17316 51221 17325 51255
rect 17325 51221 17359 51255
rect 17359 51221 17368 51255
rect 17316 51212 17368 51221
rect 20076 51212 20128 51264
rect 21180 51212 21232 51264
rect 22100 51255 22152 51264
rect 22100 51221 22109 51255
rect 22109 51221 22143 51255
rect 22143 51221 22152 51255
rect 22100 51212 22152 51221
rect 23480 51212 23532 51264
rect 28908 51212 28960 51264
rect 30288 51212 30340 51264
rect 34152 51255 34204 51264
rect 34152 51221 34161 51255
rect 34161 51221 34195 51255
rect 34195 51221 34204 51255
rect 34152 51212 34204 51221
rect 36084 51255 36136 51264
rect 36084 51221 36093 51255
rect 36093 51221 36127 51255
rect 36127 51221 36136 51255
rect 36084 51212 36136 51221
rect 37924 51255 37976 51264
rect 37924 51221 37933 51255
rect 37933 51221 37967 51255
rect 37967 51221 37976 51255
rect 37924 51212 37976 51221
rect 41788 51212 41840 51264
rect 47216 51255 47268 51264
rect 47216 51221 47225 51255
rect 47225 51221 47259 51255
rect 47259 51221 47268 51255
rect 47216 51212 47268 51221
rect 52276 51255 52328 51264
rect 52276 51221 52285 51255
rect 52285 51221 52319 51255
rect 52319 51221 52328 51255
rect 52276 51212 52328 51221
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 3424 51051 3476 51060
rect 3424 51017 3433 51051
rect 3433 51017 3467 51051
rect 3467 51017 3476 51051
rect 3424 51008 3476 51017
rect 9128 51051 9180 51060
rect 9128 51017 9137 51051
rect 9137 51017 9171 51051
rect 9171 51017 9180 51051
rect 9128 51008 9180 51017
rect 10968 51051 11020 51060
rect 10968 51017 10977 51051
rect 10977 51017 11011 51051
rect 11011 51017 11020 51051
rect 10968 51008 11020 51017
rect 12164 51008 12216 51060
rect 18052 51051 18104 51060
rect 18052 51017 18061 51051
rect 18061 51017 18095 51051
rect 18095 51017 18104 51051
rect 18052 51008 18104 51017
rect 21272 51051 21324 51060
rect 21272 51017 21281 51051
rect 21281 51017 21315 51051
rect 21315 51017 21324 51051
rect 21272 51008 21324 51017
rect 23204 51051 23256 51060
rect 23204 51017 23213 51051
rect 23213 51017 23247 51051
rect 23247 51017 23256 51051
rect 23204 51008 23256 51017
rect 25044 51051 25096 51060
rect 25044 51017 25053 51051
rect 25053 51017 25087 51051
rect 25087 51017 25096 51051
rect 25044 51008 25096 51017
rect 34612 51051 34664 51060
rect 34612 51017 34621 51051
rect 34621 51017 34655 51051
rect 34655 51017 34664 51051
rect 34612 51008 34664 51017
rect 39948 51008 40000 51060
rect 48964 51051 49016 51060
rect 48964 51017 48973 51051
rect 48973 51017 49007 51051
rect 49007 51017 49016 51051
rect 48964 51008 49016 51017
rect 57152 51051 57204 51060
rect 57152 51017 57161 51051
rect 57161 51017 57195 51051
rect 57195 51017 57204 51051
rect 57152 51008 57204 51017
rect 6552 50940 6604 50992
rect 11612 50940 11664 50992
rect 15476 50940 15528 50992
rect 22100 50983 22152 50992
rect 22100 50949 22134 50983
rect 22134 50949 22152 50983
rect 22100 50940 22152 50949
rect 23940 50983 23992 50992
rect 23940 50949 23974 50983
rect 23974 50949 23992 50983
rect 23940 50940 23992 50949
rect 28356 50940 28408 50992
rect 3240 50872 3292 50924
rect 4436 50915 4488 50924
rect 4436 50881 4445 50915
rect 4445 50881 4479 50915
rect 4479 50881 4488 50915
rect 4436 50872 4488 50881
rect 10140 50872 10192 50924
rect 11244 50872 11296 50924
rect 17408 50872 17460 50924
rect 23112 50872 23164 50924
rect 23664 50915 23716 50924
rect 23664 50881 23673 50915
rect 23673 50881 23707 50915
rect 23707 50881 23716 50915
rect 23664 50872 23716 50881
rect 1584 50804 1636 50856
rect 11704 50847 11756 50856
rect 5816 50711 5868 50720
rect 5816 50677 5825 50711
rect 5825 50677 5859 50711
rect 5859 50677 5868 50711
rect 5816 50668 5868 50677
rect 8116 50668 8168 50720
rect 11704 50813 11713 50847
rect 11713 50813 11747 50847
rect 11747 50813 11756 50847
rect 11704 50804 11756 50813
rect 14096 50847 14148 50856
rect 14096 50813 14105 50847
rect 14105 50813 14139 50847
rect 14139 50813 14148 50847
rect 14096 50804 14148 50813
rect 16672 50847 16724 50856
rect 16672 50813 16681 50847
rect 16681 50813 16715 50847
rect 16715 50813 16724 50847
rect 16672 50804 16724 50813
rect 26976 50847 27028 50856
rect 15476 50711 15528 50720
rect 15476 50677 15485 50711
rect 15485 50677 15519 50711
rect 15519 50677 15528 50711
rect 15476 50668 15528 50677
rect 17040 50668 17092 50720
rect 19248 50668 19300 50720
rect 20076 50668 20128 50720
rect 26976 50813 26985 50847
rect 26985 50813 27019 50847
rect 27019 50813 27028 50847
rect 26976 50804 27028 50813
rect 30104 50940 30156 50992
rect 34152 50940 34204 50992
rect 36084 50940 36136 50992
rect 37924 50940 37976 50992
rect 28908 50872 28960 50924
rect 33232 50915 33284 50924
rect 33232 50881 33241 50915
rect 33241 50881 33275 50915
rect 33275 50881 33284 50915
rect 33232 50872 33284 50881
rect 36544 50872 36596 50924
rect 37188 50872 37240 50924
rect 38752 50872 38804 50924
rect 22468 50668 22520 50720
rect 23664 50668 23716 50720
rect 28356 50711 28408 50720
rect 28356 50677 28365 50711
rect 28365 50677 28399 50711
rect 28399 50677 28408 50711
rect 28356 50668 28408 50677
rect 29092 50668 29144 50720
rect 36452 50711 36504 50720
rect 36452 50677 36461 50711
rect 36461 50677 36495 50711
rect 36495 50677 36504 50711
rect 36452 50668 36504 50677
rect 38660 50711 38712 50720
rect 38660 50677 38669 50711
rect 38669 50677 38703 50711
rect 38703 50677 38712 50711
rect 38660 50668 38712 50677
rect 41696 50804 41748 50856
rect 43168 50940 43220 50992
rect 47216 50940 47268 50992
rect 52276 50940 52328 50992
rect 55956 50940 56008 50992
rect 43720 50872 43772 50924
rect 44272 50915 44324 50924
rect 44272 50881 44281 50915
rect 44281 50881 44315 50915
rect 44315 50881 44324 50915
rect 44272 50872 44324 50881
rect 46388 50872 46440 50924
rect 57428 50872 57480 50924
rect 47584 50847 47636 50856
rect 47584 50813 47593 50847
rect 47593 50813 47627 50847
rect 47627 50813 47636 50847
rect 47584 50804 47636 50813
rect 50620 50804 50672 50856
rect 39856 50668 39908 50720
rect 43812 50711 43864 50720
rect 43812 50677 43821 50711
rect 43821 50677 43855 50711
rect 43855 50677 43864 50711
rect 43812 50668 43864 50677
rect 45652 50711 45704 50720
rect 45652 50677 45661 50711
rect 45661 50677 45695 50711
rect 45695 50677 45704 50711
rect 45652 50668 45704 50677
rect 52184 50711 52236 50720
rect 52184 50677 52193 50711
rect 52193 50677 52227 50711
rect 52227 50677 52236 50711
rect 52184 50668 52236 50677
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 3240 50507 3292 50516
rect 3240 50473 3249 50507
rect 3249 50473 3283 50507
rect 3283 50473 3292 50507
rect 3240 50464 3292 50473
rect 5172 50464 5224 50516
rect 6184 50464 6236 50516
rect 11244 50507 11296 50516
rect 11244 50473 11253 50507
rect 11253 50473 11287 50507
rect 11287 50473 11296 50507
rect 11244 50464 11296 50473
rect 14096 50464 14148 50516
rect 15568 50507 15620 50516
rect 15568 50473 15577 50507
rect 15577 50473 15611 50507
rect 15611 50473 15620 50507
rect 15568 50464 15620 50473
rect 17408 50507 17460 50516
rect 17408 50473 17417 50507
rect 17417 50473 17451 50507
rect 17451 50473 17460 50507
rect 17408 50464 17460 50473
rect 23112 50507 23164 50516
rect 23112 50473 23121 50507
rect 23121 50473 23155 50507
rect 23155 50473 23164 50507
rect 23112 50464 23164 50473
rect 25688 50464 25740 50516
rect 30472 50464 30524 50516
rect 37832 50464 37884 50516
rect 47768 50464 47820 50516
rect 57428 50507 57480 50516
rect 57428 50473 57437 50507
rect 57437 50473 57471 50507
rect 57471 50473 57480 50507
rect 57428 50464 57480 50473
rect 1584 50260 1636 50312
rect 5540 50260 5592 50312
rect 2872 50192 2924 50244
rect 19248 50328 19300 50380
rect 21732 50371 21784 50380
rect 21732 50337 21741 50371
rect 21741 50337 21775 50371
rect 21775 50337 21784 50371
rect 21732 50328 21784 50337
rect 36544 50371 36596 50380
rect 36544 50337 36553 50371
rect 36553 50337 36587 50371
rect 36587 50337 36596 50371
rect 36544 50328 36596 50337
rect 39856 50371 39908 50380
rect 39856 50337 39865 50371
rect 39865 50337 39899 50371
rect 39899 50337 39908 50371
rect 39856 50328 39908 50337
rect 55956 50328 56008 50380
rect 7932 50260 7984 50312
rect 8944 50260 8996 50312
rect 13820 50260 13872 50312
rect 15476 50260 15528 50312
rect 17316 50260 17368 50312
rect 6368 50124 6420 50176
rect 7012 50192 7064 50244
rect 8116 50192 8168 50244
rect 10784 50192 10836 50244
rect 16120 50192 16172 50244
rect 21088 50192 21140 50244
rect 13544 50167 13596 50176
rect 13544 50133 13553 50167
rect 13553 50133 13587 50167
rect 13587 50133 13596 50167
rect 13544 50124 13596 50133
rect 24952 50260 25004 50312
rect 26976 50303 27028 50312
rect 26976 50269 26985 50303
rect 26985 50269 27019 50303
rect 27019 50269 27028 50303
rect 26976 50260 27028 50269
rect 28356 50260 28408 50312
rect 29000 50260 29052 50312
rect 29552 50303 29604 50312
rect 29552 50269 29561 50303
rect 29561 50269 29595 50303
rect 29595 50269 29604 50303
rect 29552 50260 29604 50269
rect 30196 50260 30248 50312
rect 24860 50192 24912 50244
rect 30104 50192 30156 50244
rect 34704 50303 34756 50312
rect 34704 50269 34713 50303
rect 34713 50269 34747 50303
rect 34747 50269 34756 50303
rect 34704 50260 34756 50269
rect 36452 50260 36504 50312
rect 36636 50260 36688 50312
rect 40132 50303 40184 50312
rect 40132 50269 40166 50303
rect 40166 50269 40184 50303
rect 40132 50260 40184 50269
rect 41696 50303 41748 50312
rect 41696 50269 41705 50303
rect 41705 50269 41739 50303
rect 41739 50269 41748 50303
rect 41696 50260 41748 50269
rect 41788 50260 41840 50312
rect 44272 50260 44324 50312
rect 47584 50260 47636 50312
rect 50620 50260 50672 50312
rect 52184 50260 52236 50312
rect 31300 50192 31352 50244
rect 46296 50192 46348 50244
rect 28356 50167 28408 50176
rect 28356 50133 28365 50167
rect 28365 50133 28399 50167
rect 28399 50133 28408 50167
rect 28356 50124 28408 50133
rect 32772 50167 32824 50176
rect 32772 50133 32781 50167
rect 32781 50133 32815 50167
rect 32815 50133 32824 50167
rect 32772 50124 32824 50133
rect 36084 50167 36136 50176
rect 36084 50133 36093 50167
rect 36093 50133 36127 50167
rect 36127 50133 36136 50167
rect 36084 50124 36136 50133
rect 41236 50167 41288 50176
rect 41236 50133 41245 50167
rect 41245 50133 41279 50167
rect 41279 50133 41288 50167
rect 41236 50124 41288 50133
rect 41420 50124 41472 50176
rect 56600 50192 56652 50244
rect 52092 50167 52144 50176
rect 52092 50133 52101 50167
rect 52101 50133 52135 50167
rect 52135 50133 52144 50167
rect 52092 50124 52144 50133
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 16120 49963 16172 49972
rect 16120 49929 16129 49963
rect 16129 49929 16163 49963
rect 16163 49929 16172 49963
rect 16120 49920 16172 49929
rect 21088 49963 21140 49972
rect 21088 49929 21097 49963
rect 21097 49929 21131 49963
rect 21131 49929 21140 49963
rect 21088 49920 21140 49929
rect 24492 49963 24544 49972
rect 24492 49929 24501 49963
rect 24501 49929 24535 49963
rect 24535 49929 24544 49963
rect 24492 49920 24544 49929
rect 26240 49920 26292 49972
rect 29920 49920 29972 49972
rect 33232 49920 33284 49972
rect 44272 49920 44324 49972
rect 5816 49852 5868 49904
rect 16028 49852 16080 49904
rect 19248 49852 19300 49904
rect 20076 49852 20128 49904
rect 23480 49852 23532 49904
rect 28356 49852 28408 49904
rect 29092 49895 29144 49904
rect 29092 49861 29126 49895
rect 29126 49861 29144 49895
rect 29092 49852 29144 49861
rect 32496 49895 32548 49904
rect 32496 49861 32505 49895
rect 32505 49861 32539 49895
rect 32539 49861 32548 49895
rect 32496 49852 32548 49861
rect 34796 49852 34848 49904
rect 36084 49852 36136 49904
rect 38660 49852 38712 49904
rect 41236 49852 41288 49904
rect 43076 49852 43128 49904
rect 43812 49852 43864 49904
rect 55404 49920 55456 49972
rect 52092 49852 52144 49904
rect 3516 49784 3568 49836
rect 6460 49784 6512 49836
rect 10232 49784 10284 49836
rect 13728 49784 13780 49836
rect 13912 49784 13964 49836
rect 19340 49784 19392 49836
rect 19708 49827 19760 49836
rect 19708 49793 19717 49827
rect 19717 49793 19751 49827
rect 19751 49793 19760 49827
rect 19708 49784 19760 49793
rect 21088 49784 21140 49836
rect 24860 49784 24912 49836
rect 26424 49784 26476 49836
rect 26976 49827 27028 49836
rect 26976 49793 26985 49827
rect 26985 49793 27019 49827
rect 27019 49793 27028 49827
rect 26976 49784 27028 49793
rect 29552 49784 29604 49836
rect 34704 49827 34756 49836
rect 34704 49793 34713 49827
rect 34713 49793 34747 49827
rect 34747 49793 34756 49827
rect 34704 49784 34756 49793
rect 36544 49784 36596 49836
rect 37280 49827 37332 49836
rect 37280 49793 37289 49827
rect 37289 49793 37323 49827
rect 37323 49793 37332 49827
rect 37280 49784 37332 49793
rect 48780 49827 48832 49836
rect 1584 49759 1636 49768
rect 1584 49725 1593 49759
rect 1593 49725 1627 49759
rect 1627 49725 1636 49759
rect 1584 49716 1636 49725
rect 6368 49759 6420 49768
rect 2964 49623 3016 49632
rect 2964 49589 2973 49623
rect 2973 49589 3007 49623
rect 3007 49589 3016 49623
rect 2964 49580 3016 49589
rect 6368 49725 6377 49759
rect 6377 49725 6411 49759
rect 6411 49725 6420 49759
rect 6368 49716 6420 49725
rect 8944 49716 8996 49768
rect 14740 49759 14792 49768
rect 14740 49725 14749 49759
rect 14749 49725 14783 49759
rect 14783 49725 14792 49759
rect 14740 49716 14792 49725
rect 21732 49716 21784 49768
rect 5448 49648 5500 49700
rect 28724 49716 28776 49768
rect 35992 49716 36044 49768
rect 38752 49716 38804 49768
rect 48780 49793 48789 49827
rect 48789 49793 48823 49827
rect 48823 49793 48832 49827
rect 48780 49784 48832 49793
rect 45008 49716 45060 49768
rect 50620 49759 50672 49768
rect 50620 49725 50629 49759
rect 50629 49725 50663 49759
rect 50663 49725 50672 49759
rect 50620 49716 50672 49725
rect 52736 49716 52788 49768
rect 53932 49784 53984 49836
rect 56784 49784 56836 49836
rect 40408 49648 40460 49700
rect 5816 49623 5868 49632
rect 5816 49589 5825 49623
rect 5825 49589 5859 49623
rect 5859 49589 5868 49623
rect 5816 49580 5868 49589
rect 7748 49623 7800 49632
rect 7748 49589 7757 49623
rect 7757 49589 7791 49623
rect 7791 49589 7800 49623
rect 7748 49580 7800 49589
rect 10416 49623 10468 49632
rect 10416 49589 10425 49623
rect 10425 49589 10459 49623
rect 10459 49589 10468 49623
rect 10416 49580 10468 49589
rect 14372 49580 14424 49632
rect 40500 49623 40552 49632
rect 40500 49589 40509 49623
rect 40509 49589 40543 49623
rect 40543 49589 40552 49623
rect 40500 49580 40552 49589
rect 46756 49623 46808 49632
rect 46756 49589 46765 49623
rect 46765 49589 46799 49623
rect 46799 49589 46808 49623
rect 46756 49580 46808 49589
rect 50160 49623 50212 49632
rect 50160 49589 50169 49623
rect 50169 49589 50203 49623
rect 50203 49589 50212 49623
rect 50160 49580 50212 49589
rect 56324 49623 56376 49632
rect 56324 49589 56333 49623
rect 56333 49589 56367 49623
rect 56367 49589 56376 49623
rect 56324 49580 56376 49589
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 2872 49376 2924 49428
rect 6460 49376 6512 49428
rect 13912 49376 13964 49428
rect 13820 49308 13872 49360
rect 14740 49376 14792 49428
rect 21088 49419 21140 49428
rect 21088 49385 21097 49419
rect 21097 49385 21131 49419
rect 21131 49385 21140 49419
rect 21088 49376 21140 49385
rect 26424 49419 26476 49428
rect 26424 49385 26433 49419
rect 26433 49385 26467 49419
rect 26467 49385 26476 49419
rect 26424 49376 26476 49385
rect 31300 49419 31352 49428
rect 31300 49385 31309 49419
rect 31309 49385 31343 49419
rect 31343 49385 31352 49419
rect 31300 49376 31352 49385
rect 36544 49376 36596 49428
rect 41144 49376 41196 49428
rect 46296 49376 46348 49428
rect 4988 49240 5040 49292
rect 5448 49283 5500 49292
rect 5448 49249 5457 49283
rect 5457 49249 5491 49283
rect 5491 49249 5500 49283
rect 5448 49240 5500 49249
rect 55956 49376 56008 49428
rect 58532 49419 58584 49428
rect 17040 49240 17092 49292
rect 19432 49240 19484 49292
rect 19708 49283 19760 49292
rect 19708 49249 19717 49283
rect 19717 49249 19751 49283
rect 19751 49249 19760 49283
rect 19708 49240 19760 49249
rect 21732 49240 21784 49292
rect 24860 49240 24912 49292
rect 29552 49240 29604 49292
rect 39856 49283 39908 49292
rect 39856 49249 39865 49283
rect 39865 49249 39899 49283
rect 39899 49249 39908 49283
rect 39856 49240 39908 49249
rect 48228 49283 48280 49292
rect 48228 49249 48237 49283
rect 48237 49249 48271 49283
rect 48271 49249 48280 49283
rect 55312 49283 55364 49292
rect 48228 49240 48280 49249
rect 1584 49215 1636 49224
rect 1584 49181 1593 49215
rect 1593 49181 1627 49215
rect 1627 49181 1636 49215
rect 1584 49172 1636 49181
rect 2964 49172 3016 49224
rect 7748 49172 7800 49224
rect 8944 49215 8996 49224
rect 8944 49181 8953 49215
rect 8953 49181 8987 49215
rect 8987 49181 8996 49215
rect 8944 49172 8996 49181
rect 12164 49215 12216 49224
rect 12164 49181 12173 49215
rect 12173 49181 12207 49215
rect 12207 49181 12216 49215
rect 12164 49172 12216 49181
rect 13544 49172 13596 49224
rect 14372 49215 14424 49224
rect 14372 49181 14406 49215
rect 14406 49181 14424 49215
rect 14372 49172 14424 49181
rect 17776 49172 17828 49224
rect 31760 49215 31812 49224
rect 31760 49181 31769 49215
rect 31769 49181 31803 49215
rect 31803 49181 31812 49215
rect 31760 49172 31812 49181
rect 32772 49172 32824 49224
rect 34796 49172 34848 49224
rect 1860 49036 1912 49088
rect 10324 49079 10376 49088
rect 10324 49045 10333 49079
rect 10333 49045 10367 49079
rect 10367 49045 10376 49079
rect 10324 49036 10376 49045
rect 20996 49104 21048 49156
rect 24032 49104 24084 49156
rect 26332 49104 26384 49156
rect 30288 49104 30340 49156
rect 18604 49079 18656 49088
rect 18604 49045 18613 49079
rect 18613 49045 18647 49079
rect 18647 49045 18656 49079
rect 18604 49036 18656 49045
rect 23112 49036 23164 49088
rect 33140 49079 33192 49088
rect 33140 49045 33149 49079
rect 33149 49045 33183 49079
rect 33183 49045 33192 49079
rect 33140 49036 33192 49045
rect 40500 49172 40552 49224
rect 41696 49215 41748 49224
rect 41696 49181 41705 49215
rect 41705 49181 41739 49215
rect 41739 49181 41748 49215
rect 41696 49172 41748 49181
rect 45008 49215 45060 49224
rect 45008 49181 45017 49215
rect 45017 49181 45051 49215
rect 45051 49181 45060 49215
rect 45008 49172 45060 49181
rect 45652 49172 45704 49224
rect 55312 49249 55321 49283
rect 55321 49249 55355 49283
rect 55355 49249 55364 49283
rect 55312 49240 55364 49249
rect 58532 49385 58541 49419
rect 58541 49385 58575 49419
rect 58575 49385 58584 49419
rect 58532 49376 58584 49385
rect 41788 49104 41840 49156
rect 50068 49172 50120 49224
rect 52736 49215 52788 49224
rect 52736 49181 52745 49215
rect 52745 49181 52779 49215
rect 52779 49181 52788 49215
rect 52736 49172 52788 49181
rect 56324 49172 56376 49224
rect 48780 49104 48832 49156
rect 40316 49036 40368 49088
rect 43076 49079 43128 49088
rect 43076 49045 43085 49079
rect 43085 49045 43119 49079
rect 43119 49045 43128 49079
rect 43076 49036 43128 49045
rect 50620 49104 50672 49156
rect 53380 49104 53432 49156
rect 49792 49036 49844 49088
rect 53840 49036 53892 49088
rect 56692 49079 56744 49088
rect 56692 49045 56701 49079
rect 56701 49045 56735 49079
rect 56735 49045 56744 49079
rect 56692 49036 56744 49045
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 3516 48875 3568 48884
rect 3516 48841 3525 48875
rect 3525 48841 3559 48875
rect 3559 48841 3568 48875
rect 3516 48832 3568 48841
rect 10232 48832 10284 48884
rect 20996 48875 21048 48884
rect 20996 48841 21005 48875
rect 21005 48841 21039 48875
rect 21039 48841 21048 48875
rect 20996 48832 21048 48841
rect 26332 48832 26384 48884
rect 41788 48875 41840 48884
rect 41788 48841 41797 48875
rect 41797 48841 41831 48875
rect 41831 48841 41840 48875
rect 41788 48832 41840 48841
rect 46388 48875 46440 48884
rect 46388 48841 46397 48875
rect 46397 48841 46431 48875
rect 46431 48841 46440 48875
rect 46388 48832 46440 48841
rect 56784 48875 56836 48884
rect 56784 48841 56793 48875
rect 56793 48841 56827 48875
rect 56827 48841 56836 48875
rect 56784 48832 56836 48841
rect 5816 48764 5868 48816
rect 10324 48764 10376 48816
rect 4988 48696 5040 48748
rect 5540 48696 5592 48748
rect 8116 48696 8168 48748
rect 12164 48764 12216 48816
rect 12900 48696 12952 48748
rect 18604 48764 18656 48816
rect 33140 48764 33192 48816
rect 13636 48696 13688 48748
rect 15476 48696 15528 48748
rect 17040 48696 17092 48748
rect 19432 48696 19484 48748
rect 20812 48696 20864 48748
rect 22468 48739 22520 48748
rect 22468 48705 22477 48739
rect 22477 48705 22511 48739
rect 22511 48705 22520 48739
rect 22468 48696 22520 48705
rect 24400 48696 24452 48748
rect 24860 48696 24912 48748
rect 26424 48696 26476 48748
rect 32956 48696 33008 48748
rect 34336 48764 34388 48816
rect 41420 48764 41472 48816
rect 43076 48764 43128 48816
rect 50160 48764 50212 48816
rect 55404 48764 55456 48816
rect 35624 48696 35676 48748
rect 37280 48739 37332 48748
rect 37280 48705 37289 48739
rect 37289 48705 37323 48739
rect 37323 48705 37332 48739
rect 37280 48696 37332 48705
rect 38752 48696 38804 48748
rect 41696 48696 41748 48748
rect 42432 48696 42484 48748
rect 1860 48492 1912 48544
rect 30104 48628 30156 48680
rect 11888 48492 11940 48544
rect 14188 48492 14240 48544
rect 14924 48535 14976 48544
rect 14924 48501 14933 48535
rect 14933 48501 14967 48535
rect 14967 48501 14976 48535
rect 14924 48492 14976 48501
rect 18328 48535 18380 48544
rect 18328 48501 18337 48535
rect 18337 48501 18371 48535
rect 18371 48501 18380 48535
rect 18328 48492 18380 48501
rect 23848 48535 23900 48544
rect 23848 48501 23857 48535
rect 23857 48501 23891 48535
rect 23891 48501 23900 48535
rect 23848 48492 23900 48501
rect 31760 48628 31812 48680
rect 40408 48671 40460 48680
rect 40408 48637 40417 48671
rect 40417 48637 40451 48671
rect 40451 48637 40460 48671
rect 40408 48628 40460 48637
rect 44456 48696 44508 48748
rect 48780 48739 48832 48748
rect 48780 48705 48789 48739
rect 48789 48705 48823 48739
rect 48823 48705 48832 48739
rect 48780 48696 48832 48705
rect 53196 48739 53248 48748
rect 53196 48705 53205 48739
rect 53205 48705 53239 48739
rect 53239 48705 53248 48739
rect 53196 48696 53248 48705
rect 56048 48696 56100 48748
rect 45008 48671 45060 48680
rect 45008 48637 45017 48671
rect 45017 48637 45051 48671
rect 45051 48637 45060 48671
rect 45008 48628 45060 48637
rect 55312 48628 55364 48680
rect 50068 48560 50120 48612
rect 31576 48535 31628 48544
rect 31576 48501 31585 48535
rect 31585 48501 31619 48535
rect 31619 48501 31628 48535
rect 31576 48492 31628 48501
rect 33508 48535 33560 48544
rect 33508 48501 33517 48535
rect 33517 48501 33551 48535
rect 33551 48501 33560 48535
rect 33508 48492 33560 48501
rect 34244 48492 34296 48544
rect 38016 48492 38068 48544
rect 42984 48492 43036 48544
rect 52736 48492 52788 48544
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 14832 48288 14884 48340
rect 17040 48288 17092 48340
rect 22468 48288 22520 48340
rect 24860 48288 24912 48340
rect 10784 48263 10836 48272
rect 10784 48229 10793 48263
rect 10793 48229 10827 48263
rect 10827 48229 10836 48263
rect 10784 48220 10836 48229
rect 12900 48263 12952 48272
rect 12900 48229 12909 48263
rect 12909 48229 12943 48263
rect 12943 48229 12952 48263
rect 12900 48220 12952 48229
rect 16028 48263 16080 48272
rect 16028 48229 16037 48263
rect 16037 48229 16071 48263
rect 16071 48229 16080 48263
rect 16028 48220 16080 48229
rect 4988 48195 5040 48204
rect 4988 48161 4997 48195
rect 4997 48161 5031 48195
rect 5031 48161 5040 48195
rect 4988 48152 5040 48161
rect 20812 48263 20864 48272
rect 20812 48229 20821 48263
rect 20821 48229 20855 48263
rect 20855 48229 20864 48263
rect 20812 48220 20864 48229
rect 32956 48288 33008 48340
rect 48228 48288 48280 48340
rect 53380 48331 53432 48340
rect 43720 48220 43772 48272
rect 53380 48297 53389 48331
rect 53389 48297 53423 48331
rect 53423 48297 53432 48331
rect 53380 48288 53432 48297
rect 50068 48220 50120 48272
rect 19432 48195 19484 48204
rect 19432 48161 19441 48195
rect 19441 48161 19475 48195
rect 19475 48161 19484 48195
rect 19432 48152 19484 48161
rect 36544 48195 36596 48204
rect 8944 48084 8996 48136
rect 5908 48016 5960 48068
rect 10416 48084 10468 48136
rect 11520 48127 11572 48136
rect 11520 48093 11529 48127
rect 11529 48093 11563 48127
rect 11563 48093 11572 48127
rect 11520 48084 11572 48093
rect 14924 48127 14976 48136
rect 14924 48093 14958 48127
rect 14958 48093 14976 48127
rect 12900 48016 12952 48068
rect 14924 48084 14976 48093
rect 18328 48084 18380 48136
rect 21180 48084 21232 48136
rect 25780 48084 25832 48136
rect 30104 48084 30156 48136
rect 31576 48084 31628 48136
rect 32220 48127 32272 48136
rect 32220 48093 32229 48127
rect 32229 48093 32263 48127
rect 32263 48093 32272 48127
rect 32220 48084 32272 48093
rect 33508 48084 33560 48136
rect 34336 48084 34388 48136
rect 36544 48161 36553 48195
rect 36553 48161 36587 48195
rect 36587 48161 36596 48195
rect 36544 48152 36596 48161
rect 42432 48195 42484 48204
rect 42432 48161 42441 48195
rect 42441 48161 42475 48195
rect 42475 48161 42484 48195
rect 42432 48152 42484 48161
rect 45008 48152 45060 48204
rect 48228 48195 48280 48204
rect 48228 48161 48237 48195
rect 48237 48161 48271 48195
rect 48271 48161 48280 48195
rect 48228 48152 48280 48161
rect 56600 48220 56652 48272
rect 40408 48084 40460 48136
rect 42984 48084 43036 48136
rect 49792 48084 49844 48136
rect 52736 48084 52788 48136
rect 55312 48127 55364 48136
rect 55312 48093 55321 48127
rect 55321 48093 55355 48127
rect 55355 48093 55364 48127
rect 55312 48084 55364 48093
rect 56692 48084 56744 48136
rect 14832 48016 14884 48068
rect 20904 48016 20956 48068
rect 35992 48016 36044 48068
rect 6368 47991 6420 48000
rect 6368 47957 6377 47991
rect 6377 47957 6411 47991
rect 6411 47957 6420 47991
rect 6368 47948 6420 47957
rect 18420 47991 18472 48000
rect 18420 47957 18429 47991
rect 18429 47957 18463 47991
rect 18463 47957 18472 47991
rect 18420 47948 18472 47957
rect 31760 47991 31812 48000
rect 31760 47957 31769 47991
rect 31769 47957 31803 47991
rect 31803 47957 31812 47991
rect 31760 47948 31812 47957
rect 41144 48016 41196 48068
rect 46388 48016 46440 48068
rect 49700 48016 49752 48068
rect 54116 48016 54168 48068
rect 37924 47991 37976 48000
rect 37924 47957 37933 47991
rect 37933 47957 37967 47991
rect 37967 47957 37976 47991
rect 37924 47948 37976 47957
rect 41788 47948 41840 48000
rect 47860 47948 47912 48000
rect 49608 47991 49660 48000
rect 49608 47957 49617 47991
rect 49617 47957 49651 47991
rect 49651 47957 49660 47991
rect 49608 47948 49660 47957
rect 50896 47948 50948 48000
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 15476 47787 15528 47796
rect 15476 47753 15485 47787
rect 15485 47753 15519 47787
rect 15519 47753 15528 47787
rect 15476 47744 15528 47753
rect 20904 47787 20956 47796
rect 20904 47753 20913 47787
rect 20913 47753 20947 47787
rect 20947 47753 20956 47787
rect 20904 47744 20956 47753
rect 24400 47787 24452 47796
rect 24400 47753 24409 47787
rect 24409 47753 24443 47787
rect 24443 47753 24452 47787
rect 24400 47744 24452 47753
rect 26424 47787 26476 47796
rect 26424 47753 26433 47787
rect 26433 47753 26467 47787
rect 26467 47753 26476 47787
rect 26424 47744 26476 47753
rect 35624 47787 35676 47796
rect 35624 47753 35633 47787
rect 35633 47753 35667 47787
rect 35667 47753 35676 47787
rect 35624 47744 35676 47753
rect 44456 47787 44508 47796
rect 44456 47753 44465 47787
rect 44465 47753 44499 47787
rect 44499 47753 44508 47787
rect 44456 47744 44508 47753
rect 50068 47787 50120 47796
rect 50068 47753 50077 47787
rect 50077 47753 50111 47787
rect 50111 47753 50120 47787
rect 50068 47744 50120 47753
rect 54116 47787 54168 47796
rect 54116 47753 54125 47787
rect 54125 47753 54159 47787
rect 54159 47753 54168 47787
rect 54116 47744 54168 47753
rect 4988 47676 5040 47728
rect 11888 47719 11940 47728
rect 11888 47685 11897 47719
rect 11897 47685 11931 47719
rect 11931 47685 11940 47719
rect 11888 47676 11940 47685
rect 18420 47676 18472 47728
rect 26240 47676 26292 47728
rect 29000 47676 29052 47728
rect 31760 47676 31812 47728
rect 40316 47676 40368 47728
rect 46756 47676 46808 47728
rect 53196 47676 53248 47728
rect 5172 47608 5224 47660
rect 7748 47608 7800 47660
rect 14188 47608 14240 47660
rect 17040 47608 17092 47660
rect 19432 47608 19484 47660
rect 20904 47608 20956 47660
rect 22468 47608 22520 47660
rect 24860 47608 24912 47660
rect 26792 47608 26844 47660
rect 32220 47608 32272 47660
rect 34336 47608 34388 47660
rect 34520 47651 34572 47660
rect 34520 47617 34554 47651
rect 34554 47617 34572 47651
rect 34520 47608 34572 47617
rect 36544 47608 36596 47660
rect 37372 47608 37424 47660
rect 42432 47608 42484 47660
rect 45652 47608 45704 47660
rect 52552 47608 52604 47660
rect 4988 47540 5040 47592
rect 5448 47540 5500 47592
rect 13636 47583 13688 47592
rect 13636 47549 13645 47583
rect 13645 47549 13679 47583
rect 13679 47549 13688 47583
rect 13636 47540 13688 47549
rect 5724 47404 5776 47456
rect 7288 47404 7340 47456
rect 27620 47540 27672 47592
rect 41328 47583 41380 47592
rect 41328 47549 41337 47583
rect 41337 47549 41371 47583
rect 41371 47549 41380 47583
rect 41328 47540 41380 47549
rect 52736 47583 52788 47592
rect 52736 47549 52745 47583
rect 52745 47549 52779 47583
rect 52779 47549 52788 47583
rect 52736 47540 52788 47549
rect 14832 47404 14884 47456
rect 18328 47447 18380 47456
rect 18328 47413 18337 47447
rect 18337 47413 18371 47447
rect 18371 47413 18380 47447
rect 18328 47404 18380 47413
rect 30012 47447 30064 47456
rect 30012 47413 30021 47447
rect 30021 47413 30055 47447
rect 30055 47413 30064 47447
rect 30012 47404 30064 47413
rect 33784 47447 33836 47456
rect 33784 47413 33793 47447
rect 33793 47413 33827 47447
rect 33827 47413 33836 47447
rect 33784 47404 33836 47413
rect 38660 47447 38712 47456
rect 38660 47413 38669 47447
rect 38669 47413 38703 47447
rect 38703 47413 38712 47447
rect 38660 47404 38712 47413
rect 44548 47404 44600 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 5172 47243 5224 47252
rect 5172 47209 5181 47243
rect 5181 47209 5215 47243
rect 5215 47209 5224 47243
rect 5172 47200 5224 47209
rect 5816 47200 5868 47252
rect 20904 47243 20956 47252
rect 20904 47209 20913 47243
rect 20913 47209 20947 47243
rect 20947 47209 20956 47243
rect 20904 47200 20956 47209
rect 26792 47243 26844 47252
rect 26792 47209 26801 47243
rect 26801 47209 26835 47243
rect 26835 47209 26844 47243
rect 26792 47200 26844 47209
rect 35992 47200 36044 47252
rect 46388 47243 46440 47252
rect 46388 47209 46397 47243
rect 46397 47209 46431 47243
rect 46431 47209 46440 47243
rect 46388 47200 46440 47209
rect 49700 47200 49752 47252
rect 53932 47243 53984 47252
rect 53932 47209 53941 47243
rect 53941 47209 53975 47243
rect 53975 47209 53984 47243
rect 53932 47200 53984 47209
rect 29184 47132 29236 47184
rect 5448 47064 5500 47116
rect 19432 47064 19484 47116
rect 22468 47107 22520 47116
rect 22468 47073 22477 47107
rect 22477 47073 22511 47107
rect 22511 47073 22520 47107
rect 22468 47064 22520 47073
rect 24860 47064 24912 47116
rect 27620 47107 27672 47116
rect 4344 46996 4396 47048
rect 5724 46996 5776 47048
rect 11428 46996 11480 47048
rect 14832 47039 14884 47048
rect 14832 47005 14841 47039
rect 14841 47005 14875 47039
rect 14875 47005 14884 47039
rect 14832 46996 14884 47005
rect 16948 46996 17000 47048
rect 18328 46996 18380 47048
rect 23848 46996 23900 47048
rect 27620 47073 27629 47107
rect 27629 47073 27663 47107
rect 27663 47073 27672 47107
rect 27620 47064 27672 47073
rect 48228 47107 48280 47116
rect 48228 47073 48237 47107
rect 48237 47073 48271 47107
rect 48271 47073 48280 47107
rect 48228 47064 48280 47073
rect 30012 46996 30064 47048
rect 30104 46996 30156 47048
rect 33784 46996 33836 47048
rect 34428 46996 34480 47048
rect 5540 46928 5592 46980
rect 12164 46928 12216 46980
rect 17960 46928 18012 46980
rect 20996 46928 21048 46980
rect 26424 46928 26476 46980
rect 35348 46928 35400 46980
rect 37924 46996 37976 47048
rect 40408 46996 40460 47048
rect 41328 46996 41380 47048
rect 41788 46996 41840 47048
rect 46940 46996 46992 47048
rect 49608 46996 49660 47048
rect 50620 47039 50672 47048
rect 50620 47005 50629 47039
rect 50629 47005 50663 47039
rect 50663 47005 50672 47039
rect 50620 46996 50672 47005
rect 50896 47039 50948 47048
rect 50896 47005 50930 47039
rect 50930 47005 50948 47039
rect 50896 46996 50948 47005
rect 37464 46928 37516 46980
rect 40132 46971 40184 46980
rect 40132 46937 40166 46971
rect 40166 46937 40184 46971
rect 40132 46928 40184 46937
rect 46204 46928 46256 46980
rect 52460 46928 52512 46980
rect 53840 46996 53892 47048
rect 52736 46928 52788 46980
rect 53656 46928 53708 46980
rect 55312 46928 55364 46980
rect 11980 46903 12032 46912
rect 11980 46869 11989 46903
rect 11989 46869 12023 46903
rect 12023 46869 12032 46903
rect 11980 46860 12032 46869
rect 16212 46903 16264 46912
rect 16212 46869 16221 46903
rect 16221 46869 16255 46903
rect 16255 46869 16264 46903
rect 16212 46860 16264 46869
rect 18236 46903 18288 46912
rect 18236 46869 18245 46903
rect 18245 46869 18279 46903
rect 18279 46869 18288 46903
rect 18236 46860 18288 46869
rect 23848 46903 23900 46912
rect 23848 46869 23857 46903
rect 23857 46869 23891 46903
rect 23891 46869 23900 46903
rect 23848 46860 23900 46869
rect 32496 46903 32548 46912
rect 32496 46869 32505 46903
rect 32505 46869 32539 46903
rect 32539 46869 32548 46903
rect 32496 46860 32548 46869
rect 37280 46860 37332 46912
rect 41236 46903 41288 46912
rect 41236 46869 41245 46903
rect 41245 46869 41279 46903
rect 41279 46869 41288 46903
rect 41236 46860 41288 46869
rect 43076 46903 43128 46912
rect 43076 46869 43085 46903
rect 43085 46869 43119 46903
rect 43119 46869 43128 46903
rect 43076 46860 43128 46869
rect 52000 46903 52052 46912
rect 52000 46869 52009 46903
rect 52009 46869 52043 46903
rect 52043 46869 52052 46903
rect 52000 46860 52052 46869
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 5540 46656 5592 46708
rect 7748 46699 7800 46708
rect 7748 46665 7757 46699
rect 7757 46665 7791 46699
rect 7791 46665 7800 46699
rect 7748 46656 7800 46665
rect 12900 46699 12952 46708
rect 12900 46665 12909 46699
rect 12909 46665 12943 46699
rect 12943 46665 12952 46699
rect 12900 46656 12952 46665
rect 20996 46699 21048 46708
rect 20996 46665 21005 46699
rect 21005 46665 21039 46699
rect 21039 46665 21048 46699
rect 20996 46656 21048 46665
rect 24032 46699 24084 46708
rect 24032 46665 24041 46699
rect 24041 46665 24075 46699
rect 24075 46665 24084 46699
rect 24032 46656 24084 46665
rect 26424 46699 26476 46708
rect 26424 46665 26433 46699
rect 26433 46665 26467 46699
rect 26467 46665 26476 46699
rect 26424 46656 26476 46665
rect 35348 46699 35400 46708
rect 35348 46665 35357 46699
rect 35357 46665 35391 46699
rect 35391 46665 35400 46699
rect 35348 46656 35400 46665
rect 45652 46699 45704 46708
rect 45652 46665 45661 46699
rect 45661 46665 45695 46699
rect 45695 46665 45704 46699
rect 45652 46656 45704 46665
rect 4620 46588 4672 46640
rect 6368 46588 6420 46640
rect 11980 46588 12032 46640
rect 16212 46588 16264 46640
rect 18236 46588 18288 46640
rect 23848 46588 23900 46640
rect 32496 46588 32548 46640
rect 34244 46631 34296 46640
rect 34244 46597 34278 46631
rect 34278 46597 34296 46631
rect 34244 46588 34296 46597
rect 34428 46588 34480 46640
rect 38660 46588 38712 46640
rect 41236 46588 41288 46640
rect 47860 46631 47912 46640
rect 47860 46597 47894 46631
rect 47894 46597 47912 46631
rect 47860 46588 47912 46597
rect 3240 46520 3292 46572
rect 4344 46520 4396 46572
rect 7840 46520 7892 46572
rect 13636 46520 13688 46572
rect 19432 46520 19484 46572
rect 21088 46520 21140 46572
rect 22560 46520 22612 46572
rect 24860 46520 24912 46572
rect 26240 46520 26292 46572
rect 29092 46563 29144 46572
rect 29092 46529 29126 46563
rect 29126 46529 29144 46563
rect 29092 46520 29144 46529
rect 1860 46452 1912 46504
rect 5448 46452 5500 46504
rect 11520 46495 11572 46504
rect 11520 46461 11529 46495
rect 11529 46461 11563 46495
rect 11563 46461 11572 46495
rect 11520 46452 11572 46461
rect 8944 46316 8996 46368
rect 9588 46359 9640 46368
rect 9588 46325 9597 46359
rect 9597 46325 9631 46359
rect 9631 46325 9640 46359
rect 9588 46316 9640 46325
rect 16120 46359 16172 46368
rect 16120 46325 16129 46359
rect 16129 46325 16163 46359
rect 16163 46325 16172 46359
rect 16120 46316 16172 46325
rect 18144 46359 18196 46368
rect 18144 46325 18153 46359
rect 18153 46325 18187 46359
rect 18187 46325 18196 46359
rect 18144 46316 18196 46325
rect 30012 46316 30064 46368
rect 30196 46359 30248 46368
rect 30196 46325 30205 46359
rect 30205 46325 30239 46359
rect 30239 46325 30248 46359
rect 30196 46316 30248 46325
rect 33508 46359 33560 46368
rect 33508 46325 33517 46359
rect 33517 46325 33551 46359
rect 33551 46325 33560 46359
rect 33508 46316 33560 46325
rect 40408 46520 40460 46572
rect 42432 46563 42484 46572
rect 42432 46529 42441 46563
rect 42441 46529 42475 46563
rect 42475 46529 42484 46563
rect 42432 46520 42484 46529
rect 43812 46520 43864 46572
rect 44180 46520 44232 46572
rect 46940 46520 46992 46572
rect 48228 46520 48280 46572
rect 50620 46656 50672 46708
rect 52000 46588 52052 46640
rect 53656 46563 53708 46572
rect 53656 46529 53665 46563
rect 53665 46529 53699 46563
rect 53699 46529 53708 46563
rect 53656 46520 53708 46529
rect 55496 46520 55548 46572
rect 56692 46520 56744 46572
rect 44272 46495 44324 46504
rect 44272 46461 44281 46495
rect 44281 46461 44315 46495
rect 44315 46461 44324 46495
rect 44272 46452 44324 46461
rect 55312 46452 55364 46504
rect 38752 46384 38804 46436
rect 37464 46316 37516 46368
rect 40684 46316 40736 46368
rect 42800 46316 42852 46368
rect 48964 46359 49016 46368
rect 48964 46325 48973 46359
rect 48973 46325 49007 46359
rect 49007 46325 49016 46359
rect 48964 46316 49016 46325
rect 51540 46359 51592 46368
rect 51540 46325 51549 46359
rect 51549 46325 51583 46359
rect 51583 46325 51592 46359
rect 51540 46316 51592 46325
rect 55036 46359 55088 46368
rect 55036 46325 55045 46359
rect 55045 46325 55079 46359
rect 55079 46325 55088 46359
rect 55036 46316 55088 46325
rect 57244 46316 57296 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 3240 46155 3292 46164
rect 3240 46121 3249 46155
rect 3249 46121 3283 46155
rect 3283 46121 3292 46155
rect 3240 46112 3292 46121
rect 5448 46112 5500 46164
rect 5908 46155 5960 46164
rect 5908 46121 5917 46155
rect 5917 46121 5951 46155
rect 5951 46121 5960 46155
rect 5908 46112 5960 46121
rect 7840 46155 7892 46164
rect 7840 46121 7849 46155
rect 7849 46121 7883 46155
rect 7883 46121 7892 46155
rect 7840 46112 7892 46121
rect 12164 46155 12216 46164
rect 12164 46121 12173 46155
rect 12173 46121 12207 46155
rect 12207 46121 12216 46155
rect 12164 46112 12216 46121
rect 1860 46019 1912 46028
rect 1860 45985 1869 46019
rect 1869 45985 1903 46019
rect 1903 45985 1912 46019
rect 1860 45976 1912 45985
rect 4528 46019 4580 46028
rect 4528 45985 4537 46019
rect 4537 45985 4571 46019
rect 4571 45985 4580 46019
rect 4528 45976 4580 45985
rect 16948 46112 17000 46164
rect 21088 46155 21140 46164
rect 21088 46121 21097 46155
rect 21097 46121 21131 46155
rect 21131 46121 21140 46155
rect 21088 46112 21140 46121
rect 23756 46112 23808 46164
rect 26240 46155 26292 46164
rect 26240 46121 26249 46155
rect 26249 46121 26283 46155
rect 26283 46121 26292 46155
rect 29000 46155 29052 46164
rect 26240 46112 26292 46121
rect 29000 46121 29009 46155
rect 29009 46121 29043 46155
rect 29043 46121 29052 46155
rect 29000 46112 29052 46121
rect 34520 46112 34572 46164
rect 37372 46112 37424 46164
rect 40132 46112 40184 46164
rect 43812 46155 43864 46164
rect 43812 46121 43821 46155
rect 43821 46121 43855 46155
rect 43855 46121 43864 46155
rect 43812 46112 43864 46121
rect 46204 46112 46256 46164
rect 52552 46112 52604 46164
rect 56692 46155 56744 46164
rect 56692 46121 56701 46155
rect 56701 46121 56735 46155
rect 56735 46121 56744 46155
rect 56692 46112 56744 46121
rect 5816 45908 5868 45960
rect 7288 45908 7340 45960
rect 8944 45951 8996 45960
rect 8944 45917 8953 45951
rect 8953 45917 8987 45951
rect 8987 45917 8996 45951
rect 8944 45908 8996 45917
rect 11520 45908 11572 45960
rect 4620 45840 4672 45892
rect 8576 45840 8628 45892
rect 12900 45840 12952 45892
rect 16120 45908 16172 45960
rect 14832 45840 14884 45892
rect 19432 45976 19484 46028
rect 24860 46019 24912 46028
rect 24860 45985 24869 46019
rect 24869 45985 24903 46019
rect 24903 45985 24912 46019
rect 24860 45976 24912 45985
rect 27620 46019 27672 46028
rect 27620 45985 27629 46019
rect 27629 45985 27663 46019
rect 27663 45985 27672 46019
rect 27620 45976 27672 45985
rect 30012 45976 30064 46028
rect 18144 45908 18196 45960
rect 22560 45908 22612 45960
rect 23112 45908 23164 45960
rect 30196 45908 30248 45960
rect 34428 45976 34480 46028
rect 37464 46019 37516 46028
rect 37464 45985 37473 46019
rect 37473 45985 37507 46019
rect 37507 45985 37516 46019
rect 37464 45976 37516 45985
rect 44272 45976 44324 46028
rect 33508 45908 33560 45960
rect 37280 45908 37332 45960
rect 38016 45908 38068 45960
rect 40592 45951 40644 45960
rect 21272 45840 21324 45892
rect 24952 45840 25004 45892
rect 31208 45840 31260 45892
rect 40592 45917 40601 45951
rect 40601 45917 40635 45951
rect 40635 45917 40644 45951
rect 40592 45908 40644 45917
rect 40684 45908 40736 45960
rect 41328 45908 41380 45960
rect 42432 45951 42484 45960
rect 42432 45917 42441 45951
rect 42441 45917 42475 45951
rect 42475 45917 42484 45951
rect 42432 45908 42484 45917
rect 43076 45908 43128 45960
rect 50068 45976 50120 46028
rect 55312 46019 55364 46028
rect 55312 45985 55321 46019
rect 55321 45985 55355 46019
rect 55355 45985 55364 46019
rect 55312 45976 55364 45985
rect 45744 45908 45796 45960
rect 46940 45908 46992 45960
rect 48964 45908 49016 45960
rect 51540 45908 51592 45960
rect 52460 45908 52512 45960
rect 45652 45840 45704 45892
rect 53380 45840 53432 45892
rect 56692 45840 56744 45892
rect 10324 45815 10376 45824
rect 10324 45781 10333 45815
rect 10333 45781 10367 45815
rect 10367 45781 10376 45815
rect 10324 45772 10376 45781
rect 15752 45815 15804 45824
rect 15752 45781 15761 45815
rect 15761 45781 15795 45815
rect 15795 45781 15804 45815
rect 15752 45772 15804 45781
rect 18052 45815 18104 45824
rect 18052 45781 18061 45815
rect 18061 45781 18095 45815
rect 18095 45781 18104 45815
rect 18052 45772 18104 45781
rect 30288 45772 30340 45824
rect 41972 45815 42024 45824
rect 41972 45781 41981 45815
rect 41981 45781 42015 45815
rect 42015 45781 42024 45815
rect 41972 45772 42024 45781
rect 48228 45815 48280 45824
rect 48228 45781 48237 45815
rect 48237 45781 48271 45815
rect 48271 45781 48280 45815
rect 48228 45772 48280 45781
rect 53748 45815 53800 45824
rect 53748 45781 53757 45815
rect 53757 45781 53791 45815
rect 53791 45781 53800 45815
rect 53748 45772 53800 45781
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 4620 45568 4672 45620
rect 8576 45611 8628 45620
rect 8576 45577 8585 45611
rect 8585 45577 8619 45611
rect 8619 45577 8628 45611
rect 8576 45568 8628 45577
rect 12900 45611 12952 45620
rect 12900 45577 12909 45611
rect 12909 45577 12943 45611
rect 12943 45577 12952 45611
rect 12900 45568 12952 45577
rect 21272 45611 21324 45620
rect 21272 45577 21281 45611
rect 21281 45577 21315 45611
rect 21315 45577 21324 45611
rect 21272 45568 21324 45577
rect 45652 45611 45704 45620
rect 45652 45577 45661 45611
rect 45661 45577 45695 45611
rect 45695 45577 45704 45611
rect 45652 45568 45704 45577
rect 55496 45568 55548 45620
rect 10324 45500 10376 45552
rect 13636 45500 13688 45552
rect 3148 45432 3200 45484
rect 1676 45364 1728 45416
rect 9588 45432 9640 45484
rect 11520 45475 11572 45484
rect 11520 45441 11529 45475
rect 11529 45441 11563 45475
rect 11563 45441 11572 45475
rect 11520 45432 11572 45441
rect 12900 45432 12952 45484
rect 15752 45500 15804 45552
rect 18052 45500 18104 45552
rect 19984 45432 20036 45484
rect 21364 45432 21416 45484
rect 23204 45432 23256 45484
rect 25044 45500 25096 45552
rect 25780 45432 25832 45484
rect 30104 45432 30156 45484
rect 31484 45432 31536 45484
rect 7196 45407 7248 45416
rect 7196 45373 7205 45407
rect 7205 45373 7239 45407
rect 7239 45373 7248 45407
rect 7196 45364 7248 45373
rect 9036 45407 9088 45416
rect 9036 45373 9045 45407
rect 9045 45373 9079 45407
rect 9079 45373 9088 45407
rect 9036 45364 9088 45373
rect 16672 45407 16724 45416
rect 16672 45373 16681 45407
rect 16681 45373 16715 45407
rect 16715 45373 16724 45407
rect 16672 45364 16724 45373
rect 21824 45407 21876 45416
rect 21824 45373 21833 45407
rect 21833 45373 21867 45407
rect 21867 45373 21876 45407
rect 21824 45364 21876 45373
rect 27712 45364 27764 45416
rect 17960 45296 18012 45348
rect 6368 45228 6420 45280
rect 7196 45228 7248 45280
rect 10416 45271 10468 45280
rect 10416 45237 10425 45271
rect 10425 45237 10459 45271
rect 10459 45237 10468 45271
rect 10416 45228 10468 45237
rect 15476 45271 15528 45280
rect 15476 45237 15485 45271
rect 15485 45237 15519 45271
rect 15519 45237 15528 45271
rect 15476 45228 15528 45237
rect 20260 45228 20312 45280
rect 25688 45271 25740 45280
rect 25688 45237 25697 45271
rect 25697 45237 25731 45271
rect 25731 45237 25740 45271
rect 25688 45228 25740 45237
rect 29736 45271 29788 45280
rect 29736 45237 29745 45271
rect 29745 45237 29779 45271
rect 29779 45237 29788 45271
rect 29736 45228 29788 45237
rect 31668 45364 31720 45416
rect 34796 45432 34848 45484
rect 36544 45432 36596 45484
rect 39212 45432 39264 45484
rect 40592 45500 40644 45552
rect 42800 45500 42852 45552
rect 44548 45543 44600 45552
rect 44548 45509 44582 45543
rect 44582 45509 44600 45543
rect 44548 45500 44600 45509
rect 48228 45500 48280 45552
rect 41972 45432 42024 45484
rect 42432 45475 42484 45484
rect 42432 45441 42441 45475
rect 42441 45441 42475 45475
rect 42475 45441 42484 45475
rect 42432 45432 42484 45441
rect 42524 45432 42576 45484
rect 46940 45432 46992 45484
rect 47584 45475 47636 45484
rect 47584 45441 47593 45475
rect 47593 45441 47627 45475
rect 47627 45441 47636 45475
rect 47584 45432 47636 45441
rect 51540 45432 51592 45484
rect 54024 45432 54076 45484
rect 37924 45364 37976 45416
rect 49424 45364 49476 45416
rect 52736 45407 52788 45416
rect 52736 45373 52745 45407
rect 52745 45373 52779 45407
rect 52779 45373 52788 45407
rect 52736 45364 52788 45373
rect 41144 45296 41196 45348
rect 44180 45296 44232 45348
rect 30380 45228 30432 45280
rect 31576 45271 31628 45280
rect 31576 45237 31585 45271
rect 31585 45237 31619 45271
rect 31619 45237 31628 45271
rect 31576 45228 31628 45237
rect 33784 45228 33836 45280
rect 35348 45228 35400 45280
rect 39396 45271 39448 45280
rect 39396 45237 39405 45271
rect 39405 45237 39439 45271
rect 39439 45237 39448 45271
rect 39396 45228 39448 45237
rect 48964 45271 49016 45280
rect 48964 45237 48973 45271
rect 48973 45237 49007 45271
rect 49007 45237 49016 45271
rect 48964 45228 49016 45237
rect 52092 45228 52144 45280
rect 56508 45228 56560 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 3148 45067 3200 45076
rect 3148 45033 3157 45067
rect 3157 45033 3191 45067
rect 3191 45033 3200 45067
rect 3148 45024 3200 45033
rect 21364 45067 21416 45076
rect 21364 45033 21373 45067
rect 21373 45033 21407 45067
rect 21407 45033 21416 45067
rect 21364 45024 21416 45033
rect 23204 45067 23256 45076
rect 23204 45033 23213 45067
rect 23213 45033 23247 45067
rect 23247 45033 23256 45067
rect 23204 45024 23256 45033
rect 29092 45024 29144 45076
rect 31208 45024 31260 45076
rect 51540 45067 51592 45076
rect 51540 45033 51549 45067
rect 51549 45033 51583 45067
rect 51583 45033 51592 45067
rect 51540 45024 51592 45033
rect 53380 45067 53432 45076
rect 53380 45033 53389 45067
rect 53389 45033 53423 45067
rect 53423 45033 53432 45067
rect 53380 45024 53432 45033
rect 56692 45067 56744 45076
rect 56692 45033 56701 45067
rect 56701 45033 56735 45067
rect 56735 45033 56744 45067
rect 56692 45024 56744 45033
rect 16672 44888 16724 44940
rect 19984 44931 20036 44940
rect 19984 44897 19993 44931
rect 19993 44897 20027 44931
rect 20027 44897 20036 44931
rect 19984 44888 20036 44897
rect 45744 44931 45796 44940
rect 45744 44897 45753 44931
rect 45753 44897 45787 44931
rect 45787 44897 45796 44931
rect 45744 44888 45796 44897
rect 47584 44931 47636 44940
rect 47584 44897 47593 44931
rect 47593 44897 47627 44931
rect 47627 44897 47636 44931
rect 47584 44888 47636 44897
rect 56508 44888 56560 44940
rect 1676 44820 1728 44872
rect 6368 44863 6420 44872
rect 6368 44829 6377 44863
rect 6377 44829 6411 44863
rect 6411 44829 6420 44863
rect 6368 44820 6420 44829
rect 9036 44820 9088 44872
rect 9496 44820 9548 44872
rect 10784 44863 10836 44872
rect 10784 44829 10793 44863
rect 10793 44829 10827 44863
rect 10827 44829 10836 44863
rect 10784 44820 10836 44829
rect 14096 44863 14148 44872
rect 14096 44829 14105 44863
rect 14105 44829 14139 44863
rect 14139 44829 14148 44863
rect 14096 44820 14148 44829
rect 15476 44820 15528 44872
rect 20260 44863 20312 44872
rect 20260 44829 20294 44863
rect 20294 44829 20312 44863
rect 20260 44820 20312 44829
rect 21548 44820 21600 44872
rect 3056 44752 3108 44804
rect 7656 44752 7708 44804
rect 9588 44752 9640 44804
rect 7748 44727 7800 44736
rect 7748 44693 7757 44727
rect 7757 44693 7791 44727
rect 7791 44693 7800 44727
rect 7748 44684 7800 44693
rect 23020 44820 23072 44872
rect 27712 44820 27764 44872
rect 29736 44820 29788 44872
rect 30380 44820 30432 44872
rect 31668 44820 31720 44872
rect 37924 44863 37976 44872
rect 37924 44829 37933 44863
rect 37933 44829 37967 44863
rect 37967 44829 37976 44863
rect 37924 44820 37976 44829
rect 40408 44820 40460 44872
rect 42432 44863 42484 44872
rect 42432 44829 42441 44863
rect 42441 44829 42475 44863
rect 42475 44829 42484 44863
rect 42432 44820 42484 44829
rect 48964 44820 49016 44872
rect 52736 44820 52788 44872
rect 54576 44820 54628 44872
rect 57244 44820 57296 44872
rect 23112 44752 23164 44804
rect 27528 44752 27580 44804
rect 32036 44752 32088 44804
rect 34060 44752 34112 44804
rect 38016 44752 38068 44804
rect 39120 44752 39172 44804
rect 41880 44752 41932 44804
rect 42708 44795 42760 44804
rect 42708 44761 42742 44795
rect 42742 44761 42760 44795
rect 42708 44752 42760 44761
rect 48872 44752 48924 44804
rect 51356 44752 51408 44804
rect 53380 44752 53432 44804
rect 55956 44752 56008 44804
rect 12164 44727 12216 44736
rect 12164 44693 12173 44727
rect 12173 44693 12207 44727
rect 12207 44693 12216 44727
rect 12164 44684 12216 44693
rect 15476 44727 15528 44736
rect 15476 44693 15485 44727
rect 15485 44693 15519 44727
rect 15519 44693 15528 44727
rect 15476 44684 15528 44693
rect 18236 44727 18288 44736
rect 18236 44693 18245 44727
rect 18245 44693 18279 44727
rect 18279 44693 18288 44727
rect 18236 44684 18288 44693
rect 27160 44727 27212 44736
rect 27160 44693 27169 44727
rect 27169 44693 27203 44727
rect 27203 44693 27212 44727
rect 27160 44684 27212 44693
rect 31944 44684 31996 44736
rect 36728 44684 36780 44736
rect 39304 44727 39356 44736
rect 39304 44693 39313 44727
rect 39313 44693 39347 44727
rect 39347 44693 39356 44727
rect 39304 44684 39356 44693
rect 41052 44684 41104 44736
rect 43812 44727 43864 44736
rect 43812 44693 43821 44727
rect 43821 44693 43855 44727
rect 43855 44693 43864 44727
rect 43812 44684 43864 44693
rect 47124 44727 47176 44736
rect 47124 44693 47133 44727
rect 47133 44693 47167 44727
rect 47167 44693 47176 44727
rect 47124 44684 47176 44693
rect 48964 44727 49016 44736
rect 48964 44693 48973 44727
rect 48973 44693 49007 44727
rect 49007 44693 49016 44727
rect 48964 44684 49016 44693
rect 58532 44727 58584 44736
rect 58532 44693 58541 44727
rect 58541 44693 58575 44727
rect 58575 44693 58584 44727
rect 58532 44684 58584 44693
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 3056 44523 3108 44532
rect 3056 44489 3065 44523
rect 3065 44489 3099 44523
rect 3099 44489 3108 44523
rect 3056 44480 3108 44489
rect 7656 44480 7708 44532
rect 9588 44523 9640 44532
rect 9588 44489 9597 44523
rect 9597 44489 9631 44523
rect 9631 44489 9640 44523
rect 9588 44480 9640 44489
rect 12900 44523 12952 44532
rect 12900 44489 12909 44523
rect 12909 44489 12943 44523
rect 12943 44489 12952 44523
rect 12900 44480 12952 44489
rect 23112 44480 23164 44532
rect 31484 44480 31536 44532
rect 54024 44480 54076 44532
rect 55956 44523 56008 44532
rect 55956 44489 55965 44523
rect 55965 44489 55999 44523
rect 55999 44489 56008 44523
rect 55956 44480 56008 44489
rect 1676 44387 1728 44396
rect 1676 44353 1685 44387
rect 1685 44353 1719 44387
rect 1719 44353 1728 44387
rect 1676 44344 1728 44353
rect 3056 44344 3108 44396
rect 5356 44344 5408 44396
rect 7196 44412 7248 44464
rect 7472 44344 7524 44396
rect 10416 44412 10468 44464
rect 12164 44412 12216 44464
rect 15476 44412 15528 44464
rect 18236 44412 18288 44464
rect 30288 44412 30340 44464
rect 30380 44412 30432 44464
rect 33784 44455 33836 44464
rect 33784 44421 33818 44455
rect 33818 44421 33836 44455
rect 33784 44412 33836 44421
rect 43812 44412 43864 44464
rect 45744 44412 45796 44464
rect 10784 44344 10836 44396
rect 13636 44387 13688 44396
rect 13636 44353 13645 44387
rect 13645 44353 13679 44387
rect 13679 44353 13688 44387
rect 13636 44344 13688 44353
rect 16672 44344 16724 44396
rect 21824 44387 21876 44396
rect 21824 44353 21833 44387
rect 21833 44353 21867 44387
rect 21867 44353 21876 44387
rect 21824 44344 21876 44353
rect 23848 44344 23900 44396
rect 25044 44387 25096 44396
rect 25044 44353 25053 44387
rect 25053 44353 25087 44387
rect 25087 44353 25096 44387
rect 25044 44344 25096 44353
rect 27068 44344 27120 44396
rect 32220 44344 32272 44396
rect 6368 44319 6420 44328
rect 6368 44285 6377 44319
rect 6377 44285 6411 44319
rect 6411 44285 6420 44319
rect 6368 44276 6420 44285
rect 9496 44276 9548 44328
rect 11428 44276 11480 44328
rect 27712 44276 27764 44328
rect 32772 44276 32824 44328
rect 35440 44344 35492 44396
rect 36636 44344 36688 44396
rect 41788 44344 41840 44396
rect 42432 44344 42484 44396
rect 44456 44344 44508 44396
rect 46664 44344 46716 44396
rect 48964 44412 49016 44464
rect 53748 44412 53800 44464
rect 55036 44412 55088 44464
rect 48320 44344 48372 44396
rect 37924 44276 37976 44328
rect 40408 44276 40460 44328
rect 45284 44276 45336 44328
rect 52736 44387 52788 44396
rect 52736 44353 52745 44387
rect 52745 44353 52779 44387
rect 52779 44353 52788 44387
rect 52736 44344 52788 44353
rect 53288 44344 53340 44396
rect 54576 44387 54628 44396
rect 54576 44353 54585 44387
rect 54585 44353 54619 44387
rect 54619 44353 54628 44387
rect 54576 44344 54628 44353
rect 49424 44319 49476 44328
rect 49424 44285 49433 44319
rect 49433 44285 49467 44319
rect 49467 44285 49476 44319
rect 49424 44276 49476 44285
rect 5724 44183 5776 44192
rect 5724 44149 5733 44183
rect 5733 44149 5767 44183
rect 5767 44149 5776 44183
rect 5724 44140 5776 44149
rect 14372 44140 14424 44192
rect 18328 44183 18380 44192
rect 18328 44149 18337 44183
rect 18337 44149 18371 44183
rect 18371 44149 18380 44183
rect 18328 44140 18380 44149
rect 26424 44183 26476 44192
rect 26424 44149 26433 44183
rect 26433 44149 26467 44183
rect 26467 44149 26476 44183
rect 26424 44140 26476 44149
rect 29736 44183 29788 44192
rect 29736 44149 29745 44183
rect 29745 44149 29779 44183
rect 29779 44149 29788 44183
rect 29736 44140 29788 44149
rect 33324 44140 33376 44192
rect 36360 44140 36412 44192
rect 40040 44183 40092 44192
rect 40040 44149 40049 44183
rect 40049 44149 40083 44183
rect 40083 44149 40092 44183
rect 40040 44140 40092 44149
rect 40776 44140 40828 44192
rect 42800 44140 42852 44192
rect 47860 44140 47912 44192
rect 49700 44140 49752 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 6368 43936 6420 43988
rect 6828 43936 6880 43988
rect 23848 43979 23900 43988
rect 23848 43945 23857 43979
rect 23857 43945 23891 43979
rect 23891 43945 23900 43979
rect 23848 43936 23900 43945
rect 27068 43979 27120 43988
rect 27068 43945 27077 43979
rect 27077 43945 27111 43979
rect 27111 43945 27120 43979
rect 27068 43936 27120 43945
rect 27528 43936 27580 43988
rect 32220 43979 32272 43988
rect 32220 43945 32229 43979
rect 32229 43945 32263 43979
rect 32263 43945 32272 43979
rect 32220 43936 32272 43945
rect 35440 43936 35492 43988
rect 39212 43936 39264 43988
rect 42708 43936 42760 43988
rect 1676 43800 1728 43852
rect 14096 43843 14148 43852
rect 14096 43809 14105 43843
rect 14105 43809 14139 43843
rect 14139 43809 14148 43843
rect 14096 43800 14148 43809
rect 16672 43800 16724 43852
rect 17132 43843 17184 43852
rect 17132 43809 17141 43843
rect 17141 43809 17175 43843
rect 17175 43809 17184 43843
rect 17132 43800 17184 43809
rect 25044 43800 25096 43852
rect 25596 43800 25648 43852
rect 30380 43800 30432 43852
rect 45652 43936 45704 43988
rect 46664 43979 46716 43988
rect 46664 43945 46673 43979
rect 46673 43945 46707 43979
rect 46707 43945 46716 43979
rect 46664 43936 46716 43945
rect 53380 43979 53432 43988
rect 53380 43945 53389 43979
rect 53389 43945 53423 43979
rect 53423 43945 53432 43979
rect 53380 43936 53432 43945
rect 44456 43911 44508 43920
rect 44456 43877 44465 43911
rect 44465 43877 44499 43911
rect 44499 43877 44508 43911
rect 44456 43868 44508 43877
rect 56508 43843 56560 43852
rect 7748 43732 7800 43784
rect 9588 43775 9640 43784
rect 9588 43741 9597 43775
rect 9597 43741 9631 43775
rect 9631 43741 9640 43775
rect 9588 43732 9640 43741
rect 11428 43732 11480 43784
rect 14372 43775 14424 43784
rect 14372 43741 14406 43775
rect 14406 43741 14424 43775
rect 14372 43732 14424 43741
rect 18328 43732 18380 43784
rect 21548 43732 21600 43784
rect 27160 43732 27212 43784
rect 29184 43732 29236 43784
rect 5632 43707 5684 43716
rect 5632 43673 5641 43707
rect 5641 43673 5675 43707
rect 5675 43673 5684 43707
rect 5632 43664 5684 43673
rect 9680 43664 9732 43716
rect 10876 43664 10928 43716
rect 14832 43664 14884 43716
rect 20536 43664 20588 43716
rect 23204 43664 23256 43716
rect 27712 43664 27764 43716
rect 56508 43809 56517 43843
rect 56517 43809 56551 43843
rect 56551 43809 56560 43843
rect 56508 43800 56560 43809
rect 31944 43732 31996 43784
rect 32772 43775 32824 43784
rect 32772 43741 32781 43775
rect 32781 43741 32815 43775
rect 32815 43741 32824 43775
rect 32772 43732 32824 43741
rect 33324 43732 33376 43784
rect 37372 43732 37424 43784
rect 37924 43775 37976 43784
rect 37924 43741 37933 43775
rect 37933 43741 37967 43775
rect 37967 43741 37976 43775
rect 37924 43732 37976 43741
rect 39304 43732 39356 43784
rect 40500 43732 40552 43784
rect 42800 43732 42852 43784
rect 44456 43732 44508 43784
rect 45284 43775 45336 43784
rect 45284 43741 45293 43775
rect 45293 43741 45327 43775
rect 45327 43741 45336 43775
rect 45284 43732 45336 43741
rect 32956 43664 33008 43716
rect 39212 43664 39264 43716
rect 47124 43732 47176 43784
rect 46480 43664 46532 43716
rect 47952 43664 48004 43716
rect 49608 43664 49660 43716
rect 51632 43664 51684 43716
rect 52092 43732 52144 43784
rect 58532 43732 58584 43784
rect 53288 43664 53340 43716
rect 3240 43639 3292 43648
rect 3240 43605 3249 43639
rect 3249 43605 3283 43639
rect 3283 43605 3292 43639
rect 3240 43596 3292 43605
rect 11520 43596 11572 43648
rect 13544 43639 13596 43648
rect 13544 43605 13553 43639
rect 13553 43605 13587 43639
rect 13587 43605 13596 43639
rect 13544 43596 13596 43605
rect 15476 43639 15528 43648
rect 15476 43605 15485 43639
rect 15485 43605 15519 43639
rect 15519 43605 15528 43639
rect 15476 43596 15528 43605
rect 18512 43639 18564 43648
rect 18512 43605 18521 43639
rect 18521 43605 18555 43639
rect 18555 43605 18564 43639
rect 18512 43596 18564 43605
rect 21548 43639 21600 43648
rect 21548 43605 21557 43639
rect 21557 43605 21591 43639
rect 21591 43605 21600 43639
rect 21548 43596 21600 43605
rect 34152 43639 34204 43648
rect 34152 43605 34161 43639
rect 34161 43605 34195 43639
rect 34195 43605 34204 43639
rect 34152 43596 34204 43605
rect 48320 43596 48372 43648
rect 49424 43596 49476 43648
rect 51540 43639 51592 43648
rect 51540 43605 51549 43639
rect 51549 43605 51583 43639
rect 51583 43605 51592 43639
rect 51540 43596 51592 43605
rect 57888 43639 57940 43648
rect 57888 43605 57897 43639
rect 57897 43605 57931 43639
rect 57931 43605 57940 43639
rect 57888 43596 57940 43605
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 3056 43435 3108 43444
rect 3056 43401 3065 43435
rect 3065 43401 3099 43435
rect 3099 43401 3108 43435
rect 3056 43392 3108 43401
rect 5356 43435 5408 43444
rect 5356 43401 5365 43435
rect 5365 43401 5399 43435
rect 5399 43401 5408 43435
rect 5356 43392 5408 43401
rect 7472 43392 7524 43444
rect 14832 43435 14884 43444
rect 14832 43401 14841 43435
rect 14841 43401 14875 43435
rect 14875 43401 14884 43435
rect 14832 43392 14884 43401
rect 20536 43392 20588 43444
rect 23204 43435 23256 43444
rect 3240 43324 3292 43376
rect 5724 43324 5776 43376
rect 6828 43324 6880 43376
rect 15476 43324 15528 43376
rect 18512 43324 18564 43376
rect 1676 43299 1728 43308
rect 1676 43265 1685 43299
rect 1685 43265 1719 43299
rect 1719 43265 1728 43299
rect 1676 43256 1728 43265
rect 5172 43256 5224 43308
rect 22652 43324 22704 43376
rect 23204 43401 23213 43435
rect 23213 43401 23247 43435
rect 23247 43401 23256 43435
rect 23204 43392 23256 43401
rect 25596 43392 25648 43444
rect 30104 43392 30156 43444
rect 34796 43392 34848 43444
rect 35348 43392 35400 43444
rect 38016 43392 38068 43444
rect 46480 43435 46532 43444
rect 46480 43401 46489 43435
rect 46489 43401 46523 43435
rect 46523 43401 46532 43435
rect 46480 43392 46532 43401
rect 49608 43435 49660 43444
rect 49608 43401 49617 43435
rect 49617 43401 49651 43435
rect 49651 43401 49660 43435
rect 49608 43392 49660 43401
rect 54576 43435 54628 43444
rect 54576 43401 54585 43435
rect 54585 43401 54619 43435
rect 54619 43401 54628 43435
rect 54576 43392 54628 43401
rect 27344 43324 27396 43376
rect 10968 43256 11020 43308
rect 13360 43256 13412 43308
rect 14096 43256 14148 43308
rect 17132 43256 17184 43308
rect 19248 43299 19300 43308
rect 19248 43265 19257 43299
rect 19257 43265 19291 43299
rect 19291 43265 19300 43299
rect 19248 43256 19300 43265
rect 19340 43256 19392 43308
rect 21824 43299 21876 43308
rect 21824 43265 21833 43299
rect 21833 43265 21867 43299
rect 21867 43265 21876 43299
rect 21824 43256 21876 43265
rect 23664 43256 23716 43308
rect 27712 43324 27764 43376
rect 28908 43256 28960 43308
rect 29736 43324 29788 43376
rect 36728 43324 36780 43376
rect 39396 43324 39448 43376
rect 46204 43324 46256 43376
rect 49700 43324 49752 43376
rect 51540 43324 51592 43376
rect 32772 43256 32824 43308
rect 39212 43299 39264 43308
rect 39212 43265 39221 43299
rect 39221 43265 39255 43299
rect 39255 43265 39264 43299
rect 39212 43256 39264 43265
rect 40316 43256 40368 43308
rect 45192 43256 45244 43308
rect 46388 43256 46440 43308
rect 48320 43256 48372 43308
rect 49424 43256 49476 43308
rect 53104 43299 53156 43308
rect 53104 43265 53113 43299
rect 53113 43265 53147 43299
rect 53147 43265 53156 43299
rect 53104 43256 53156 43265
rect 55588 43256 55640 43308
rect 56508 43324 56560 43376
rect 58164 43256 58216 43308
rect 3792 43188 3844 43240
rect 9588 43231 9640 43240
rect 9588 43197 9597 43231
rect 9597 43197 9631 43231
rect 9631 43197 9640 43231
rect 9588 43188 9640 43197
rect 11428 43188 11480 43240
rect 37372 43231 37424 43240
rect 37372 43197 37381 43231
rect 37381 43197 37415 43231
rect 37415 43197 37424 43231
rect 37372 43188 37424 43197
rect 42432 43231 42484 43240
rect 42432 43197 42441 43231
rect 42441 43197 42475 43231
rect 42475 43197 42484 43231
rect 42432 43188 42484 43197
rect 36636 43120 36688 43172
rect 9496 43052 9548 43104
rect 12624 43052 12676 43104
rect 18604 43095 18656 43104
rect 18604 43061 18613 43095
rect 18613 43061 18647 43095
rect 18647 43061 18656 43095
rect 18604 43052 18656 43061
rect 18788 43052 18840 43104
rect 27436 43052 27488 43104
rect 40500 43095 40552 43104
rect 40500 43061 40509 43095
rect 40509 43061 40543 43095
rect 40543 43061 40552 43095
rect 40500 43052 40552 43061
rect 43076 43052 43128 43104
rect 51448 43095 51500 43104
rect 51448 43061 51457 43095
rect 51457 43061 51491 43095
rect 51491 43061 51500 43095
rect 51448 43052 51500 43061
rect 57336 43095 57388 43104
rect 57336 43061 57345 43095
rect 57345 43061 57379 43095
rect 57379 43061 57388 43095
rect 57336 43052 57388 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 5172 42891 5224 42900
rect 5172 42857 5181 42891
rect 5181 42857 5215 42891
rect 5215 42857 5224 42891
rect 5172 42848 5224 42857
rect 11428 42848 11480 42900
rect 23664 42891 23716 42900
rect 23664 42857 23673 42891
rect 23673 42857 23707 42891
rect 23707 42857 23716 42891
rect 23664 42848 23716 42857
rect 42524 42848 42576 42900
rect 44456 42848 44508 42900
rect 46388 42891 46440 42900
rect 46388 42857 46397 42891
rect 46397 42857 46431 42891
rect 46431 42857 46440 42891
rect 46388 42848 46440 42857
rect 19248 42780 19300 42832
rect 6828 42712 6880 42764
rect 17132 42712 17184 42764
rect 19984 42712 20036 42764
rect 48320 42848 48372 42900
rect 58164 42891 58216 42900
rect 58164 42857 58173 42891
rect 58173 42857 58207 42891
rect 58207 42857 58216 42891
rect 58164 42848 58216 42857
rect 9680 42644 9732 42696
rect 11336 42644 11388 42696
rect 15292 42644 15344 42696
rect 18604 42644 18656 42696
rect 49424 42712 49476 42764
rect 53288 42712 53340 42764
rect 56508 42712 56560 42764
rect 21548 42644 21600 42696
rect 22008 42644 22060 42696
rect 5172 42576 5224 42628
rect 8300 42576 8352 42628
rect 16028 42576 16080 42628
rect 21272 42576 21324 42628
rect 7656 42508 7708 42560
rect 16856 42551 16908 42560
rect 16856 42517 16865 42551
rect 16865 42517 16899 42551
rect 16899 42517 16908 42551
rect 16856 42508 16908 42517
rect 18696 42551 18748 42560
rect 18696 42517 18705 42551
rect 18705 42517 18739 42551
rect 18739 42517 18748 42551
rect 18696 42508 18748 42517
rect 22652 42576 22704 42628
rect 26424 42644 26476 42696
rect 27344 42576 27396 42628
rect 31576 42644 31628 42696
rect 32772 42644 32824 42696
rect 34152 42644 34204 42696
rect 32128 42576 32180 42628
rect 34704 42576 34756 42628
rect 36360 42644 36412 42696
rect 37372 42644 37424 42696
rect 37832 42644 37884 42696
rect 40040 42644 40092 42696
rect 40408 42644 40460 42696
rect 40776 42687 40828 42696
rect 40776 42653 40810 42687
rect 40810 42653 40828 42687
rect 40776 42644 40828 42653
rect 42432 42644 42484 42696
rect 44456 42644 44508 42696
rect 47860 42687 47912 42696
rect 47860 42653 47894 42687
rect 47894 42653 47912 42687
rect 47860 42644 47912 42653
rect 51448 42644 51500 42696
rect 57888 42644 57940 42696
rect 43812 42576 43864 42628
rect 46756 42576 46808 42628
rect 55128 42576 55180 42628
rect 25780 42551 25832 42560
rect 25780 42517 25789 42551
rect 25789 42517 25823 42551
rect 25823 42517 25832 42551
rect 25780 42508 25832 42517
rect 27712 42508 27764 42560
rect 32036 42508 32088 42560
rect 34060 42551 34112 42560
rect 34060 42517 34069 42551
rect 34069 42517 34103 42551
rect 34103 42517 34112 42551
rect 34060 42508 34112 42517
rect 36544 42508 36596 42560
rect 39120 42508 39172 42560
rect 40040 42508 40092 42560
rect 41880 42551 41932 42560
rect 41880 42517 41889 42551
rect 41889 42517 41923 42551
rect 41923 42517 41932 42551
rect 41880 42508 41932 42517
rect 45100 42508 45152 42560
rect 48872 42508 48924 42560
rect 51356 42508 51408 42560
rect 54760 42551 54812 42560
rect 54760 42517 54769 42551
rect 54769 42517 54803 42551
rect 54803 42517 54812 42551
rect 54760 42508 54812 42517
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 10968 42347 11020 42356
rect 10968 42313 10977 42347
rect 10977 42313 11011 42347
rect 11011 42313 11020 42347
rect 10968 42304 11020 42313
rect 13360 42304 13412 42356
rect 19340 42304 19392 42356
rect 21272 42347 21324 42356
rect 21272 42313 21281 42347
rect 21281 42313 21315 42347
rect 21315 42313 21324 42347
rect 21272 42304 21324 42313
rect 24952 42304 25004 42356
rect 28908 42304 28960 42356
rect 44456 42347 44508 42356
rect 44456 42313 44465 42347
rect 44465 42313 44499 42347
rect 44499 42313 44508 42347
rect 44456 42304 44508 42313
rect 46756 42347 46808 42356
rect 46756 42313 46765 42347
rect 46765 42313 46799 42347
rect 46799 42313 46808 42347
rect 46756 42304 46808 42313
rect 55128 42347 55180 42356
rect 55128 42313 55137 42347
rect 55137 42313 55171 42347
rect 55171 42313 55180 42347
rect 55128 42304 55180 42313
rect 56508 42304 56560 42356
rect 12808 42236 12860 42288
rect 13544 42236 13596 42288
rect 18696 42236 18748 42288
rect 25688 42236 25740 42288
rect 5448 42168 5500 42220
rect 6828 42168 6880 42220
rect 11612 42168 11664 42220
rect 14096 42168 14148 42220
rect 18604 42168 18656 42220
rect 19984 42168 20036 42220
rect 21548 42168 21600 42220
rect 22652 42211 22704 42220
rect 22652 42177 22661 42211
rect 22661 42177 22695 42211
rect 22695 42177 22704 42211
rect 22652 42168 22704 42177
rect 26148 42168 26200 42220
rect 29000 42168 29052 42220
rect 34244 42168 34296 42220
rect 37832 42168 37884 42220
rect 40224 42168 40276 42220
rect 40408 42168 40460 42220
rect 45192 42168 45244 42220
rect 46388 42168 46440 42220
rect 48320 42168 48372 42220
rect 50160 42168 50212 42220
rect 51632 42236 51684 42288
rect 55588 42279 55640 42288
rect 55588 42245 55597 42279
rect 55597 42245 55631 42279
rect 55631 42245 55640 42279
rect 55588 42236 55640 42245
rect 53656 42168 53708 42220
rect 56232 42168 56284 42220
rect 8944 42100 8996 42152
rect 9588 42143 9640 42152
rect 9588 42109 9597 42143
rect 9597 42109 9631 42143
rect 9631 42109 9640 42143
rect 9588 42100 9640 42109
rect 17316 42100 17368 42152
rect 27712 42143 27764 42152
rect 27712 42109 27721 42143
rect 27721 42109 27755 42143
rect 27755 42109 27764 42143
rect 27712 42100 27764 42109
rect 34704 42143 34756 42152
rect 34704 42109 34713 42143
rect 34713 42109 34747 42143
rect 34747 42109 34756 42143
rect 34704 42100 34756 42109
rect 53380 42100 53432 42152
rect 3792 41964 3844 42016
rect 4068 41964 4120 42016
rect 8576 42007 8628 42016
rect 8576 41973 8585 42007
rect 8585 41973 8619 42007
rect 8619 41973 8628 42007
rect 8576 41964 8628 41973
rect 16120 42007 16172 42016
rect 16120 41973 16129 42007
rect 16129 41973 16163 42007
rect 16163 41973 16172 42007
rect 16120 41964 16172 41973
rect 25872 42007 25924 42016
rect 25872 41973 25881 42007
rect 25881 41973 25915 42007
rect 25915 41973 25924 42007
rect 25872 41964 25924 41973
rect 36084 42007 36136 42016
rect 36084 41973 36093 42007
rect 36093 41973 36127 42007
rect 36127 41973 36136 42007
rect 36084 41964 36136 41973
rect 40316 41964 40368 42016
rect 49700 41964 49752 42016
rect 52184 42007 52236 42016
rect 52184 41973 52193 42007
rect 52193 41973 52227 42007
rect 52227 41973 52236 42007
rect 52184 41964 52236 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 5172 41803 5224 41812
rect 5172 41769 5181 41803
rect 5181 41769 5215 41803
rect 5215 41769 5224 41803
rect 5172 41760 5224 41769
rect 8300 41760 8352 41812
rect 11612 41803 11664 41812
rect 11612 41769 11621 41803
rect 11621 41769 11655 41803
rect 11655 41769 11664 41803
rect 11612 41760 11664 41769
rect 21548 41803 21600 41812
rect 11336 41692 11388 41744
rect 6828 41624 6880 41676
rect 11428 41624 11480 41676
rect 3792 41599 3844 41608
rect 3792 41565 3801 41599
rect 3801 41565 3835 41599
rect 3835 41565 3844 41599
rect 3792 41556 3844 41565
rect 4068 41599 4120 41608
rect 4068 41565 4102 41599
rect 4102 41565 4120 41599
rect 4068 41556 4120 41565
rect 8576 41556 8628 41608
rect 12624 41556 12676 41608
rect 21548 41769 21557 41803
rect 21557 41769 21591 41803
rect 21591 41769 21600 41803
rect 21548 41760 21600 41769
rect 29000 41803 29052 41812
rect 29000 41769 29009 41803
rect 29009 41769 29043 41803
rect 29043 41769 29052 41803
rect 29000 41760 29052 41769
rect 41788 41760 41840 41812
rect 43812 41803 43864 41812
rect 43812 41769 43821 41803
rect 43821 41769 43855 41803
rect 43855 41769 43864 41803
rect 43812 41760 43864 41769
rect 19984 41624 20036 41676
rect 22008 41624 22060 41676
rect 34704 41624 34756 41676
rect 35348 41667 35400 41676
rect 35348 41633 35357 41667
rect 35357 41633 35391 41667
rect 35391 41633 35400 41667
rect 35348 41624 35400 41633
rect 45192 41760 45244 41812
rect 46388 41803 46440 41812
rect 46388 41769 46397 41803
rect 46397 41769 46431 41803
rect 46431 41769 46440 41803
rect 46388 41760 46440 41769
rect 17316 41599 17368 41608
rect 17316 41565 17325 41599
rect 17325 41565 17359 41599
rect 17359 41565 17368 41599
rect 17316 41556 17368 41565
rect 18788 41556 18840 41608
rect 24952 41556 25004 41608
rect 12164 41420 12216 41472
rect 21272 41488 21324 41540
rect 23756 41488 23808 41540
rect 27436 41556 27488 41608
rect 27712 41556 27764 41608
rect 30196 41556 30248 41608
rect 32128 41599 32180 41608
rect 32128 41565 32137 41599
rect 32137 41565 32171 41599
rect 32171 41565 32180 41599
rect 32128 41556 32180 41565
rect 37832 41599 37884 41608
rect 37832 41565 37841 41599
rect 37841 41565 37875 41599
rect 37875 41565 37884 41599
rect 40500 41599 40552 41608
rect 37832 41556 37884 41565
rect 40500 41565 40509 41599
rect 40509 41565 40543 41599
rect 40543 41565 40552 41599
rect 40500 41556 40552 41565
rect 41052 41556 41104 41608
rect 42432 41599 42484 41608
rect 42432 41565 42441 41599
rect 42441 41565 42475 41599
rect 42475 41565 42484 41599
rect 42432 41556 42484 41565
rect 48320 41556 48372 41608
rect 51080 41556 51132 41608
rect 51632 41556 51684 41608
rect 52736 41556 52788 41608
rect 53380 41599 53432 41608
rect 53380 41565 53389 41599
rect 53389 41565 53423 41599
rect 53423 41565 53432 41599
rect 53380 41556 53432 41565
rect 54760 41556 54812 41608
rect 29644 41488 29696 41540
rect 31116 41488 31168 41540
rect 32404 41531 32456 41540
rect 32404 41497 32438 41531
rect 32438 41497 32456 41531
rect 32404 41488 32456 41497
rect 36544 41488 36596 41540
rect 39120 41488 39172 41540
rect 43720 41488 43772 41540
rect 46572 41488 46624 41540
rect 49332 41488 49384 41540
rect 53748 41488 53800 41540
rect 55680 41488 55732 41540
rect 57336 41556 57388 41608
rect 56508 41488 56560 41540
rect 14096 41420 14148 41472
rect 18696 41463 18748 41472
rect 18696 41429 18705 41463
rect 18705 41429 18739 41463
rect 18739 41429 18748 41463
rect 18696 41420 18748 41429
rect 23204 41420 23256 41472
rect 26608 41420 26660 41472
rect 30380 41420 30432 41472
rect 32036 41420 32088 41472
rect 36268 41420 36320 41472
rect 37740 41420 37792 41472
rect 49056 41463 49108 41472
rect 49056 41429 49065 41463
rect 49065 41429 49099 41463
rect 49099 41429 49108 41463
rect 49056 41420 49108 41429
rect 52920 41463 52972 41472
rect 52920 41429 52929 41463
rect 52929 41429 52963 41463
rect 52963 41429 52972 41463
rect 52920 41420 52972 41429
rect 54760 41463 54812 41472
rect 54760 41429 54769 41463
rect 54769 41429 54803 41463
rect 54803 41429 54812 41463
rect 54760 41420 54812 41429
rect 57336 41463 57388 41472
rect 57336 41429 57345 41463
rect 57345 41429 57379 41463
rect 57379 41429 57388 41463
rect 57336 41420 57388 41429
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 5448 41259 5500 41268
rect 5448 41225 5457 41259
rect 5457 41225 5491 41259
rect 5491 41225 5500 41259
rect 5448 41216 5500 41225
rect 21272 41259 21324 41268
rect 21272 41225 21281 41259
rect 21281 41225 21315 41259
rect 21315 41225 21324 41259
rect 21272 41216 21324 41225
rect 29644 41259 29696 41268
rect 29644 41225 29653 41259
rect 29653 41225 29687 41259
rect 29687 41225 29696 41259
rect 29644 41216 29696 41225
rect 36544 41216 36596 41268
rect 43720 41216 43772 41268
rect 46572 41259 46624 41268
rect 46572 41225 46581 41259
rect 46581 41225 46615 41259
rect 46615 41225 46624 41259
rect 46572 41216 46624 41225
rect 50160 41216 50212 41268
rect 53748 41216 53800 41268
rect 3240 41080 3292 41132
rect 7656 41148 7708 41200
rect 9496 41191 9548 41200
rect 9496 41157 9530 41191
rect 9530 41157 9548 41191
rect 9496 41148 9548 41157
rect 12164 41080 12216 41132
rect 14096 41148 14148 41200
rect 16120 41148 16172 41200
rect 18696 41148 18748 41200
rect 25872 41148 25924 41200
rect 52184 41148 52236 41200
rect 54760 41148 54812 41200
rect 57336 41148 57388 41200
rect 14832 41080 14884 41132
rect 19984 41080 20036 41132
rect 21272 41080 21324 41132
rect 22652 41080 22704 41132
rect 27160 41080 27212 41132
rect 29000 41080 29052 41132
rect 31576 41080 31628 41132
rect 34060 41080 34112 41132
rect 35348 41123 35400 41132
rect 35348 41089 35357 41123
rect 35357 41089 35391 41123
rect 35391 41089 35400 41123
rect 35348 41080 35400 41089
rect 36728 41080 36780 41132
rect 40592 41080 40644 41132
rect 41788 41080 41840 41132
rect 43812 41080 43864 41132
rect 45192 41123 45244 41132
rect 45192 41089 45201 41123
rect 45201 41089 45235 41123
rect 45235 41089 45244 41123
rect 45192 41080 45244 41089
rect 46848 41080 46900 41132
rect 48320 41080 48372 41132
rect 51540 41080 51592 41132
rect 55680 41123 55732 41132
rect 55680 41089 55689 41123
rect 55689 41089 55723 41123
rect 55723 41089 55732 41123
rect 55680 41080 55732 41089
rect 3792 41012 3844 41064
rect 6460 41055 6512 41064
rect 6460 41021 6469 41055
rect 6469 41021 6503 41055
rect 6503 41021 6512 41055
rect 6460 41012 6512 41021
rect 8944 41012 8996 41064
rect 14096 41012 14148 41064
rect 14740 41055 14792 41064
rect 14740 41021 14749 41055
rect 14749 41021 14783 41055
rect 14783 41021 14792 41055
rect 14740 41012 14792 41021
rect 17316 41012 17368 41064
rect 24952 41012 25004 41064
rect 27712 41012 27764 41064
rect 30196 41055 30248 41064
rect 30196 41021 30205 41055
rect 30205 41021 30239 41055
rect 30239 41021 30248 41055
rect 30196 41012 30248 41021
rect 32128 41012 32180 41064
rect 32496 41055 32548 41064
rect 32496 41021 32505 41055
rect 32505 41021 32539 41055
rect 32539 41021 32548 41055
rect 32496 41012 32548 41021
rect 16028 40944 16080 40996
rect 7840 40919 7892 40928
rect 7840 40885 7849 40919
rect 7849 40885 7883 40919
rect 7883 40885 7892 40919
rect 7840 40876 7892 40885
rect 10600 40919 10652 40928
rect 10600 40885 10609 40919
rect 10609 40885 10643 40919
rect 10643 40885 10652 40919
rect 10600 40876 10652 40885
rect 14280 40919 14332 40928
rect 14280 40885 14289 40919
rect 14289 40885 14323 40919
rect 14323 40885 14332 40919
rect 14280 40876 14332 40885
rect 19064 40919 19116 40928
rect 19064 40885 19073 40919
rect 19073 40885 19107 40919
rect 19107 40885 19116 40919
rect 19064 40876 19116 40885
rect 24584 40919 24636 40928
rect 24584 40885 24593 40919
rect 24593 40885 24627 40919
rect 24627 40885 24636 40919
rect 24584 40876 24636 40885
rect 26424 40919 26476 40928
rect 26424 40885 26433 40919
rect 26433 40885 26467 40919
rect 26467 40885 26476 40919
rect 26424 40876 26476 40885
rect 30012 40876 30064 40928
rect 31760 40876 31812 40928
rect 39948 41012 40000 41064
rect 42432 41055 42484 41064
rect 42432 41021 42441 41055
rect 42441 41021 42475 41055
rect 42475 41021 42484 41055
rect 42432 41012 42484 41021
rect 39396 40876 39448 40928
rect 40040 40919 40092 40928
rect 40040 40885 40049 40919
rect 40049 40885 40083 40919
rect 40083 40885 40092 40919
rect 40040 40876 40092 40885
rect 40132 40876 40184 40928
rect 52736 41012 52788 41064
rect 51080 40876 51132 40928
rect 52184 40919 52236 40928
rect 52184 40885 52193 40919
rect 52193 40885 52227 40919
rect 52227 40885 52236 40919
rect 52184 40876 52236 40885
rect 57060 40919 57112 40928
rect 57060 40885 57069 40919
rect 57069 40885 57103 40919
rect 57103 40885 57112 40919
rect 57060 40876 57112 40885
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 3240 40715 3292 40724
rect 3240 40681 3249 40715
rect 3249 40681 3283 40715
rect 3283 40681 3292 40715
rect 3240 40672 3292 40681
rect 10876 40672 10928 40724
rect 12808 40715 12860 40724
rect 12808 40681 12817 40715
rect 12817 40681 12851 40715
rect 12851 40681 12860 40715
rect 12808 40672 12860 40681
rect 18604 40672 18656 40724
rect 23756 40672 23808 40724
rect 27160 40715 27212 40724
rect 27160 40681 27169 40715
rect 27169 40681 27203 40715
rect 27203 40681 27212 40715
rect 27160 40672 27212 40681
rect 29000 40715 29052 40724
rect 29000 40681 29009 40715
rect 29009 40681 29043 40715
rect 29043 40681 29052 40715
rect 29000 40672 29052 40681
rect 30196 40672 30248 40724
rect 15292 40579 15344 40588
rect 15292 40545 15301 40579
rect 15301 40545 15335 40579
rect 15335 40545 15344 40579
rect 15292 40536 15344 40545
rect 24952 40536 25004 40588
rect 32128 40672 32180 40724
rect 41788 40715 41840 40724
rect 41788 40681 41797 40715
rect 41797 40681 41831 40715
rect 41831 40681 41840 40715
rect 41788 40672 41840 40681
rect 43812 40715 43864 40724
rect 43812 40681 43821 40715
rect 43821 40681 43855 40715
rect 43855 40681 43864 40715
rect 43812 40672 43864 40681
rect 2872 40468 2924 40520
rect 5816 40468 5868 40520
rect 7840 40468 7892 40520
rect 8944 40468 8996 40520
rect 10600 40468 10652 40520
rect 3240 40400 3292 40452
rect 11520 40468 11572 40520
rect 12164 40400 12216 40452
rect 16856 40468 16908 40520
rect 17316 40511 17368 40520
rect 17316 40477 17325 40511
rect 17325 40477 17359 40511
rect 17359 40477 17368 40511
rect 17316 40468 17368 40477
rect 19064 40468 19116 40520
rect 22560 40468 22612 40520
rect 24584 40468 24636 40520
rect 26608 40468 26660 40520
rect 27712 40468 27764 40520
rect 32036 40468 32088 40520
rect 35992 40468 36044 40520
rect 20536 40400 20588 40452
rect 29736 40400 29788 40452
rect 32312 40400 32364 40452
rect 32956 40400 33008 40452
rect 34336 40400 34388 40452
rect 37740 40468 37792 40520
rect 39396 40536 39448 40588
rect 39948 40536 40000 40588
rect 45192 40672 45244 40724
rect 46204 40672 46256 40724
rect 51080 40672 51132 40724
rect 53656 40715 53708 40724
rect 53656 40681 53665 40715
rect 53665 40681 53699 40715
rect 53699 40681 53708 40715
rect 53656 40672 53708 40681
rect 40040 40468 40092 40520
rect 51632 40536 51684 40588
rect 53380 40536 53432 40588
rect 55680 40672 55732 40724
rect 56232 40672 56284 40724
rect 42432 40511 42484 40520
rect 42432 40477 42441 40511
rect 42441 40477 42475 40511
rect 42475 40477 42484 40511
rect 42432 40468 42484 40477
rect 37832 40400 37884 40452
rect 43076 40468 43128 40520
rect 45100 40468 45152 40520
rect 48320 40468 48372 40520
rect 49700 40468 49752 40520
rect 52184 40468 52236 40520
rect 52920 40468 52972 40520
rect 57060 40468 57112 40520
rect 43720 40400 43772 40452
rect 7564 40375 7616 40384
rect 7564 40341 7573 40375
rect 7573 40341 7607 40375
rect 7607 40341 7616 40375
rect 7564 40332 7616 40341
rect 15292 40332 15344 40384
rect 21088 40375 21140 40384
rect 21088 40341 21097 40375
rect 21097 40341 21131 40375
rect 21131 40341 21140 40375
rect 21088 40332 21140 40341
rect 31944 40375 31996 40384
rect 31944 40341 31953 40375
rect 31953 40341 31987 40375
rect 31987 40341 31996 40375
rect 31944 40332 31996 40341
rect 37464 40375 37516 40384
rect 37464 40341 37473 40375
rect 37473 40341 37507 40375
rect 37507 40341 37516 40375
rect 37464 40332 37516 40341
rect 39304 40375 39356 40384
rect 39304 40341 39313 40375
rect 39313 40341 39347 40375
rect 39347 40341 39356 40375
rect 39304 40332 39356 40341
rect 49608 40375 49660 40384
rect 49608 40341 49617 40375
rect 49617 40341 49651 40375
rect 49651 40341 49660 40375
rect 49608 40332 49660 40341
rect 51816 40375 51868 40384
rect 51816 40341 51825 40375
rect 51825 40341 51859 40375
rect 51859 40341 51868 40375
rect 51816 40332 51868 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 19340 40128 19392 40180
rect 21272 40171 21324 40180
rect 21272 40137 21281 40171
rect 21281 40137 21315 40171
rect 21315 40137 21324 40171
rect 21272 40128 21324 40137
rect 26148 40171 26200 40180
rect 26148 40137 26157 40171
rect 26157 40137 26191 40171
rect 26191 40137 26200 40171
rect 26148 40128 26200 40137
rect 29736 40171 29788 40180
rect 29736 40137 29745 40171
rect 29745 40137 29779 40171
rect 29779 40137 29788 40171
rect 29736 40128 29788 40137
rect 31576 40171 31628 40180
rect 31576 40137 31585 40171
rect 31585 40137 31619 40171
rect 31619 40137 31628 40171
rect 31576 40128 31628 40137
rect 36728 40171 36780 40180
rect 36728 40137 36737 40171
rect 36737 40137 36771 40171
rect 36771 40137 36780 40171
rect 36728 40128 36780 40137
rect 40592 40128 40644 40180
rect 43720 40128 43772 40180
rect 51540 40171 51592 40180
rect 51540 40137 51549 40171
rect 51549 40137 51583 40171
rect 51583 40137 51592 40171
rect 51540 40128 51592 40137
rect 2872 40060 2924 40112
rect 3792 40060 3844 40112
rect 5632 40060 5684 40112
rect 3976 39992 4028 40044
rect 5816 39967 5868 39976
rect 5816 39933 5825 39967
rect 5825 39933 5859 39967
rect 5859 39933 5868 39967
rect 5816 39924 5868 39933
rect 3608 39831 3660 39840
rect 3608 39797 3617 39831
rect 3617 39797 3651 39831
rect 3651 39797 3660 39831
rect 3608 39788 3660 39797
rect 6460 39992 6512 40044
rect 7564 39992 7616 40044
rect 7840 39992 7892 40044
rect 12164 40035 12216 40044
rect 12164 40001 12173 40035
rect 12173 40001 12207 40035
rect 12207 40001 12216 40035
rect 12164 39992 12216 40001
rect 14280 39992 14332 40044
rect 14740 40035 14792 40044
rect 14740 40001 14749 40035
rect 14749 40001 14783 40035
rect 14783 40001 14792 40035
rect 14740 39992 14792 40001
rect 15292 39992 15344 40044
rect 17316 40060 17368 40112
rect 24952 40060 25004 40112
rect 32496 40060 32548 40112
rect 18052 39992 18104 40044
rect 19984 39992 20036 40044
rect 23020 39992 23072 40044
rect 23204 40035 23256 40044
rect 23204 40001 23238 40035
rect 23238 40001 23256 40035
rect 23204 39992 23256 40001
rect 34336 40060 34388 40112
rect 26424 39992 26476 40044
rect 27712 39992 27764 40044
rect 30288 39992 30340 40044
rect 31576 39992 31628 40044
rect 32772 40035 32824 40044
rect 32772 40001 32781 40035
rect 32781 40001 32815 40035
rect 32815 40001 32824 40035
rect 32772 39992 32824 40001
rect 8208 39967 8260 39976
rect 8208 39933 8217 39967
rect 8217 39933 8251 39967
rect 8251 39933 8260 39967
rect 8208 39924 8260 39933
rect 22560 39924 22612 39976
rect 30196 39967 30248 39976
rect 30196 39933 30205 39967
rect 30205 39933 30239 39967
rect 30239 39933 30248 39967
rect 30196 39924 30248 39933
rect 7748 39831 7800 39840
rect 7748 39797 7757 39831
rect 7757 39797 7791 39831
rect 7791 39797 7800 39831
rect 7748 39788 7800 39797
rect 8392 39788 8444 39840
rect 13544 39831 13596 39840
rect 13544 39797 13553 39831
rect 13553 39797 13587 39831
rect 13587 39797 13596 39831
rect 13544 39788 13596 39797
rect 16120 39831 16172 39840
rect 16120 39797 16129 39831
rect 16129 39797 16163 39831
rect 16163 39797 16172 39831
rect 16120 39788 16172 39797
rect 24308 39831 24360 39840
rect 24308 39797 24317 39831
rect 24317 39797 24351 39831
rect 24351 39797 24360 39831
rect 24308 39788 24360 39797
rect 34152 39831 34204 39840
rect 34152 39797 34161 39831
rect 34161 39797 34195 39831
rect 34195 39797 34204 39831
rect 34152 39788 34204 39797
rect 35992 40060 36044 40112
rect 47952 40103 48004 40112
rect 47952 40069 47961 40103
rect 47961 40069 47995 40103
rect 47995 40069 48004 40103
rect 47952 40060 48004 40069
rect 49792 40060 49844 40112
rect 37372 39992 37424 40044
rect 39396 40035 39448 40044
rect 36084 39788 36136 39840
rect 38752 39788 38804 39840
rect 38936 39831 38988 39840
rect 38936 39797 38945 39831
rect 38945 39797 38979 39831
rect 38979 39797 38988 39831
rect 38936 39788 38988 39797
rect 39396 40001 39405 40035
rect 39405 40001 39439 40035
rect 39439 40001 39448 40035
rect 39396 39992 39448 40001
rect 40132 39992 40184 40044
rect 42432 40035 42484 40044
rect 42432 40001 42441 40035
rect 42441 40001 42475 40035
rect 42475 40001 42484 40035
rect 42432 39992 42484 40001
rect 43812 39992 43864 40044
rect 45192 39992 45244 40044
rect 47768 39992 47820 40044
rect 51080 40060 51132 40112
rect 51816 39992 51868 40044
rect 40316 39788 40368 39840
rect 47032 39831 47084 39840
rect 47032 39797 47041 39831
rect 47041 39797 47075 39831
rect 47075 39797 47084 39831
rect 47032 39788 47084 39797
rect 48228 39788 48280 39840
rect 49792 39788 49844 39840
rect 53104 39788 53156 39840
rect 54668 39788 54720 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 3240 39627 3292 39636
rect 3240 39593 3249 39627
rect 3249 39593 3283 39627
rect 3283 39593 3292 39627
rect 3240 39584 3292 39593
rect 3976 39584 4028 39636
rect 7840 39584 7892 39636
rect 11336 39584 11388 39636
rect 18052 39627 18104 39636
rect 8300 39448 8352 39500
rect 8944 39491 8996 39500
rect 8944 39457 8953 39491
rect 8953 39457 8987 39491
rect 8987 39457 8996 39491
rect 8944 39448 8996 39457
rect 3608 39380 3660 39432
rect 3792 39423 3844 39432
rect 3792 39389 3801 39423
rect 3801 39389 3835 39423
rect 3835 39389 3844 39423
rect 3792 39380 3844 39389
rect 5816 39380 5868 39432
rect 4068 39355 4120 39364
rect 4068 39321 4102 39355
rect 4102 39321 4120 39355
rect 7748 39380 7800 39432
rect 4068 39312 4120 39321
rect 6828 39312 6880 39364
rect 8484 39312 8536 39364
rect 18052 39593 18061 39627
rect 18061 39593 18095 39627
rect 18095 39593 18104 39627
rect 18052 39584 18104 39593
rect 20812 39584 20864 39636
rect 29644 39584 29696 39636
rect 32404 39584 32456 39636
rect 34060 39584 34112 39636
rect 37372 39584 37424 39636
rect 39120 39584 39172 39636
rect 40408 39584 40460 39636
rect 43812 39627 43864 39636
rect 43812 39593 43821 39627
rect 43821 39593 43855 39627
rect 43855 39593 43864 39627
rect 43812 39584 43864 39593
rect 47768 39627 47820 39636
rect 47768 39593 47777 39627
rect 47777 39593 47811 39627
rect 47811 39593 47820 39627
rect 47768 39584 47820 39593
rect 12164 39491 12216 39500
rect 12164 39457 12173 39491
rect 12173 39457 12207 39491
rect 12207 39457 12216 39491
rect 12164 39448 12216 39457
rect 32772 39491 32824 39500
rect 32772 39457 32781 39491
rect 32781 39457 32815 39491
rect 32815 39457 32824 39491
rect 32772 39448 32824 39457
rect 34336 39448 34388 39500
rect 37832 39448 37884 39500
rect 42432 39491 42484 39500
rect 42432 39457 42441 39491
rect 42441 39457 42475 39491
rect 42475 39457 42484 39491
rect 42432 39448 42484 39457
rect 47952 39448 48004 39500
rect 48228 39491 48280 39500
rect 48228 39457 48237 39491
rect 48237 39457 48271 39491
rect 48271 39457 48280 39491
rect 48228 39448 48280 39457
rect 13544 39380 13596 39432
rect 13360 39312 13412 39364
rect 16120 39380 16172 39432
rect 17316 39380 17368 39432
rect 18512 39380 18564 39432
rect 19340 39380 19392 39432
rect 22560 39380 22612 39432
rect 24308 39380 24360 39432
rect 24400 39380 24452 39432
rect 30196 39380 30248 39432
rect 14740 39312 14792 39364
rect 18328 39312 18380 39364
rect 27528 39312 27580 39364
rect 30288 39312 30340 39364
rect 31760 39380 31812 39432
rect 34152 39380 34204 39432
rect 37464 39380 37516 39432
rect 38936 39380 38988 39432
rect 40316 39380 40368 39432
rect 40960 39380 41012 39432
rect 46204 39380 46256 39432
rect 49608 39380 49660 39432
rect 52736 39423 52788 39432
rect 52736 39389 52745 39423
rect 52745 39389 52779 39423
rect 52779 39389 52788 39423
rect 52736 39380 52788 39389
rect 53472 39380 53524 39432
rect 32772 39312 32824 39364
rect 43720 39312 43772 39364
rect 49056 39312 49108 39364
rect 52828 39312 52880 39364
rect 53012 39355 53064 39364
rect 53012 39321 53046 39355
rect 53046 39321 53064 39355
rect 53012 39312 53064 39321
rect 10324 39287 10376 39296
rect 10324 39253 10333 39287
rect 10333 39253 10367 39287
rect 10367 39253 10376 39287
rect 10324 39244 10376 39253
rect 13544 39287 13596 39296
rect 13544 39253 13553 39287
rect 13553 39253 13587 39287
rect 13587 39253 13596 39287
rect 13544 39244 13596 39253
rect 14832 39244 14884 39296
rect 20628 39287 20680 39296
rect 20628 39253 20637 39287
rect 20637 39253 20671 39287
rect 20671 39253 20680 39287
rect 20628 39244 20680 39253
rect 23848 39287 23900 39296
rect 23848 39253 23857 39287
rect 23857 39253 23891 39287
rect 23891 39253 23900 39287
rect 23848 39244 23900 39253
rect 27620 39244 27672 39296
rect 49608 39287 49660 39296
rect 49608 39253 49617 39287
rect 49617 39253 49651 39287
rect 49651 39253 49660 39287
rect 49608 39244 49660 39253
rect 52276 39287 52328 39296
rect 52276 39253 52285 39287
rect 52285 39253 52319 39287
rect 52319 39253 52328 39287
rect 52276 39244 52328 39253
rect 53932 39244 53984 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 8484 39083 8536 39092
rect 8484 39049 8493 39083
rect 8493 39049 8527 39083
rect 8527 39049 8536 39083
rect 8484 39040 8536 39049
rect 18328 39083 18380 39092
rect 18328 39049 18337 39083
rect 18337 39049 18371 39083
rect 18371 39049 18380 39083
rect 18328 39040 18380 39049
rect 23020 39040 23072 39092
rect 28448 39040 28500 39092
rect 31576 39083 31628 39092
rect 31576 39049 31585 39083
rect 31585 39049 31619 39083
rect 31619 39049 31628 39083
rect 31576 39040 31628 39049
rect 34244 39083 34296 39092
rect 34244 39049 34253 39083
rect 34253 39049 34287 39083
rect 34287 39049 34296 39083
rect 34244 39040 34296 39049
rect 40224 39083 40276 39092
rect 40224 39049 40233 39083
rect 40233 39049 40267 39083
rect 40267 39049 40276 39083
rect 40224 39040 40276 39049
rect 43720 39040 43772 39092
rect 49332 39083 49384 39092
rect 49332 39049 49341 39083
rect 49341 39049 49375 39083
rect 49375 39049 49384 39083
rect 49332 39040 49384 39049
rect 8392 38972 8444 39024
rect 10324 38972 10376 39024
rect 13544 38972 13596 39024
rect 20628 38972 20680 39024
rect 23848 38972 23900 39024
rect 5724 38904 5776 38956
rect 6828 38904 6880 38956
rect 8944 38947 8996 38956
rect 8944 38913 8953 38947
rect 8953 38913 8987 38947
rect 8987 38913 8996 38947
rect 8944 38904 8996 38913
rect 12164 38947 12216 38956
rect 12164 38913 12173 38947
rect 12173 38913 12207 38947
rect 12207 38913 12216 38947
rect 12164 38904 12216 38913
rect 18052 38904 18104 38956
rect 20812 38947 20864 38956
rect 20812 38913 20821 38947
rect 20821 38913 20855 38947
rect 20855 38913 20864 38947
rect 20812 38904 20864 38913
rect 24400 38904 24452 38956
rect 27712 38972 27764 39024
rect 31944 38972 31996 39024
rect 36268 38972 36320 39024
rect 39304 38972 39356 39024
rect 47032 38972 47084 39024
rect 49608 38972 49660 39024
rect 28540 38904 28592 38956
rect 30196 38947 30248 38956
rect 30196 38913 30205 38947
rect 30205 38913 30239 38947
rect 30239 38913 30248 38947
rect 30196 38904 30248 38913
rect 32772 38904 32824 38956
rect 36084 38904 36136 38956
rect 38752 38904 38804 38956
rect 43996 38904 44048 38956
rect 45192 38904 45244 38956
rect 46204 38904 46256 38956
rect 51540 38972 51592 39024
rect 52092 38904 52144 38956
rect 53472 38947 53524 38956
rect 53472 38913 53481 38947
rect 53481 38913 53515 38947
rect 53515 38913 53524 38947
rect 53472 38904 53524 38913
rect 56692 38904 56744 38956
rect 3792 38879 3844 38888
rect 3792 38845 3801 38879
rect 3801 38845 3835 38879
rect 3835 38845 3844 38879
rect 3792 38836 3844 38845
rect 16672 38836 16724 38888
rect 18512 38836 18564 38888
rect 4988 38700 5040 38752
rect 5172 38743 5224 38752
rect 5172 38709 5181 38743
rect 5181 38709 5215 38743
rect 5215 38709 5224 38743
rect 5172 38700 5224 38709
rect 10324 38743 10376 38752
rect 10324 38709 10333 38743
rect 10333 38709 10367 38743
rect 10367 38709 10376 38743
rect 10324 38700 10376 38709
rect 13544 38743 13596 38752
rect 13544 38709 13553 38743
rect 13553 38709 13587 38743
rect 13587 38709 13596 38743
rect 13544 38700 13596 38709
rect 19524 38700 19576 38752
rect 20536 38700 20588 38752
rect 34704 38879 34756 38888
rect 34704 38845 34713 38879
rect 34713 38845 34747 38879
rect 34747 38845 34756 38879
rect 34704 38836 34756 38845
rect 42432 38879 42484 38888
rect 42432 38845 42441 38879
rect 42441 38845 42475 38879
rect 42475 38845 42484 38879
rect 42432 38836 42484 38845
rect 47492 38836 47544 38888
rect 47952 38879 48004 38888
rect 47952 38845 47961 38879
rect 47961 38845 47995 38879
rect 47995 38845 48004 38879
rect 47952 38836 48004 38845
rect 55312 38879 55364 38888
rect 55312 38845 55321 38879
rect 55321 38845 55355 38879
rect 55355 38845 55364 38879
rect 55312 38836 55364 38845
rect 30840 38700 30892 38752
rect 36636 38700 36688 38752
rect 46756 38743 46808 38752
rect 46756 38709 46765 38743
rect 46765 38709 46799 38743
rect 46799 38709 46808 38743
rect 46756 38700 46808 38709
rect 49792 38743 49844 38752
rect 49792 38709 49801 38743
rect 49801 38709 49835 38743
rect 49835 38709 49844 38743
rect 49792 38700 49844 38709
rect 49884 38700 49936 38752
rect 53748 38700 53800 38752
rect 54852 38743 54904 38752
rect 54852 38709 54861 38743
rect 54861 38709 54895 38743
rect 54895 38709 54904 38743
rect 54852 38700 54904 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 27528 38496 27580 38548
rect 31116 38539 31168 38548
rect 31116 38505 31125 38539
rect 31125 38505 31159 38539
rect 31159 38505 31168 38539
rect 31116 38496 31168 38505
rect 36084 38539 36136 38548
rect 36084 38505 36093 38539
rect 36093 38505 36127 38539
rect 36127 38505 36136 38539
rect 36084 38496 36136 38505
rect 46848 38539 46900 38548
rect 46848 38505 46857 38539
rect 46857 38505 46891 38539
rect 46891 38505 46900 38539
rect 46848 38496 46900 38505
rect 53012 38496 53064 38548
rect 47492 38403 47544 38412
rect 47492 38369 47501 38403
rect 47501 38369 47535 38403
rect 47535 38369 47544 38403
rect 47492 38360 47544 38369
rect 53748 38496 53800 38548
rect 56692 38539 56744 38548
rect 56692 38505 56701 38539
rect 56701 38505 56735 38539
rect 56735 38505 56744 38539
rect 56692 38496 56744 38505
rect 4988 38335 5040 38344
rect 4988 38301 4997 38335
rect 4997 38301 5031 38335
rect 5031 38301 5040 38335
rect 4988 38292 5040 38301
rect 8944 38335 8996 38344
rect 8944 38301 8953 38335
rect 8953 38301 8987 38335
rect 8987 38301 8996 38335
rect 8944 38292 8996 38301
rect 10324 38292 10376 38344
rect 12164 38292 12216 38344
rect 13544 38292 13596 38344
rect 14740 38292 14792 38344
rect 19524 38335 19576 38344
rect 19524 38301 19558 38335
rect 19558 38301 19576 38335
rect 5816 38224 5868 38276
rect 15844 38224 15896 38276
rect 17960 38224 18012 38276
rect 18512 38224 18564 38276
rect 19524 38292 19576 38301
rect 21088 38335 21140 38344
rect 21088 38301 21097 38335
rect 21097 38301 21131 38335
rect 21131 38301 21140 38335
rect 21088 38292 21140 38301
rect 21824 38292 21876 38344
rect 24400 38335 24452 38344
rect 24400 38301 24409 38335
rect 24409 38301 24443 38335
rect 24443 38301 24452 38335
rect 24400 38292 24452 38301
rect 26240 38335 26292 38344
rect 26240 38301 26249 38335
rect 26249 38301 26283 38335
rect 26283 38301 26292 38335
rect 26240 38292 26292 38301
rect 30012 38335 30064 38344
rect 30012 38301 30046 38335
rect 30046 38301 30064 38335
rect 22376 38224 22428 38276
rect 6368 38199 6420 38208
rect 6368 38165 6377 38199
rect 6377 38165 6411 38199
rect 6411 38165 6420 38199
rect 6368 38156 6420 38165
rect 10324 38199 10376 38208
rect 10324 38165 10333 38199
rect 10333 38165 10367 38199
rect 10367 38165 10376 38199
rect 10324 38156 10376 38165
rect 13452 38199 13504 38208
rect 13452 38165 13461 38199
rect 13461 38165 13495 38199
rect 13495 38165 13504 38199
rect 13452 38156 13504 38165
rect 16948 38156 17000 38208
rect 17868 38199 17920 38208
rect 17868 38165 17877 38199
rect 17877 38165 17911 38199
rect 17911 38165 17920 38199
rect 17868 38156 17920 38165
rect 20628 38199 20680 38208
rect 20628 38165 20637 38199
rect 20637 38165 20671 38199
rect 20671 38165 20680 38199
rect 20628 38156 20680 38165
rect 22192 38156 22244 38208
rect 26332 38156 26384 38208
rect 27712 38224 27764 38276
rect 30012 38292 30064 38301
rect 31760 38292 31812 38344
rect 34704 38335 34756 38344
rect 34704 38301 34713 38335
rect 34713 38301 34747 38335
rect 34747 38301 34756 38335
rect 34704 38292 34756 38301
rect 38752 38292 38804 38344
rect 42432 38292 42484 38344
rect 45192 38292 45244 38344
rect 30196 38224 30248 38276
rect 33508 38224 33560 38276
rect 35348 38224 35400 38276
rect 37556 38224 37608 38276
rect 44456 38224 44508 38276
rect 46756 38292 46808 38344
rect 51540 38335 51592 38344
rect 51540 38301 51549 38335
rect 51549 38301 51583 38335
rect 51583 38301 51592 38335
rect 51540 38292 51592 38301
rect 54852 38292 54904 38344
rect 55312 38335 55364 38344
rect 55312 38301 55321 38335
rect 55321 38301 55355 38335
rect 55355 38301 55364 38335
rect 55312 38292 55364 38301
rect 47492 38224 47544 38276
rect 51448 38224 51500 38276
rect 53748 38224 53800 38276
rect 56692 38224 56744 38276
rect 27804 38156 27856 38208
rect 34796 38156 34848 38208
rect 37924 38199 37976 38208
rect 37924 38165 37933 38199
rect 37933 38165 37967 38199
rect 37967 38165 37976 38199
rect 37924 38156 37976 38165
rect 44272 38199 44324 38208
rect 44272 38165 44281 38199
rect 44281 38165 44315 38199
rect 44315 38165 44324 38199
rect 44272 38156 44324 38165
rect 47032 38156 47084 38208
rect 53840 38156 53892 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 4068 37952 4120 38004
rect 5724 37952 5776 38004
rect 15844 37995 15896 38004
rect 15844 37961 15853 37995
rect 15853 37961 15887 37995
rect 15887 37961 15896 37995
rect 15844 37952 15896 37961
rect 18052 37995 18104 38004
rect 18052 37961 18061 37995
rect 18061 37961 18095 37995
rect 18095 37961 18104 37995
rect 18052 37952 18104 37961
rect 28540 37995 28592 38004
rect 28540 37961 28549 37995
rect 28549 37961 28583 37995
rect 28583 37961 28592 37995
rect 28540 37952 28592 37961
rect 30288 37952 30340 38004
rect 33508 37995 33560 38004
rect 33508 37961 33517 37995
rect 33517 37961 33551 37995
rect 33551 37961 33560 37995
rect 33508 37952 33560 37961
rect 35348 37995 35400 38004
rect 35348 37961 35357 37995
rect 35357 37961 35391 37995
rect 35391 37961 35400 37995
rect 35348 37952 35400 37961
rect 44456 37995 44508 38004
rect 44456 37961 44465 37995
rect 44465 37961 44499 37995
rect 44499 37961 44508 37995
rect 44456 37952 44508 37961
rect 6368 37884 6420 37936
rect 10324 37884 10376 37936
rect 13452 37884 13504 37936
rect 5172 37816 5224 37868
rect 15292 37816 15344 37868
rect 6644 37748 6696 37800
rect 11520 37748 11572 37800
rect 17868 37884 17920 37936
rect 20628 37884 20680 37936
rect 18512 37859 18564 37868
rect 18512 37825 18521 37859
rect 18521 37825 18555 37859
rect 18555 37825 18564 37859
rect 18512 37816 18564 37825
rect 21824 37859 21876 37868
rect 21824 37825 21833 37859
rect 21833 37825 21867 37859
rect 21867 37825 21876 37859
rect 21824 37816 21876 37825
rect 23204 37816 23256 37868
rect 24400 37884 24452 37936
rect 27620 37884 27672 37936
rect 24952 37816 25004 37868
rect 30932 37816 30984 37868
rect 16672 37791 16724 37800
rect 16672 37757 16681 37791
rect 16681 37757 16715 37791
rect 16715 37757 16724 37791
rect 16672 37748 16724 37757
rect 26240 37748 26292 37800
rect 29092 37791 29144 37800
rect 29092 37757 29101 37791
rect 29101 37757 29135 37791
rect 29135 37757 29144 37791
rect 29092 37748 29144 37757
rect 31760 37748 31812 37800
rect 33140 37816 33192 37868
rect 34704 37884 34756 37936
rect 35348 37816 35400 37868
rect 38752 37884 38804 37936
rect 38660 37816 38712 37868
rect 39120 37859 39172 37868
rect 39120 37825 39129 37859
rect 39129 37825 39163 37859
rect 39163 37825 39172 37859
rect 39120 37816 39172 37825
rect 39396 37859 39448 37868
rect 39396 37825 39430 37859
rect 39430 37825 39448 37859
rect 39396 37816 39448 37825
rect 44456 37816 44508 37868
rect 49884 37884 49936 37936
rect 52276 37884 52328 37936
rect 54668 37884 54720 37936
rect 47124 37816 47176 37868
rect 47492 37816 47544 37868
rect 48228 37816 48280 37868
rect 45560 37791 45612 37800
rect 45560 37757 45569 37791
rect 45569 37757 45603 37791
rect 45603 37757 45612 37791
rect 50804 37791 50856 37800
rect 45560 37748 45612 37757
rect 50804 37757 50813 37791
rect 50813 37757 50847 37791
rect 50847 37757 50856 37791
rect 50804 37748 50856 37757
rect 4620 37612 4672 37664
rect 9772 37655 9824 37664
rect 9772 37621 9781 37655
rect 9781 37621 9815 37655
rect 9815 37621 9824 37655
rect 9772 37612 9824 37621
rect 13176 37655 13228 37664
rect 13176 37621 13185 37655
rect 13185 37621 13219 37655
rect 13219 37621 13228 37655
rect 13176 37612 13228 37621
rect 19892 37655 19944 37664
rect 19892 37621 19901 37655
rect 19901 37621 19935 37655
rect 19935 37621 19944 37655
rect 19892 37612 19944 37621
rect 22100 37612 22152 37664
rect 25044 37655 25096 37664
rect 25044 37621 25053 37655
rect 25053 37621 25087 37655
rect 25087 37621 25096 37655
rect 25044 37612 25096 37621
rect 38752 37612 38804 37664
rect 40500 37655 40552 37664
rect 40500 37621 40509 37655
rect 40509 37621 40543 37655
rect 40543 37621 40552 37655
rect 40500 37612 40552 37621
rect 46940 37655 46992 37664
rect 46940 37621 46949 37655
rect 46949 37621 46983 37655
rect 46983 37621 46992 37655
rect 46940 37612 46992 37621
rect 49884 37612 49936 37664
rect 52184 37655 52236 37664
rect 52184 37621 52193 37655
rect 52193 37621 52227 37655
rect 52227 37621 52236 37655
rect 52184 37612 52236 37621
rect 55312 37612 55364 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 17960 37408 18012 37460
rect 22376 37408 22428 37460
rect 27712 37408 27764 37460
rect 30932 37451 30984 37460
rect 30932 37417 30941 37451
rect 30941 37417 30975 37451
rect 30975 37417 30984 37451
rect 30932 37408 30984 37417
rect 33140 37451 33192 37460
rect 33140 37417 33149 37451
rect 33149 37417 33183 37451
rect 33183 37417 33192 37451
rect 33140 37408 33192 37417
rect 37556 37408 37608 37460
rect 42432 37408 42484 37460
rect 8944 37315 8996 37324
rect 8944 37281 8953 37315
rect 8953 37281 8987 37315
rect 8987 37281 8996 37315
rect 8944 37272 8996 37281
rect 14740 37272 14792 37324
rect 34704 37315 34756 37324
rect 34704 37281 34713 37315
rect 34713 37281 34747 37315
rect 34747 37281 34756 37315
rect 34704 37272 34756 37281
rect 48228 37315 48280 37324
rect 48228 37281 48237 37315
rect 48237 37281 48271 37315
rect 48271 37281 48280 37315
rect 48228 37272 48280 37281
rect 4988 37204 5040 37256
rect 6828 37204 6880 37256
rect 9772 37204 9824 37256
rect 11520 37247 11572 37256
rect 6736 37136 6788 37188
rect 9680 37136 9732 37188
rect 6552 37111 6604 37120
rect 6552 37077 6561 37111
rect 6561 37077 6595 37111
rect 6595 37077 6604 37111
rect 6552 37068 6604 37077
rect 9036 37068 9088 37120
rect 9128 37068 9180 37120
rect 11520 37213 11529 37247
rect 11529 37213 11563 37247
rect 11563 37213 11572 37247
rect 11520 37204 11572 37213
rect 13176 37204 13228 37256
rect 16672 37247 16724 37256
rect 16672 37213 16681 37247
rect 16681 37213 16715 37247
rect 16715 37213 16724 37247
rect 16672 37204 16724 37213
rect 16948 37247 17000 37256
rect 16948 37213 16982 37247
rect 16982 37213 17000 37247
rect 16948 37204 17000 37213
rect 15292 37136 15344 37188
rect 19892 37204 19944 37256
rect 21088 37247 21140 37256
rect 21088 37213 21097 37247
rect 21097 37213 21131 37247
rect 21131 37213 21140 37247
rect 21088 37204 21140 37213
rect 24400 37247 24452 37256
rect 24400 37213 24409 37247
rect 24409 37213 24443 37247
rect 24443 37213 24452 37247
rect 24400 37204 24452 37213
rect 25044 37204 25096 37256
rect 20260 37136 20312 37188
rect 26332 37204 26384 37256
rect 29552 37247 29604 37256
rect 29552 37213 29561 37247
rect 29561 37213 29595 37247
rect 29595 37213 29604 37247
rect 29552 37204 29604 37213
rect 29644 37204 29696 37256
rect 31760 37247 31812 37256
rect 31760 37213 31769 37247
rect 31769 37213 31803 37247
rect 31803 37213 31812 37247
rect 31760 37204 31812 37213
rect 34796 37204 34848 37256
rect 35440 37204 35492 37256
rect 36636 37204 36688 37256
rect 40408 37204 40460 37256
rect 45560 37204 45612 37256
rect 47032 37204 47084 37256
rect 55312 37408 55364 37460
rect 56692 37451 56744 37460
rect 56692 37417 56701 37451
rect 56701 37417 56735 37451
rect 56735 37417 56744 37451
rect 56692 37408 56744 37417
rect 55312 37247 55364 37256
rect 55312 37213 55321 37247
rect 55321 37213 55355 37247
rect 55355 37213 55364 37247
rect 55312 37204 55364 37213
rect 33508 37136 33560 37188
rect 50160 37136 50212 37188
rect 53840 37136 53892 37188
rect 56416 37136 56468 37188
rect 10324 37111 10376 37120
rect 10324 37077 10333 37111
rect 10333 37077 10367 37111
rect 10367 37077 10376 37111
rect 10324 37068 10376 37077
rect 12900 37111 12952 37120
rect 12900 37077 12909 37111
rect 12909 37077 12943 37111
rect 12943 37077 12952 37111
rect 12900 37068 12952 37077
rect 15660 37068 15712 37120
rect 20628 37111 20680 37120
rect 20628 37077 20637 37111
rect 20637 37077 20671 37111
rect 20671 37077 20680 37111
rect 20628 37068 20680 37077
rect 25780 37111 25832 37120
rect 25780 37077 25789 37111
rect 25789 37077 25823 37111
rect 25823 37077 25832 37111
rect 25780 37068 25832 37077
rect 26240 37068 26292 37120
rect 35348 37068 35400 37120
rect 47768 37111 47820 37120
rect 47768 37077 47777 37111
rect 47777 37077 47811 37111
rect 47811 37077 47820 37111
rect 47768 37068 47820 37077
rect 50068 37068 50120 37120
rect 52828 37068 52880 37120
rect 53564 37068 53616 37120
rect 53748 37068 53800 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 5816 36907 5868 36916
rect 5816 36873 5825 36907
rect 5825 36873 5859 36907
rect 5859 36873 5868 36907
rect 5816 36864 5868 36873
rect 9680 36864 9732 36916
rect 14740 36864 14792 36916
rect 19432 36864 19484 36916
rect 20260 36907 20312 36916
rect 20260 36873 20269 36907
rect 20269 36873 20303 36907
rect 20303 36873 20312 36907
rect 20260 36864 20312 36873
rect 23204 36907 23256 36916
rect 23204 36873 23213 36907
rect 23213 36873 23247 36907
rect 23247 36873 23256 36907
rect 23204 36864 23256 36873
rect 24952 36864 25004 36916
rect 33508 36907 33560 36916
rect 33508 36873 33517 36907
rect 33517 36873 33551 36907
rect 33551 36873 33560 36907
rect 33508 36864 33560 36873
rect 38660 36907 38712 36916
rect 38660 36873 38669 36907
rect 38669 36873 38703 36907
rect 38703 36873 38712 36907
rect 38660 36864 38712 36873
rect 50160 36864 50212 36916
rect 56416 36907 56468 36916
rect 56416 36873 56425 36907
rect 56425 36873 56459 36907
rect 56459 36873 56468 36907
rect 56416 36864 56468 36873
rect 6552 36796 6604 36848
rect 8484 36796 8536 36848
rect 10324 36796 10376 36848
rect 12900 36796 12952 36848
rect 13360 36796 13412 36848
rect 4528 36728 4580 36780
rect 4988 36728 5040 36780
rect 6644 36728 6696 36780
rect 11520 36771 11572 36780
rect 11520 36737 11529 36771
rect 11529 36737 11563 36771
rect 11563 36737 11572 36771
rect 11520 36728 11572 36737
rect 16672 36771 16724 36780
rect 16672 36737 16681 36771
rect 16681 36737 16715 36771
rect 16715 36737 16724 36771
rect 16672 36728 16724 36737
rect 18052 36728 18104 36780
rect 20628 36796 20680 36848
rect 27344 36839 27396 36848
rect 27344 36805 27353 36839
rect 27353 36805 27387 36839
rect 27387 36805 27396 36839
rect 27344 36796 27396 36805
rect 21088 36728 21140 36780
rect 22468 36728 22520 36780
rect 25044 36728 25096 36780
rect 29092 36728 29144 36780
rect 30932 36728 30984 36780
rect 33508 36728 33560 36780
rect 35440 36728 35492 36780
rect 37924 36796 37976 36848
rect 47768 36796 47820 36848
rect 49884 36796 49936 36848
rect 52184 36796 52236 36848
rect 8392 36703 8444 36712
rect 8392 36669 8401 36703
rect 8401 36669 8435 36703
rect 8435 36669 8444 36703
rect 8392 36660 8444 36669
rect 23664 36703 23716 36712
rect 23664 36669 23673 36703
rect 23673 36669 23707 36703
rect 23707 36669 23716 36703
rect 23664 36660 23716 36669
rect 31760 36660 31812 36712
rect 38660 36728 38712 36780
rect 42432 36728 42484 36780
rect 46940 36728 46992 36780
rect 50160 36728 50212 36780
rect 50804 36771 50856 36780
rect 50804 36737 50813 36771
rect 50813 36737 50847 36771
rect 50847 36737 50856 36771
rect 50804 36728 50856 36737
rect 55220 36796 55272 36848
rect 56692 36728 56744 36780
rect 38844 36660 38896 36712
rect 39120 36703 39172 36712
rect 39120 36669 39129 36703
rect 39129 36669 39163 36703
rect 39163 36669 39172 36703
rect 39120 36660 39172 36669
rect 45560 36660 45612 36712
rect 48228 36660 48280 36712
rect 52092 36592 52144 36644
rect 7932 36567 7984 36576
rect 7932 36533 7941 36567
rect 7941 36533 7975 36567
rect 7975 36533 7984 36567
rect 7932 36524 7984 36533
rect 12900 36567 12952 36576
rect 12900 36533 12909 36567
rect 12909 36533 12943 36567
rect 12943 36533 12952 36567
rect 12900 36524 12952 36533
rect 28908 36524 28960 36576
rect 29828 36524 29880 36576
rect 36728 36567 36780 36576
rect 36728 36533 36737 36567
rect 36737 36533 36771 36567
rect 36771 36533 36780 36567
rect 36728 36524 36780 36533
rect 39488 36524 39540 36576
rect 45652 36524 45704 36576
rect 47032 36567 47084 36576
rect 47032 36533 47041 36567
rect 47041 36533 47075 36567
rect 47075 36533 47084 36567
rect 47032 36524 47084 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 8484 36320 8536 36372
rect 18052 36363 18104 36372
rect 18052 36329 18061 36363
rect 18061 36329 18095 36363
rect 18095 36329 18104 36363
rect 18052 36320 18104 36329
rect 22468 36363 22520 36372
rect 22468 36329 22477 36363
rect 22477 36329 22511 36363
rect 22511 36329 22520 36363
rect 22468 36320 22520 36329
rect 27804 36320 27856 36372
rect 30932 36363 30984 36372
rect 30932 36329 30941 36363
rect 30941 36329 30975 36363
rect 30975 36329 30984 36363
rect 30932 36320 30984 36329
rect 31760 36320 31812 36372
rect 38660 36363 38712 36372
rect 38660 36329 38669 36363
rect 38669 36329 38703 36363
rect 38703 36329 38712 36363
rect 38660 36320 38712 36329
rect 51448 36320 51500 36372
rect 56692 36363 56744 36372
rect 56692 36329 56701 36363
rect 56701 36329 56735 36363
rect 56735 36329 56744 36363
rect 56692 36320 56744 36329
rect 8392 36184 8444 36236
rect 8944 36227 8996 36236
rect 8944 36193 8953 36227
rect 8953 36193 8987 36227
rect 8987 36193 8996 36227
rect 8944 36184 8996 36193
rect 11520 36227 11572 36236
rect 11520 36193 11529 36227
rect 11529 36193 11563 36227
rect 11563 36193 11572 36227
rect 11520 36184 11572 36193
rect 16672 36227 16724 36236
rect 16672 36193 16681 36227
rect 16681 36193 16715 36227
rect 16715 36193 16724 36227
rect 16672 36184 16724 36193
rect 21088 36227 21140 36236
rect 21088 36193 21097 36227
rect 21097 36193 21131 36227
rect 21131 36193 21140 36227
rect 21088 36184 21140 36193
rect 29092 36184 29144 36236
rect 6368 36116 6420 36168
rect 6644 36116 6696 36168
rect 7932 36116 7984 36168
rect 9036 36116 9088 36168
rect 12900 36116 12952 36168
rect 14004 36116 14056 36168
rect 14740 36116 14792 36168
rect 17868 36116 17920 36168
rect 22192 36116 22244 36168
rect 24400 36159 24452 36168
rect 24400 36125 24409 36159
rect 24409 36125 24443 36159
rect 24443 36125 24452 36159
rect 24400 36116 24452 36125
rect 25780 36116 25832 36168
rect 26240 36159 26292 36168
rect 26240 36125 26249 36159
rect 26249 36125 26283 36159
rect 26283 36125 26292 36159
rect 26240 36116 26292 36125
rect 27068 36116 27120 36168
rect 13820 36048 13872 36100
rect 17776 36048 17828 36100
rect 20536 36048 20588 36100
rect 7932 36023 7984 36032
rect 7932 35989 7941 36023
rect 7941 35989 7975 36023
rect 7975 35989 7984 36023
rect 7932 35980 7984 35989
rect 12900 36023 12952 36032
rect 12900 35989 12909 36023
rect 12909 35989 12943 36023
rect 12943 35989 12952 36023
rect 12900 35980 12952 35989
rect 15200 35980 15252 36032
rect 20168 35980 20220 36032
rect 39120 36184 39172 36236
rect 46848 36184 46900 36236
rect 48228 36227 48280 36236
rect 48228 36193 48237 36227
rect 48237 36193 48271 36227
rect 48271 36193 48280 36227
rect 48228 36184 48280 36193
rect 34612 36116 34664 36168
rect 35440 36116 35492 36168
rect 38752 36116 38804 36168
rect 39948 36116 40000 36168
rect 40500 36116 40552 36168
rect 31024 36048 31076 36100
rect 32312 36091 32364 36100
rect 32312 36057 32321 36091
rect 32321 36057 32355 36091
rect 32355 36057 32364 36091
rect 32312 36048 32364 36057
rect 36084 36048 36136 36100
rect 42432 36116 42484 36168
rect 50160 36159 50212 36168
rect 50160 36125 50176 36159
rect 50176 36125 50210 36159
rect 50210 36125 50212 36159
rect 50160 36116 50212 36125
rect 52736 36116 52788 36168
rect 55312 36159 55364 36168
rect 55312 36125 55321 36159
rect 55321 36125 55355 36159
rect 55355 36125 55364 36159
rect 55312 36116 55364 36125
rect 29920 35980 29972 36032
rect 35992 35980 36044 36032
rect 37372 35980 37424 36032
rect 49792 36048 49844 36100
rect 50068 36048 50120 36100
rect 51264 36048 51316 36100
rect 56600 36048 56652 36100
rect 41420 35980 41472 36032
rect 52552 35980 52604 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 6736 35776 6788 35828
rect 7932 35708 7984 35760
rect 12900 35708 12952 35760
rect 3976 35683 4028 35692
rect 3976 35649 3985 35683
rect 3985 35649 4019 35683
rect 4019 35649 4028 35683
rect 3976 35640 4028 35649
rect 11520 35683 11572 35692
rect 11520 35649 11529 35683
rect 11529 35649 11563 35683
rect 11563 35649 11572 35683
rect 11520 35640 11572 35649
rect 6368 35615 6420 35624
rect 6368 35581 6377 35615
rect 6377 35581 6411 35615
rect 6411 35581 6420 35615
rect 6368 35572 6420 35581
rect 14004 35708 14056 35760
rect 22100 35751 22152 35760
rect 22100 35717 22134 35751
rect 22134 35717 22152 35751
rect 22100 35708 22152 35717
rect 23664 35776 23716 35828
rect 24400 35776 24452 35828
rect 25044 35819 25096 35828
rect 25044 35785 25053 35819
rect 25053 35785 25087 35819
rect 25087 35785 25096 35819
rect 25044 35776 25096 35785
rect 28908 35776 28960 35828
rect 29552 35776 29604 35828
rect 29920 35776 29972 35828
rect 31760 35776 31812 35828
rect 33508 35819 33560 35828
rect 33508 35785 33517 35819
rect 33517 35785 33551 35819
rect 33551 35785 33560 35819
rect 33508 35776 33560 35785
rect 36084 35819 36136 35828
rect 36084 35785 36093 35819
rect 36093 35785 36127 35819
rect 36127 35785 36136 35819
rect 36084 35776 36136 35785
rect 39396 35819 39448 35828
rect 39396 35785 39405 35819
rect 39405 35785 39439 35819
rect 39439 35785 39448 35819
rect 39396 35776 39448 35785
rect 13452 35640 13504 35692
rect 20720 35640 20772 35692
rect 21088 35640 21140 35692
rect 23664 35683 23716 35692
rect 23664 35649 23673 35683
rect 23673 35649 23707 35683
rect 23707 35649 23716 35683
rect 23664 35640 23716 35649
rect 28356 35640 28408 35692
rect 30196 35640 30248 35692
rect 36728 35708 36780 35760
rect 39488 35708 39540 35760
rect 41420 35708 41472 35760
rect 47032 35708 47084 35760
rect 36360 35640 36412 35692
rect 42524 35640 42576 35692
rect 50804 35640 50856 35692
rect 53932 35640 53984 35692
rect 55312 35708 55364 35760
rect 56784 35640 56836 35692
rect 27068 35615 27120 35624
rect 27068 35581 27077 35615
rect 27077 35581 27111 35615
rect 27111 35581 27120 35615
rect 27068 35572 27120 35581
rect 28908 35615 28960 35624
rect 4988 35436 5040 35488
rect 12900 35479 12952 35488
rect 12900 35445 12909 35479
rect 12909 35445 12943 35479
rect 12943 35445 12952 35479
rect 12900 35436 12952 35445
rect 13636 35436 13688 35488
rect 16672 35436 16724 35488
rect 17868 35436 17920 35488
rect 19248 35436 19300 35488
rect 27068 35436 27120 35488
rect 28908 35581 28917 35615
rect 28917 35581 28951 35615
rect 28951 35581 28960 35615
rect 28908 35572 28960 35581
rect 34612 35572 34664 35624
rect 37740 35572 37792 35624
rect 39856 35572 39908 35624
rect 45560 35572 45612 35624
rect 52736 35615 52788 35624
rect 28448 35479 28500 35488
rect 28448 35445 28457 35479
rect 28457 35445 28491 35479
rect 28491 35445 28500 35479
rect 28448 35436 28500 35445
rect 30288 35479 30340 35488
rect 30288 35445 30297 35479
rect 30297 35445 30331 35479
rect 30331 35445 30340 35479
rect 30288 35436 30340 35445
rect 40684 35436 40736 35488
rect 47032 35479 47084 35488
rect 47032 35445 47041 35479
rect 47041 35445 47075 35479
rect 47075 35445 47084 35479
rect 47032 35436 47084 35445
rect 52736 35581 52745 35615
rect 52745 35581 52779 35615
rect 52779 35581 52788 35615
rect 52736 35572 52788 35581
rect 50160 35436 50212 35488
rect 51172 35436 51224 35488
rect 54116 35479 54168 35488
rect 54116 35445 54125 35479
rect 54125 35445 54159 35479
rect 54159 35445 54168 35479
rect 54116 35436 54168 35445
rect 55956 35479 56008 35488
rect 55956 35445 55965 35479
rect 55965 35445 55999 35479
rect 55999 35445 56008 35479
rect 55956 35436 56008 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 13820 35232 13872 35284
rect 6828 35096 6880 35148
rect 11520 35139 11572 35148
rect 11520 35105 11529 35139
rect 11529 35105 11563 35139
rect 11563 35105 11572 35139
rect 11520 35096 11572 35105
rect 16672 35232 16724 35284
rect 17776 35275 17828 35284
rect 17776 35241 17785 35275
rect 17785 35241 17819 35275
rect 17819 35241 17828 35275
rect 17776 35232 17828 35241
rect 28356 35232 28408 35284
rect 31024 35275 31076 35284
rect 31024 35241 31033 35275
rect 31033 35241 31067 35275
rect 31067 35241 31076 35275
rect 31024 35232 31076 35241
rect 19248 35139 19300 35148
rect 19248 35105 19257 35139
rect 19257 35105 19291 35139
rect 19291 35105 19300 35139
rect 19248 35096 19300 35105
rect 21088 35139 21140 35148
rect 21088 35105 21097 35139
rect 21097 35105 21131 35139
rect 21131 35105 21140 35139
rect 21088 35096 21140 35105
rect 28908 35096 28960 35148
rect 31760 35232 31812 35284
rect 44456 35275 44508 35284
rect 44456 35241 44465 35275
rect 44465 35241 44499 35275
rect 44499 35241 44508 35275
rect 44456 35232 44508 35241
rect 45560 35232 45612 35284
rect 37740 35139 37792 35148
rect 37740 35105 37749 35139
rect 37749 35105 37783 35139
rect 37783 35105 37792 35139
rect 37740 35096 37792 35105
rect 39948 35096 40000 35148
rect 47124 35232 47176 35284
rect 46848 35164 46900 35216
rect 12900 35028 12952 35080
rect 14004 35028 14056 35080
rect 19524 35071 19576 35080
rect 19524 35037 19558 35071
rect 19558 35037 19576 35071
rect 19524 35028 19576 35037
rect 24400 35028 24452 35080
rect 26240 35028 26292 35080
rect 27068 35071 27120 35080
rect 27068 35037 27077 35071
rect 27077 35037 27111 35071
rect 27111 35037 27120 35071
rect 27068 35028 27120 35037
rect 30288 35028 30340 35080
rect 40684 35071 40736 35080
rect 40684 35037 40718 35071
rect 40718 35037 40736 35071
rect 40684 35028 40736 35037
rect 44180 35028 44232 35080
rect 55312 35139 55364 35148
rect 55312 35105 55321 35139
rect 55321 35105 55355 35139
rect 55355 35105 55364 35139
rect 55312 35096 55364 35105
rect 47032 35028 47084 35080
rect 50160 35071 50212 35080
rect 50160 35037 50169 35071
rect 50169 35037 50203 35071
rect 50203 35037 50212 35071
rect 50160 35028 50212 35037
rect 55956 35028 56008 35080
rect 57152 35071 57204 35080
rect 57152 35037 57161 35071
rect 57161 35037 57195 35071
rect 57195 35037 57204 35071
rect 57152 35028 57204 35037
rect 9588 34960 9640 35012
rect 14740 34960 14792 35012
rect 18236 34960 18288 35012
rect 22836 34960 22888 35012
rect 26976 34960 27028 35012
rect 28356 34960 28408 35012
rect 31852 34960 31904 35012
rect 35992 35003 36044 35012
rect 35992 34969 36001 35003
rect 36001 34969 36035 35003
rect 36035 34969 36044 35003
rect 35992 34960 36044 34969
rect 40132 34960 40184 35012
rect 46848 34960 46900 35012
rect 48964 34960 49016 35012
rect 51908 34960 51960 35012
rect 54024 34960 54076 35012
rect 56876 34960 56928 35012
rect 8300 34935 8352 34944
rect 8300 34901 8309 34935
rect 8309 34901 8343 34935
rect 8343 34901 8352 34935
rect 8300 34892 8352 34901
rect 15476 34935 15528 34944
rect 15476 34901 15485 34935
rect 15485 34901 15519 34935
rect 15519 34901 15528 34935
rect 15476 34892 15528 34901
rect 20628 34935 20680 34944
rect 20628 34901 20637 34935
rect 20637 34901 20671 34935
rect 20671 34901 20680 34935
rect 20628 34892 20680 34901
rect 22468 34935 22520 34944
rect 22468 34901 22477 34935
rect 22477 34901 22511 34935
rect 22511 34901 22520 34935
rect 22468 34892 22520 34901
rect 26608 34935 26660 34944
rect 26608 34901 26617 34935
rect 26617 34901 26651 34935
rect 26651 34901 26660 34935
rect 26608 34892 26660 34901
rect 30380 34892 30432 34944
rect 41788 34935 41840 34944
rect 41788 34901 41797 34935
rect 41797 34901 41831 34935
rect 41831 34901 41840 34935
rect 41788 34892 41840 34901
rect 49700 34892 49752 34944
rect 52092 34892 52144 34944
rect 53012 34892 53064 34944
rect 56692 34935 56744 34944
rect 56692 34901 56701 34935
rect 56701 34901 56735 34935
rect 56735 34901 56744 34935
rect 56692 34892 56744 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 11060 34688 11112 34740
rect 13452 34688 13504 34740
rect 14740 34731 14792 34740
rect 14740 34697 14749 34731
rect 14749 34697 14783 34731
rect 14783 34697 14792 34731
rect 14740 34688 14792 34697
rect 18236 34731 18288 34740
rect 18236 34697 18245 34731
rect 18245 34697 18279 34731
rect 18279 34697 18288 34731
rect 18236 34688 18288 34697
rect 24492 34688 24544 34740
rect 24676 34688 24728 34740
rect 28356 34731 28408 34740
rect 28356 34697 28365 34731
rect 28365 34697 28399 34731
rect 28399 34697 28408 34731
rect 28356 34688 28408 34697
rect 30196 34731 30248 34740
rect 30196 34697 30205 34731
rect 30205 34697 30239 34731
rect 30239 34697 30248 34731
rect 30196 34688 30248 34697
rect 36360 34731 36412 34740
rect 36360 34697 36369 34731
rect 36369 34697 36403 34731
rect 36403 34697 36412 34731
rect 36360 34688 36412 34697
rect 38844 34688 38896 34740
rect 39120 34688 39172 34740
rect 45652 34688 45704 34740
rect 46848 34731 46900 34740
rect 3976 34620 4028 34672
rect 11888 34620 11940 34672
rect 13636 34663 13688 34672
rect 13636 34629 13670 34663
rect 13670 34629 13688 34663
rect 13636 34620 13688 34629
rect 20628 34620 20680 34672
rect 8944 34595 8996 34604
rect 8944 34561 8953 34595
rect 8953 34561 8987 34595
rect 8987 34561 8996 34595
rect 8944 34552 8996 34561
rect 10324 34552 10376 34604
rect 15200 34552 15252 34604
rect 16672 34552 16724 34604
rect 18512 34552 18564 34604
rect 23756 34620 23808 34672
rect 28448 34620 28500 34672
rect 23848 34552 23900 34604
rect 25044 34552 25096 34604
rect 28356 34552 28408 34604
rect 29920 34552 29972 34604
rect 31760 34552 31812 34604
rect 32128 34552 32180 34604
rect 34704 34552 34756 34604
rect 10784 34484 10836 34536
rect 13084 34484 13136 34536
rect 19248 34527 19300 34536
rect 19248 34493 19257 34527
rect 19257 34493 19291 34527
rect 19291 34493 19300 34527
rect 19248 34484 19300 34493
rect 23756 34527 23808 34536
rect 23756 34493 23765 34527
rect 23765 34493 23799 34527
rect 23799 34493 23808 34527
rect 23756 34484 23808 34493
rect 26884 34484 26936 34536
rect 34612 34484 34664 34536
rect 36084 34552 36136 34604
rect 37372 34620 37424 34672
rect 37740 34620 37792 34672
rect 41788 34620 41840 34672
rect 44180 34620 44232 34672
rect 46848 34697 46857 34731
rect 46857 34697 46891 34731
rect 46891 34697 46900 34731
rect 46848 34688 46900 34697
rect 48964 34731 49016 34740
rect 48964 34697 48973 34731
rect 48973 34697 49007 34731
rect 49007 34697 49016 34731
rect 48964 34688 49016 34697
rect 49792 34620 49844 34672
rect 46296 34552 46348 34604
rect 48964 34552 49016 34604
rect 53380 34552 53432 34604
rect 54116 34620 54168 34672
rect 6368 34416 6420 34468
rect 6828 34416 6880 34468
rect 20628 34391 20680 34400
rect 20628 34357 20637 34391
rect 20637 34357 20671 34391
rect 20671 34357 20680 34391
rect 20628 34348 20680 34357
rect 34796 34348 34848 34400
rect 37924 34348 37976 34400
rect 44916 34484 44968 34536
rect 45468 34527 45520 34536
rect 45468 34493 45477 34527
rect 45477 34493 45511 34527
rect 45511 34493 45520 34527
rect 45468 34484 45520 34493
rect 47584 34527 47636 34536
rect 47584 34493 47593 34527
rect 47593 34493 47627 34527
rect 47627 34493 47636 34527
rect 47584 34484 47636 34493
rect 52736 34527 52788 34536
rect 52736 34493 52745 34527
rect 52745 34493 52779 34527
rect 52779 34493 52788 34527
rect 52736 34484 52788 34493
rect 54024 34484 54076 34536
rect 39856 34348 39908 34400
rect 45008 34391 45060 34400
rect 45008 34357 45017 34391
rect 45017 34357 45051 34391
rect 45051 34357 45060 34391
rect 45008 34348 45060 34357
rect 50160 34348 50212 34400
rect 55956 34391 56008 34400
rect 55956 34357 55965 34391
rect 55965 34357 55999 34391
rect 55999 34357 56008 34391
rect 55956 34348 56008 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 10324 34187 10376 34196
rect 10324 34153 10333 34187
rect 10333 34153 10367 34187
rect 10367 34153 10376 34187
rect 10324 34144 10376 34153
rect 15292 34144 15344 34196
rect 18512 34187 18564 34196
rect 18512 34153 18521 34187
rect 18521 34153 18555 34187
rect 18555 34153 18564 34187
rect 18512 34144 18564 34153
rect 21088 34144 21140 34196
rect 21824 34144 21876 34196
rect 26976 34144 27028 34196
rect 31852 34144 31904 34196
rect 36084 34187 36136 34196
rect 36084 34153 36093 34187
rect 36093 34153 36127 34187
rect 36127 34153 36136 34187
rect 36084 34144 36136 34153
rect 50804 34144 50856 34196
rect 53380 34187 53432 34196
rect 53380 34153 53389 34187
rect 53389 34153 53423 34187
rect 53423 34153 53432 34187
rect 53380 34144 53432 34153
rect 56600 34144 56652 34196
rect 8944 34051 8996 34060
rect 8944 34017 8953 34051
rect 8953 34017 8987 34051
rect 8987 34017 8996 34051
rect 8944 34008 8996 34017
rect 16672 34008 16724 34060
rect 26240 34051 26292 34060
rect 26240 34017 26249 34051
rect 26249 34017 26283 34051
rect 26283 34017 26292 34051
rect 26240 34008 26292 34017
rect 28908 34008 28960 34060
rect 39856 34051 39908 34060
rect 39856 34017 39865 34051
rect 39865 34017 39899 34051
rect 39899 34017 39908 34051
rect 39856 34008 39908 34017
rect 57152 34051 57204 34060
rect 57152 34017 57161 34051
rect 57161 34017 57195 34051
rect 57195 34017 57204 34051
rect 57152 34008 57204 34017
rect 3792 33940 3844 33992
rect 6368 33940 6420 33992
rect 10784 33983 10836 33992
rect 10784 33949 10793 33983
rect 10793 33949 10827 33983
rect 10827 33949 10836 33983
rect 10784 33940 10836 33949
rect 14004 33940 14056 33992
rect 15476 33940 15528 33992
rect 19248 33983 19300 33992
rect 19248 33949 19257 33983
rect 19257 33949 19291 33983
rect 19291 33949 19300 33983
rect 19248 33940 19300 33949
rect 20628 33940 20680 33992
rect 24400 33983 24452 33992
rect 24400 33949 24409 33983
rect 24409 33949 24443 33983
rect 24443 33949 24452 33983
rect 24400 33940 24452 33949
rect 29828 33983 29880 33992
rect 29828 33949 29862 33983
rect 29862 33949 29880 33983
rect 31668 33983 31720 33992
rect 29828 33940 29880 33949
rect 31668 33949 31677 33983
rect 31677 33949 31711 33983
rect 31711 33949 31720 33983
rect 31668 33940 31720 33949
rect 34612 33940 34664 33992
rect 34796 33940 34848 33992
rect 37924 33983 37976 33992
rect 37924 33949 37933 33983
rect 37933 33949 37967 33983
rect 37967 33949 37976 33983
rect 37924 33940 37976 33949
rect 39120 33940 39172 33992
rect 42616 33940 42668 33992
rect 44916 33940 44968 33992
rect 47584 33940 47636 33992
rect 50160 33983 50212 33992
rect 50160 33949 50169 33983
rect 50169 33949 50203 33983
rect 50203 33949 50212 33983
rect 50160 33940 50212 33949
rect 52092 33940 52144 33992
rect 6000 33872 6052 33924
rect 7748 33872 7800 33924
rect 10324 33872 10376 33924
rect 12072 33872 12124 33924
rect 18420 33872 18472 33924
rect 20720 33872 20772 33924
rect 6276 33847 6328 33856
rect 6276 33813 6285 33847
rect 6285 33813 6319 33847
rect 6319 33813 6328 33847
rect 6276 33804 6328 33813
rect 8116 33847 8168 33856
rect 8116 33813 8125 33847
rect 8125 33813 8159 33847
rect 8159 33813 8168 33847
rect 8116 33804 8168 33813
rect 12532 33804 12584 33856
rect 20628 33847 20680 33856
rect 20628 33813 20637 33847
rect 20637 33813 20671 33847
rect 20671 33813 20680 33847
rect 20628 33804 20680 33813
rect 25688 33872 25740 33924
rect 26332 33872 26384 33924
rect 33508 33872 33560 33924
rect 39672 33872 39724 33924
rect 43812 33872 43864 33924
rect 45560 33872 45612 33924
rect 48872 33872 48924 33924
rect 50804 33872 50856 33924
rect 51080 33872 51132 33924
rect 52736 33872 52788 33924
rect 56692 33940 56744 33992
rect 57152 33872 57204 33924
rect 58440 33872 58492 33924
rect 24860 33804 24912 33856
rect 25780 33847 25832 33856
rect 25780 33813 25789 33847
rect 25789 33813 25823 33847
rect 25823 33813 25832 33847
rect 25780 33804 25832 33813
rect 33048 33847 33100 33856
rect 33048 33813 33057 33847
rect 33057 33813 33091 33847
rect 33091 33813 33100 33847
rect 33048 33804 33100 33813
rect 39304 33847 39356 33856
rect 39304 33813 39313 33847
rect 39313 33813 39347 33847
rect 39347 33813 39356 33847
rect 39304 33804 39356 33813
rect 40592 33804 40644 33856
rect 43904 33847 43956 33856
rect 43904 33813 43913 33847
rect 43913 33813 43947 33847
rect 43947 33813 43956 33847
rect 43904 33804 43956 33813
rect 46388 33847 46440 33856
rect 46388 33813 46397 33847
rect 46397 33813 46431 33847
rect 46431 33813 46440 33847
rect 46388 33804 46440 33813
rect 48228 33847 48280 33856
rect 48228 33813 48237 33847
rect 48237 33813 48271 33847
rect 48271 33813 48280 33847
rect 48228 33804 48280 33813
rect 58532 33847 58584 33856
rect 58532 33813 58541 33847
rect 58541 33813 58575 33847
rect 58575 33813 58584 33847
rect 58532 33804 58584 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 7748 33643 7800 33652
rect 7748 33609 7757 33643
rect 7757 33609 7791 33643
rect 7791 33609 7800 33643
rect 7748 33600 7800 33609
rect 9588 33643 9640 33652
rect 9588 33609 9597 33643
rect 9597 33609 9631 33643
rect 9631 33609 9640 33643
rect 9588 33600 9640 33609
rect 18420 33643 18472 33652
rect 18420 33609 18429 33643
rect 18429 33609 18463 33643
rect 18463 33609 18472 33643
rect 18420 33600 18472 33609
rect 25044 33643 25096 33652
rect 25044 33609 25053 33643
rect 25053 33609 25087 33643
rect 25087 33609 25096 33643
rect 25044 33600 25096 33609
rect 28356 33643 28408 33652
rect 28356 33609 28365 33643
rect 28365 33609 28399 33643
rect 28399 33609 28408 33643
rect 28356 33600 28408 33609
rect 33508 33643 33560 33652
rect 33508 33609 33517 33643
rect 33517 33609 33551 33643
rect 33551 33609 33560 33643
rect 33508 33600 33560 33609
rect 34704 33600 34756 33652
rect 39672 33643 39724 33652
rect 39672 33609 39681 33643
rect 39681 33609 39715 33643
rect 39715 33609 39724 33643
rect 39672 33600 39724 33609
rect 43812 33643 43864 33652
rect 43812 33609 43821 33643
rect 43821 33609 43855 33643
rect 43855 33609 43864 33643
rect 43812 33600 43864 33609
rect 48964 33643 49016 33652
rect 48964 33609 48973 33643
rect 48973 33609 49007 33643
rect 49007 33609 49016 33643
rect 48964 33600 49016 33609
rect 50804 33643 50856 33652
rect 50804 33609 50813 33643
rect 50813 33609 50847 33643
rect 50847 33609 50856 33643
rect 50804 33600 50856 33609
rect 53932 33600 53984 33652
rect 6276 33532 6328 33584
rect 8576 33532 8628 33584
rect 11888 33575 11940 33584
rect 11888 33541 11897 33575
rect 11897 33541 11931 33575
rect 11931 33541 11940 33575
rect 11888 33532 11940 33541
rect 13360 33532 13412 33584
rect 5172 33464 5224 33516
rect 6368 33507 6420 33516
rect 6368 33473 6377 33507
rect 6377 33473 6411 33507
rect 6411 33473 6420 33507
rect 6368 33464 6420 33473
rect 6920 33464 6972 33516
rect 8944 33464 8996 33516
rect 14740 33464 14792 33516
rect 19248 33532 19300 33584
rect 20628 33532 20680 33584
rect 25780 33532 25832 33584
rect 26608 33532 26660 33584
rect 30380 33532 30432 33584
rect 39304 33532 39356 33584
rect 40132 33575 40184 33584
rect 40132 33541 40141 33575
rect 40141 33541 40175 33575
rect 40175 33541 40184 33575
rect 40132 33532 40184 33541
rect 43904 33532 43956 33584
rect 48228 33532 48280 33584
rect 49700 33575 49752 33584
rect 49700 33541 49734 33575
rect 49734 33541 49752 33575
rect 49700 33532 49752 33541
rect 53012 33575 53064 33584
rect 53012 33541 53046 33575
rect 53046 33541 53064 33575
rect 53012 33532 53064 33541
rect 54668 33532 54720 33584
rect 57152 33532 57204 33584
rect 18880 33464 18932 33516
rect 21824 33507 21876 33516
rect 21824 33473 21833 33507
rect 21833 33473 21867 33507
rect 21867 33473 21876 33507
rect 21824 33464 21876 33473
rect 22100 33507 22152 33516
rect 22100 33473 22134 33507
rect 22134 33473 22152 33507
rect 22100 33464 22152 33473
rect 23756 33464 23808 33516
rect 24400 33464 24452 33516
rect 29920 33464 29972 33516
rect 31760 33464 31812 33516
rect 33876 33464 33928 33516
rect 43812 33464 43864 33516
rect 3792 33396 3844 33448
rect 14004 33396 14056 33448
rect 19248 33439 19300 33448
rect 19248 33405 19257 33439
rect 19257 33405 19291 33439
rect 19291 33405 19300 33439
rect 19248 33396 19300 33405
rect 26976 33439 27028 33448
rect 26976 33405 26985 33439
rect 26985 33405 27019 33439
rect 27019 33405 27028 33439
rect 26976 33396 27028 33405
rect 32128 33439 32180 33448
rect 32128 33405 32137 33439
rect 32137 33405 32171 33439
rect 32171 33405 32180 33439
rect 32128 33396 32180 33405
rect 20536 33328 20588 33380
rect 5908 33260 5960 33312
rect 13084 33260 13136 33312
rect 15476 33303 15528 33312
rect 15476 33269 15485 33303
rect 15485 33269 15519 33303
rect 15519 33269 15528 33303
rect 15476 33260 15528 33269
rect 23204 33303 23256 33312
rect 23204 33269 23213 33303
rect 23213 33269 23247 33303
rect 23247 33269 23256 33303
rect 23204 33260 23256 33269
rect 31208 33303 31260 33312
rect 31208 33269 31217 33303
rect 31217 33269 31251 33303
rect 31251 33269 31260 33303
rect 31208 33260 31260 33269
rect 31668 33260 31720 33312
rect 37924 33396 37976 33448
rect 34704 33260 34756 33312
rect 39856 33260 39908 33312
rect 42156 33396 42208 33448
rect 44180 33396 44232 33448
rect 47584 33439 47636 33448
rect 47584 33405 47593 33439
rect 47593 33405 47627 33439
rect 47627 33405 47636 33439
rect 47584 33396 47636 33405
rect 51080 33396 51132 33448
rect 52736 33439 52788 33448
rect 52736 33405 52745 33439
rect 52745 33405 52779 33439
rect 52779 33405 52788 33439
rect 52736 33396 52788 33405
rect 45652 33303 45704 33312
rect 45652 33269 45661 33303
rect 45661 33269 45695 33303
rect 45695 33269 45704 33303
rect 45652 33260 45704 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 5172 33099 5224 33108
rect 5172 33065 5181 33099
rect 5181 33065 5215 33099
rect 5215 33065 5224 33099
rect 5172 33056 5224 33065
rect 6000 33056 6052 33108
rect 10324 33099 10376 33108
rect 10324 33065 10333 33099
rect 10333 33065 10367 33099
rect 10367 33065 10376 33099
rect 10324 33056 10376 33065
rect 12072 33056 12124 33108
rect 22100 33056 22152 33108
rect 22836 33099 22888 33108
rect 22836 33065 22845 33099
rect 22845 33065 22879 33099
rect 22879 33065 22888 33099
rect 22836 33056 22888 33065
rect 26332 33056 26384 33108
rect 37004 33056 37056 33108
rect 46296 33056 46348 33108
rect 51908 33056 51960 33108
rect 56784 33056 56836 33108
rect 58440 33056 58492 33108
rect 8944 32963 8996 32972
rect 8944 32929 8953 32963
rect 8953 32929 8987 32963
rect 8987 32929 8996 32963
rect 8944 32920 8996 32929
rect 14004 32920 14056 32972
rect 16672 32963 16724 32972
rect 16672 32929 16681 32963
rect 16681 32929 16715 32963
rect 16715 32929 16724 32963
rect 16672 32920 16724 32929
rect 29920 32963 29972 32972
rect 29920 32929 29929 32963
rect 29929 32929 29963 32963
rect 29963 32929 29972 32963
rect 29920 32920 29972 32929
rect 39856 32920 39908 32972
rect 42156 32963 42208 32972
rect 42156 32929 42165 32963
rect 42165 32929 42199 32963
rect 42199 32929 42208 32963
rect 42156 32920 42208 32929
rect 52736 32920 52788 32972
rect 57152 32963 57204 32972
rect 3332 32852 3384 32904
rect 3792 32895 3844 32904
rect 3792 32861 3801 32895
rect 3801 32861 3835 32895
rect 3835 32861 3844 32895
rect 3792 32852 3844 32861
rect 4712 32784 4764 32836
rect 5908 32827 5960 32836
rect 5908 32793 5942 32827
rect 5942 32793 5960 32827
rect 5908 32784 5960 32793
rect 10232 32852 10284 32904
rect 11060 32895 11112 32904
rect 11060 32861 11094 32895
rect 11094 32861 11112 32895
rect 11060 32852 11112 32861
rect 19248 32852 19300 32904
rect 6920 32784 6972 32836
rect 9588 32784 9640 32836
rect 16580 32784 16632 32836
rect 17960 32784 18012 32836
rect 20168 32852 20220 32904
rect 23204 32852 23256 32904
rect 24400 32895 24452 32904
rect 24400 32861 24409 32895
rect 24409 32861 24443 32895
rect 24443 32861 24452 32895
rect 24400 32852 24452 32861
rect 24676 32895 24728 32904
rect 24676 32861 24710 32895
rect 24710 32861 24728 32895
rect 24676 32852 24728 32861
rect 26976 32895 27028 32904
rect 26976 32861 26985 32895
rect 26985 32861 27019 32895
rect 27019 32861 27028 32895
rect 26976 32852 27028 32861
rect 27528 32852 27580 32904
rect 31208 32852 31260 32904
rect 21824 32784 21876 32836
rect 23296 32784 23348 32836
rect 25044 32784 25096 32836
rect 28632 32784 28684 32836
rect 33048 32852 33100 32904
rect 35900 32852 35952 32904
rect 40592 32895 40644 32904
rect 40592 32861 40626 32895
rect 40626 32861 40644 32895
rect 40592 32852 40644 32861
rect 32128 32784 32180 32836
rect 34612 32784 34664 32836
rect 38660 32784 38712 32836
rect 41788 32784 41840 32836
rect 45652 32852 45704 32904
rect 47584 32852 47636 32904
rect 50804 32852 50856 32904
rect 50988 32852 51040 32904
rect 51172 32895 51224 32904
rect 51172 32861 51206 32895
rect 51206 32861 51224 32895
rect 51172 32852 51224 32861
rect 57152 32929 57161 32963
rect 57161 32929 57195 32963
rect 57195 32929 57204 32963
rect 57152 32920 57204 32929
rect 55956 32852 56008 32904
rect 16212 32759 16264 32768
rect 16212 32725 16221 32759
rect 16221 32725 16255 32759
rect 16255 32725 16264 32759
rect 16212 32716 16264 32725
rect 18052 32759 18104 32768
rect 18052 32725 18061 32759
rect 18061 32725 18095 32759
rect 18095 32725 18104 32759
rect 18052 32716 18104 32725
rect 28356 32759 28408 32768
rect 28356 32725 28365 32759
rect 28365 32725 28399 32759
rect 28399 32725 28408 32759
rect 28356 32716 28408 32725
rect 31300 32759 31352 32768
rect 31300 32725 31309 32759
rect 31309 32725 31343 32759
rect 31343 32725 31352 32759
rect 31300 32716 31352 32725
rect 33324 32759 33376 32768
rect 33324 32725 33333 32759
rect 33333 32725 33367 32759
rect 33367 32725 33376 32759
rect 33324 32716 33376 32725
rect 36452 32716 36504 32768
rect 41696 32759 41748 32768
rect 41696 32725 41705 32759
rect 41705 32725 41739 32759
rect 41739 32725 41748 32759
rect 41696 32716 41748 32725
rect 43536 32759 43588 32768
rect 43536 32725 43545 32759
rect 43545 32725 43579 32759
rect 43579 32725 43588 32759
rect 43536 32716 43588 32725
rect 46480 32784 46532 32836
rect 57428 32827 57480 32836
rect 57428 32793 57462 32827
rect 57462 32793 57480 32827
rect 57428 32784 57480 32793
rect 45652 32716 45704 32768
rect 48228 32759 48280 32768
rect 48228 32725 48237 32759
rect 48237 32725 48271 32759
rect 48271 32725 48280 32759
rect 48228 32716 48280 32725
rect 52368 32716 52420 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 4712 32555 4764 32564
rect 4712 32521 4721 32555
rect 4721 32521 4755 32555
rect 4755 32521 4764 32555
rect 4712 32512 4764 32521
rect 8576 32512 8628 32564
rect 9588 32555 9640 32564
rect 9588 32521 9597 32555
rect 9597 32521 9631 32555
rect 9631 32521 9640 32555
rect 9588 32512 9640 32521
rect 18880 32512 18932 32564
rect 23848 32512 23900 32564
rect 25688 32512 25740 32564
rect 31760 32512 31812 32564
rect 38660 32555 38712 32564
rect 38660 32521 38669 32555
rect 38669 32521 38703 32555
rect 38703 32521 38712 32555
rect 38660 32512 38712 32521
rect 43812 32555 43864 32564
rect 43812 32521 43821 32555
rect 43821 32521 43855 32555
rect 43855 32521 43864 32555
rect 43812 32512 43864 32521
rect 45560 32512 45612 32564
rect 48872 32512 48924 32564
rect 57428 32512 57480 32564
rect 8116 32444 8168 32496
rect 8300 32444 8352 32496
rect 12532 32487 12584 32496
rect 12532 32453 12566 32487
rect 12566 32453 12584 32487
rect 12532 32444 12584 32453
rect 18052 32444 18104 32496
rect 22468 32444 22520 32496
rect 31300 32444 31352 32496
rect 33324 32444 33376 32496
rect 37924 32444 37976 32496
rect 3332 32419 3384 32428
rect 3332 32385 3341 32419
rect 3341 32385 3375 32419
rect 3375 32385 3384 32419
rect 3332 32376 3384 32385
rect 5172 32376 5224 32428
rect 6920 32376 6972 32428
rect 12072 32308 12124 32360
rect 13084 32376 13136 32428
rect 13820 32376 13872 32428
rect 16672 32419 16724 32428
rect 16672 32385 16681 32419
rect 16681 32385 16715 32419
rect 16715 32385 16724 32419
rect 16672 32376 16724 32385
rect 17316 32376 17368 32428
rect 19248 32376 19300 32428
rect 21824 32376 21876 32428
rect 24492 32376 24544 32428
rect 29092 32376 29144 32428
rect 29920 32376 29972 32428
rect 31668 32376 31720 32428
rect 34704 32376 34756 32428
rect 36360 32376 36412 32428
rect 39304 32376 39356 32428
rect 41696 32444 41748 32496
rect 40408 32376 40460 32428
rect 42156 32376 42208 32428
rect 44180 32444 44232 32496
rect 43628 32376 43680 32428
rect 45008 32444 45060 32496
rect 48228 32444 48280 32496
rect 58532 32444 58584 32496
rect 47584 32419 47636 32428
rect 47584 32385 47593 32419
rect 47593 32385 47627 32419
rect 47627 32385 47636 32419
rect 47584 32376 47636 32385
rect 52276 32376 52328 32428
rect 52736 32376 52788 32428
rect 57888 32376 57940 32428
rect 27528 32308 27580 32360
rect 35900 32308 35952 32360
rect 37280 32351 37332 32360
rect 37280 32317 37289 32351
rect 37289 32317 37323 32351
rect 37323 32317 37332 32351
rect 37280 32308 37332 32317
rect 50804 32351 50856 32360
rect 50804 32317 50813 32351
rect 50813 32317 50847 32351
rect 50847 32317 50856 32351
rect 50804 32308 50856 32317
rect 17960 32240 18012 32292
rect 10508 32172 10560 32224
rect 13912 32172 13964 32224
rect 29276 32215 29328 32224
rect 29276 32181 29285 32215
rect 29285 32181 29319 32215
rect 29319 32181 29328 32215
rect 29276 32172 29328 32181
rect 33508 32215 33560 32224
rect 33508 32181 33517 32215
rect 33517 32181 33551 32215
rect 33551 32181 33560 32215
rect 33508 32172 33560 32181
rect 35992 32215 36044 32224
rect 35992 32181 36001 32215
rect 36001 32181 36035 32215
rect 36035 32181 36044 32215
rect 35992 32172 36044 32181
rect 41236 32215 41288 32224
rect 41236 32181 41245 32215
rect 41245 32181 41279 32215
rect 41279 32181 41288 32215
rect 41236 32172 41288 32181
rect 51080 32172 51132 32224
rect 55496 32215 55548 32224
rect 55496 32181 55505 32215
rect 55505 32181 55539 32215
rect 55539 32181 55548 32215
rect 55496 32172 55548 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2872 31764 2924 31816
rect 4988 31968 5040 32020
rect 5172 32011 5224 32020
rect 5172 31977 5181 32011
rect 5181 31977 5215 32011
rect 5215 31977 5224 32011
rect 5172 31968 5224 31977
rect 16580 31968 16632 32020
rect 27528 32011 27580 32020
rect 27528 31977 27537 32011
rect 27537 31977 27571 32011
rect 27571 31977 27580 32011
rect 27528 31968 27580 31977
rect 33876 31968 33928 32020
rect 39304 32011 39356 32020
rect 39304 31977 39313 32011
rect 39313 31977 39347 32011
rect 39347 31977 39356 32011
rect 39304 31968 39356 31977
rect 41788 32011 41840 32020
rect 41788 31977 41797 32011
rect 41797 31977 41831 32011
rect 41831 31977 41840 32011
rect 41788 31968 41840 31977
rect 43628 32011 43680 32020
rect 43628 31977 43637 32011
rect 43637 31977 43671 32011
rect 43671 31977 43680 32011
rect 43628 31968 43680 31977
rect 46480 31968 46532 32020
rect 10232 31875 10284 31884
rect 10232 31841 10241 31875
rect 10241 31841 10275 31875
rect 10275 31841 10284 31875
rect 10232 31832 10284 31841
rect 31208 31900 31260 31952
rect 10508 31807 10560 31816
rect 4252 31696 4304 31748
rect 10508 31773 10542 31807
rect 10542 31773 10560 31807
rect 10508 31764 10560 31773
rect 11520 31764 11572 31816
rect 12072 31807 12124 31816
rect 12072 31773 12081 31807
rect 12081 31773 12115 31807
rect 12115 31773 12124 31807
rect 12072 31764 12124 31773
rect 13084 31832 13136 31884
rect 19248 31832 19300 31884
rect 35900 31875 35952 31884
rect 35900 31841 35909 31875
rect 35909 31841 35943 31875
rect 35943 31841 35952 31875
rect 35900 31832 35952 31841
rect 37280 31832 37332 31884
rect 37924 31875 37976 31884
rect 37924 31841 37933 31875
rect 37933 31841 37967 31875
rect 37967 31841 37976 31875
rect 37924 31832 37976 31841
rect 40408 31875 40460 31884
rect 40408 31841 40417 31875
rect 40417 31841 40451 31875
rect 40451 31841 40460 31875
rect 40408 31832 40460 31841
rect 42156 31832 42208 31884
rect 44916 31832 44968 31884
rect 50804 31968 50856 32020
rect 56876 31968 56928 32020
rect 57888 32011 57940 32020
rect 57888 31977 57897 32011
rect 57897 31977 57931 32011
rect 57931 31977 57940 32011
rect 57888 31968 57940 31977
rect 50804 31832 50856 31884
rect 52736 31832 52788 31884
rect 15476 31764 15528 31816
rect 16672 31764 16724 31816
rect 21272 31764 21324 31816
rect 22468 31764 22520 31816
rect 23664 31764 23716 31816
rect 24860 31764 24912 31816
rect 15568 31696 15620 31748
rect 31484 31764 31536 31816
rect 32128 31807 32180 31816
rect 32128 31773 32137 31807
rect 32137 31773 32171 31807
rect 32171 31773 32180 31807
rect 32128 31764 32180 31773
rect 33508 31764 33560 31816
rect 36452 31764 36504 31816
rect 39304 31764 39356 31816
rect 41236 31764 41288 31816
rect 43536 31764 43588 31816
rect 46388 31764 46440 31816
rect 50160 31764 50212 31816
rect 52368 31764 52420 31816
rect 55496 31764 55548 31816
rect 58532 31764 58584 31816
rect 57060 31696 57112 31748
rect 13452 31671 13504 31680
rect 13452 31637 13461 31671
rect 13461 31637 13495 31671
rect 13495 31637 13504 31671
rect 13452 31628 13504 31637
rect 15476 31671 15528 31680
rect 15476 31637 15485 31671
rect 15485 31637 15519 31671
rect 15519 31637 15528 31671
rect 15476 31628 15528 31637
rect 20996 31671 21048 31680
rect 20996 31637 21005 31671
rect 21005 31637 21039 31671
rect 21039 31637 21048 31671
rect 20996 31628 21048 31637
rect 23756 31671 23808 31680
rect 23756 31637 23765 31671
rect 23765 31637 23799 31671
rect 23799 31637 23808 31671
rect 23756 31628 23808 31637
rect 37280 31671 37332 31680
rect 37280 31637 37289 31671
rect 37289 31637 37323 31671
rect 37323 31637 37332 31671
rect 37280 31628 37332 31637
rect 49608 31671 49660 31680
rect 49608 31637 49617 31671
rect 49617 31637 49651 31671
rect 49651 31637 49660 31671
rect 49608 31628 49660 31637
rect 52460 31628 52512 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 4252 31467 4304 31476
rect 4252 31433 4261 31467
rect 4261 31433 4295 31467
rect 4295 31433 4304 31467
rect 4252 31424 4304 31433
rect 14740 31467 14792 31476
rect 14740 31433 14749 31467
rect 14749 31433 14783 31467
rect 14783 31433 14792 31467
rect 14740 31424 14792 31433
rect 21272 31467 21324 31476
rect 21272 31433 21281 31467
rect 21281 31433 21315 31467
rect 21315 31433 21324 31467
rect 21272 31424 21324 31433
rect 30840 31424 30892 31476
rect 31116 31467 31168 31476
rect 31116 31433 31125 31467
rect 31125 31433 31159 31467
rect 31159 31433 31168 31467
rect 34612 31467 34664 31476
rect 31116 31424 31168 31433
rect 3700 31356 3752 31408
rect 33600 31356 33652 31408
rect 34612 31433 34621 31467
rect 34621 31433 34655 31467
rect 34655 31433 34664 31467
rect 34612 31424 34664 31433
rect 36360 31424 36412 31476
rect 43996 31467 44048 31476
rect 43996 31433 44005 31467
rect 44005 31433 44039 31467
rect 44039 31433 44048 31467
rect 43996 31424 44048 31433
rect 51264 31424 51316 31476
rect 2872 31331 2924 31340
rect 2872 31297 2881 31331
rect 2881 31297 2915 31331
rect 2915 31297 2924 31331
rect 2872 31288 2924 31297
rect 3976 31288 4028 31340
rect 11520 31331 11572 31340
rect 11520 31297 11529 31331
rect 11529 31297 11563 31331
rect 11563 31297 11572 31331
rect 11520 31288 11572 31297
rect 13452 31288 13504 31340
rect 13912 31288 13964 31340
rect 16672 31288 16724 31340
rect 19340 31288 19392 31340
rect 21272 31288 21324 31340
rect 22468 31288 22520 31340
rect 23296 31288 23348 31340
rect 13084 31220 13136 31272
rect 19248 31220 19300 31272
rect 12900 31127 12952 31136
rect 12900 31093 12909 31127
rect 12909 31093 12943 31127
rect 12943 31093 12952 31127
rect 12900 31084 12952 31093
rect 19432 31127 19484 31136
rect 19432 31093 19441 31127
rect 19441 31093 19475 31127
rect 19475 31093 19484 31127
rect 19432 31084 19484 31093
rect 24584 31127 24636 31136
rect 24584 31093 24593 31127
rect 24593 31093 24627 31127
rect 24627 31093 24636 31127
rect 24584 31084 24636 31093
rect 27068 31288 27120 31340
rect 29736 31288 29788 31340
rect 34704 31288 34756 31340
rect 37280 31356 37332 31408
rect 40500 31356 40552 31408
rect 44272 31356 44324 31408
rect 37924 31288 37976 31340
rect 40592 31288 40644 31340
rect 42432 31288 42484 31340
rect 42616 31331 42668 31340
rect 42616 31297 42625 31331
rect 42625 31297 42659 31331
rect 42659 31297 42668 31331
rect 42616 31288 42668 31297
rect 45652 31331 45704 31340
rect 45652 31297 45661 31331
rect 45661 31297 45695 31331
rect 45695 31297 45704 31331
rect 45652 31288 45704 31297
rect 46940 31288 46992 31340
rect 47584 31288 47636 31340
rect 50804 31331 50856 31340
rect 50804 31297 50813 31331
rect 50813 31297 50847 31331
rect 50847 31297 50856 31331
rect 50804 31288 50856 31297
rect 52184 31288 52236 31340
rect 56692 31288 56744 31340
rect 25044 31263 25096 31272
rect 25044 31229 25053 31263
rect 25053 31229 25087 31263
rect 25087 31229 25096 31263
rect 25044 31220 25096 31229
rect 27528 31220 27580 31272
rect 33232 31263 33284 31272
rect 33232 31229 33241 31263
rect 33241 31229 33275 31263
rect 33275 31229 33284 31263
rect 33232 31220 33284 31229
rect 39580 31220 39632 31272
rect 52736 31220 52788 31272
rect 26240 31084 26292 31136
rect 26424 31127 26476 31136
rect 26424 31093 26433 31127
rect 26433 31093 26467 31127
rect 26467 31093 26476 31127
rect 26424 31084 26476 31093
rect 29368 31127 29420 31136
rect 29368 31093 29377 31127
rect 29377 31093 29411 31127
rect 29411 31093 29420 31127
rect 29368 31084 29420 31093
rect 39672 31127 39724 31136
rect 39672 31093 39681 31127
rect 39681 31093 39715 31127
rect 39715 31093 39724 31127
rect 39672 31084 39724 31093
rect 41696 31084 41748 31136
rect 47032 31127 47084 31136
rect 47032 31093 47041 31127
rect 47041 31093 47075 31127
rect 47075 31093 47084 31127
rect 47032 31084 47084 31093
rect 55588 31127 55640 31136
rect 55588 31093 55597 31127
rect 55597 31093 55631 31127
rect 55631 31093 55640 31127
rect 55588 31084 55640 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 13820 30880 13872 30932
rect 15568 30880 15620 30932
rect 17316 30923 17368 30932
rect 17316 30889 17325 30923
rect 17325 30889 17359 30923
rect 17359 30889 17368 30923
rect 17316 30880 17368 30889
rect 33232 30880 33284 30932
rect 39304 30923 39356 30932
rect 39304 30889 39313 30923
rect 39313 30889 39347 30923
rect 39347 30889 39356 30923
rect 39304 30880 39356 30889
rect 52276 30923 52328 30932
rect 52276 30889 52285 30923
rect 52285 30889 52319 30923
rect 52319 30889 52328 30923
rect 52276 30880 52328 30889
rect 58532 30923 58584 30932
rect 58532 30889 58541 30923
rect 58541 30889 58575 30923
rect 58575 30889 58584 30923
rect 58532 30880 58584 30889
rect 41236 30812 41288 30864
rect 11520 30744 11572 30796
rect 22468 30787 22520 30796
rect 22468 30753 22477 30787
rect 22477 30753 22511 30787
rect 22511 30753 22520 30787
rect 22468 30744 22520 30753
rect 42800 30744 42852 30796
rect 47584 30744 47636 30796
rect 4528 30676 4580 30728
rect 7012 30676 7064 30728
rect 9312 30719 9364 30728
rect 9312 30685 9321 30719
rect 9321 30685 9355 30719
rect 9355 30685 9364 30719
rect 9312 30676 9364 30685
rect 12900 30676 12952 30728
rect 14096 30719 14148 30728
rect 14096 30685 14105 30719
rect 14105 30685 14139 30719
rect 14139 30685 14148 30719
rect 14096 30676 14148 30685
rect 15476 30676 15528 30728
rect 15936 30719 15988 30728
rect 15936 30685 15945 30719
rect 15945 30685 15979 30719
rect 15979 30685 15988 30719
rect 15936 30676 15988 30685
rect 16212 30719 16264 30728
rect 16212 30685 16246 30719
rect 16246 30685 16264 30719
rect 16212 30676 16264 30685
rect 20628 30719 20680 30728
rect 20628 30685 20637 30719
rect 20637 30685 20671 30719
rect 20671 30685 20680 30719
rect 20628 30676 20680 30685
rect 5816 30608 5868 30660
rect 8208 30608 8260 30660
rect 10968 30608 11020 30660
rect 23756 30676 23808 30728
rect 24952 30676 25004 30728
rect 27528 30676 27580 30728
rect 29368 30676 29420 30728
rect 32128 30676 32180 30728
rect 34704 30719 34756 30728
rect 34704 30685 34713 30719
rect 34713 30685 34747 30719
rect 34747 30685 34756 30719
rect 34704 30676 34756 30685
rect 35992 30676 36044 30728
rect 24492 30608 24544 30660
rect 29276 30608 29328 30660
rect 33508 30608 33560 30660
rect 37740 30608 37792 30660
rect 39672 30676 39724 30728
rect 42984 30676 43036 30728
rect 39580 30608 39632 30660
rect 44272 30676 44324 30728
rect 45652 30676 45704 30728
rect 49608 30676 49660 30728
rect 50804 30676 50856 30728
rect 52460 30676 52512 30728
rect 52736 30719 52788 30728
rect 52736 30685 52745 30719
rect 52745 30685 52779 30719
rect 52779 30685 52788 30719
rect 52736 30676 52788 30685
rect 55588 30719 55640 30728
rect 55588 30685 55622 30719
rect 55622 30685 55640 30719
rect 55588 30676 55640 30685
rect 57060 30676 57112 30728
rect 44364 30608 44416 30660
rect 47124 30608 47176 30660
rect 56600 30608 56652 30660
rect 56784 30608 56836 30660
rect 5264 30583 5316 30592
rect 5264 30549 5273 30583
rect 5273 30549 5307 30583
rect 5307 30549 5316 30583
rect 5264 30540 5316 30549
rect 6184 30540 6236 30592
rect 9680 30540 9732 30592
rect 22008 30583 22060 30592
rect 22008 30549 22017 30583
rect 22017 30549 22051 30583
rect 22051 30549 22060 30583
rect 22008 30540 22060 30549
rect 23848 30583 23900 30592
rect 23848 30549 23857 30583
rect 23857 30549 23891 30583
rect 23891 30549 23900 30583
rect 23848 30540 23900 30549
rect 27160 30583 27212 30592
rect 27160 30549 27169 30583
rect 27169 30549 27203 30583
rect 27203 30549 27212 30583
rect 27160 30540 27212 30549
rect 29000 30583 29052 30592
rect 29000 30549 29009 30583
rect 29009 30549 29043 30583
rect 29043 30549 29052 30583
rect 29000 30540 29052 30549
rect 31760 30540 31812 30592
rect 36084 30583 36136 30592
rect 36084 30549 36093 30583
rect 36093 30549 36127 30583
rect 36127 30549 36136 30583
rect 36084 30540 36136 30549
rect 42616 30583 42668 30592
rect 42616 30549 42625 30583
rect 42625 30549 42659 30583
rect 42659 30549 42668 30583
rect 42616 30540 42668 30549
rect 44180 30540 44232 30592
rect 47768 30583 47820 30592
rect 47768 30549 47777 30583
rect 47777 30549 47811 30583
rect 47811 30549 47820 30583
rect 47768 30540 47820 30549
rect 49608 30583 49660 30592
rect 49608 30549 49617 30583
rect 49617 30549 49651 30583
rect 49651 30549 49660 30583
rect 49608 30540 49660 30549
rect 55404 30540 55456 30592
rect 57244 30540 57296 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 3976 30379 4028 30388
rect 3976 30345 3985 30379
rect 3985 30345 4019 30379
rect 4019 30345 4028 30379
rect 3976 30336 4028 30345
rect 5816 30379 5868 30388
rect 5816 30345 5825 30379
rect 5825 30345 5859 30379
rect 5859 30345 5868 30379
rect 5816 30336 5868 30345
rect 10968 30379 11020 30388
rect 10968 30345 10977 30379
rect 10977 30345 11011 30379
rect 11011 30345 11020 30379
rect 10968 30336 11020 30345
rect 19340 30336 19392 30388
rect 21272 30379 21324 30388
rect 21272 30345 21281 30379
rect 21281 30345 21315 30379
rect 21315 30345 21324 30379
rect 21272 30336 21324 30345
rect 24492 30336 24544 30388
rect 29736 30379 29788 30388
rect 29736 30345 29745 30379
rect 29745 30345 29779 30379
rect 29779 30345 29788 30379
rect 29736 30336 29788 30345
rect 33508 30379 33560 30388
rect 33508 30345 33517 30379
rect 33517 30345 33551 30379
rect 33551 30345 33560 30379
rect 33508 30336 33560 30345
rect 40592 30336 40644 30388
rect 52184 30379 52236 30388
rect 52184 30345 52193 30379
rect 52193 30345 52227 30379
rect 52227 30345 52236 30379
rect 52184 30336 52236 30345
rect 56692 30379 56744 30388
rect 56692 30345 56701 30379
rect 56701 30345 56735 30379
rect 56735 30345 56744 30379
rect 56692 30336 56744 30345
rect 3976 30200 4028 30252
rect 4528 30200 4580 30252
rect 5816 30200 5868 30252
rect 8392 30200 8444 30252
rect 15660 30268 15712 30320
rect 26424 30268 26476 30320
rect 31208 30268 31260 30320
rect 41236 30268 41288 30320
rect 42524 30268 42576 30320
rect 42800 30268 42852 30320
rect 47768 30268 47820 30320
rect 51080 30311 51132 30320
rect 51080 30277 51114 30311
rect 51114 30277 51132 30311
rect 51080 30268 51132 30277
rect 10876 30200 10928 30252
rect 11520 30243 11572 30252
rect 11520 30209 11529 30243
rect 11529 30209 11563 30243
rect 11563 30209 11572 30243
rect 11520 30200 11572 30209
rect 13268 30200 13320 30252
rect 14004 30200 14056 30252
rect 19984 30200 20036 30252
rect 21916 30200 21968 30252
rect 25872 30200 25924 30252
rect 28908 30200 28960 30252
rect 31392 30200 31444 30252
rect 31576 30200 31628 30252
rect 37740 30243 37792 30252
rect 6920 30132 6972 30184
rect 9312 30132 9364 30184
rect 9588 30175 9640 30184
rect 9588 30141 9597 30175
rect 9597 30141 9631 30175
rect 9631 30141 9640 30175
rect 9588 30132 9640 30141
rect 15936 30132 15988 30184
rect 18052 30175 18104 30184
rect 18052 30141 18061 30175
rect 18061 30141 18095 30175
rect 18095 30141 18104 30175
rect 18052 30132 18104 30141
rect 23204 30175 23256 30184
rect 15384 30064 15436 30116
rect 9128 30039 9180 30048
rect 9128 30005 9137 30039
rect 9137 30005 9171 30039
rect 9171 30005 9180 30039
rect 9128 29996 9180 30005
rect 12440 29996 12492 30048
rect 18052 29996 18104 30048
rect 19248 29996 19300 30048
rect 23204 30141 23213 30175
rect 23213 30141 23247 30175
rect 23247 30141 23256 30175
rect 23204 30132 23256 30141
rect 24952 30132 25004 30184
rect 32128 30175 32180 30184
rect 32128 30141 32137 30175
rect 32137 30141 32171 30175
rect 32171 30141 32180 30175
rect 32128 30132 32180 30141
rect 26240 30064 26292 30116
rect 31484 30064 31536 30116
rect 34704 29996 34756 30048
rect 37740 30209 37749 30243
rect 37749 30209 37783 30243
rect 37783 30209 37792 30243
rect 37740 30200 37792 30209
rect 38844 30200 38896 30252
rect 47032 30200 47084 30252
rect 52552 30200 52604 30252
rect 53012 30243 53064 30252
rect 53012 30209 53046 30243
rect 53046 30209 53064 30243
rect 53012 30200 53064 30209
rect 56692 30200 56744 30252
rect 39580 30175 39632 30184
rect 39580 30141 39589 30175
rect 39589 30141 39623 30175
rect 39623 30141 39632 30175
rect 39580 30132 39632 30141
rect 42984 30132 43036 30184
rect 45652 30175 45704 30184
rect 45652 30141 45661 30175
rect 45661 30141 45695 30175
rect 45695 30141 45704 30175
rect 45652 30132 45704 30141
rect 46848 30132 46900 30184
rect 50804 30175 50856 30184
rect 38660 29996 38712 30048
rect 45836 29996 45888 30048
rect 47032 30039 47084 30048
rect 47032 30005 47041 30039
rect 47041 30005 47075 30039
rect 47075 30005 47084 30039
rect 47032 29996 47084 30005
rect 50804 30141 50813 30175
rect 50813 30141 50847 30175
rect 50847 30141 50856 30175
rect 50804 30132 50856 30141
rect 52736 30175 52788 30184
rect 52736 30141 52745 30175
rect 52745 30141 52779 30175
rect 52779 30141 52788 30175
rect 52736 30132 52788 30141
rect 50160 30064 50212 30116
rect 54116 30039 54168 30048
rect 54116 30005 54125 30039
rect 54125 30005 54159 30039
rect 54159 30005 54168 30039
rect 54116 29996 54168 30005
rect 57060 29996 57112 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 13268 29835 13320 29844
rect 13268 29801 13277 29835
rect 13277 29801 13311 29835
rect 13311 29801 13320 29835
rect 13268 29792 13320 29801
rect 21916 29792 21968 29844
rect 27068 29792 27120 29844
rect 29092 29792 29144 29844
rect 31392 29835 31444 29844
rect 31392 29801 31401 29835
rect 31401 29801 31435 29835
rect 31435 29801 31444 29835
rect 31392 29792 31444 29801
rect 11520 29656 11572 29708
rect 19248 29656 19300 29708
rect 20628 29699 20680 29708
rect 20628 29665 20637 29699
rect 20637 29665 20671 29699
rect 20671 29665 20680 29699
rect 20628 29656 20680 29665
rect 28816 29656 28868 29708
rect 37740 29792 37792 29844
rect 38844 29835 38896 29844
rect 38844 29801 38853 29835
rect 38853 29801 38887 29835
rect 38887 29801 38896 29835
rect 38844 29792 38896 29801
rect 42432 29792 42484 29844
rect 41236 29699 41288 29708
rect 41236 29665 41245 29699
rect 41245 29665 41279 29699
rect 41279 29665 41288 29699
rect 41236 29656 41288 29665
rect 42984 29656 43036 29708
rect 46848 29792 46900 29844
rect 47124 29835 47176 29844
rect 47124 29801 47133 29835
rect 47133 29801 47167 29835
rect 47167 29801 47176 29835
rect 47124 29792 47176 29801
rect 53012 29792 53064 29844
rect 56692 29835 56744 29844
rect 56692 29801 56701 29835
rect 56701 29801 56735 29835
rect 56735 29801 56744 29835
rect 56692 29792 56744 29801
rect 50804 29656 50856 29708
rect 52736 29656 52788 29708
rect 4436 29520 4488 29572
rect 4620 29520 4672 29572
rect 4988 29520 5040 29572
rect 6184 29588 6236 29640
rect 6920 29520 6972 29572
rect 9128 29588 9180 29640
rect 9588 29588 9640 29640
rect 14648 29631 14700 29640
rect 14648 29597 14657 29631
rect 14657 29597 14691 29631
rect 14691 29597 14700 29631
rect 14648 29588 14700 29597
rect 15936 29588 15988 29640
rect 17040 29631 17092 29640
rect 17040 29597 17049 29631
rect 17049 29597 17083 29631
rect 17083 29597 17092 29631
rect 17040 29588 17092 29597
rect 22008 29588 22060 29640
rect 10968 29520 11020 29572
rect 13544 29520 13596 29572
rect 16120 29520 16172 29572
rect 17316 29563 17368 29572
rect 17316 29529 17350 29563
rect 17350 29529 17368 29563
rect 17316 29520 17368 29529
rect 20628 29520 20680 29572
rect 23848 29588 23900 29640
rect 25044 29588 25096 29640
rect 27528 29588 27580 29640
rect 29000 29588 29052 29640
rect 31760 29588 31812 29640
rect 31944 29588 31996 29640
rect 34704 29631 34756 29640
rect 34704 29597 34713 29631
rect 34713 29597 34747 29631
rect 34747 29597 34756 29631
rect 34704 29588 34756 29597
rect 36084 29588 36136 29640
rect 42616 29588 42668 29640
rect 49608 29588 49660 29640
rect 55404 29588 55456 29640
rect 57060 29588 57112 29640
rect 57244 29588 57296 29640
rect 28356 29520 28408 29572
rect 33784 29520 33836 29572
rect 38752 29520 38804 29572
rect 45100 29520 45152 29572
rect 47952 29520 48004 29572
rect 51816 29520 51868 29572
rect 54576 29520 54628 29572
rect 6552 29495 6604 29504
rect 6552 29461 6561 29495
rect 6561 29461 6595 29495
rect 6595 29461 6604 29495
rect 6552 29452 6604 29461
rect 7104 29452 7156 29504
rect 11428 29495 11480 29504
rect 11428 29461 11437 29495
rect 11437 29461 11471 29495
rect 11471 29461 11480 29495
rect 11428 29452 11480 29461
rect 16028 29495 16080 29504
rect 16028 29461 16037 29495
rect 16037 29461 16071 29495
rect 16071 29461 16080 29495
rect 16028 29452 16080 29461
rect 17960 29452 18012 29504
rect 23848 29495 23900 29504
rect 23848 29461 23857 29495
rect 23857 29461 23891 29495
rect 23891 29461 23900 29495
rect 23848 29452 23900 29461
rect 30472 29452 30524 29504
rect 36084 29495 36136 29504
rect 36084 29461 36093 29495
rect 36093 29461 36127 29495
rect 36127 29461 36136 29495
rect 36084 29452 36136 29461
rect 44456 29495 44508 29504
rect 44456 29461 44465 29495
rect 44465 29461 44499 29495
rect 44499 29461 44508 29495
rect 44456 29452 44508 29461
rect 48320 29452 48372 29504
rect 56508 29452 56560 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 3976 29291 4028 29300
rect 3976 29257 3985 29291
rect 3985 29257 4019 29291
rect 4019 29257 4028 29291
rect 3976 29248 4028 29257
rect 5816 29291 5868 29300
rect 5816 29257 5825 29291
rect 5825 29257 5859 29291
rect 5859 29257 5868 29291
rect 5816 29248 5868 29257
rect 10876 29248 10928 29300
rect 16120 29291 16172 29300
rect 16120 29257 16129 29291
rect 16129 29257 16163 29291
rect 16163 29257 16172 29291
rect 16120 29248 16172 29257
rect 20628 29248 20680 29300
rect 25872 29291 25924 29300
rect 25872 29257 25881 29291
rect 25881 29257 25915 29291
rect 25915 29257 25924 29291
rect 25872 29248 25924 29257
rect 28632 29291 28684 29300
rect 28632 29257 28641 29291
rect 28641 29257 28675 29291
rect 28675 29257 28684 29291
rect 28632 29248 28684 29257
rect 31576 29291 31628 29300
rect 31576 29257 31585 29291
rect 31585 29257 31619 29291
rect 31619 29257 31628 29291
rect 31576 29248 31628 29257
rect 5264 29180 5316 29232
rect 4436 29155 4488 29164
rect 4436 29121 4445 29155
rect 4445 29121 4479 29155
rect 4479 29121 4488 29155
rect 4436 29112 4488 29121
rect 6368 29112 6420 29164
rect 11428 29180 11480 29232
rect 15476 29180 15528 29232
rect 23848 29180 23900 29232
rect 24584 29180 24636 29232
rect 24952 29180 25004 29232
rect 27160 29180 27212 29232
rect 30472 29223 30524 29232
rect 30472 29189 30506 29223
rect 30506 29189 30524 29223
rect 30472 29180 30524 29189
rect 10692 29112 10744 29164
rect 14096 29112 14148 29164
rect 14648 29112 14700 29164
rect 16396 29112 16448 29164
rect 18696 29112 18748 29164
rect 20076 29112 20128 29164
rect 23204 29112 23256 29164
rect 25872 29112 25924 29164
rect 32128 29112 32180 29164
rect 36084 29180 36136 29232
rect 41880 29180 41932 29232
rect 45652 29248 45704 29300
rect 35992 29112 36044 29164
rect 9588 29087 9640 29096
rect 9588 29053 9597 29087
rect 9597 29053 9631 29087
rect 9631 29053 9640 29087
rect 9588 29044 9640 29053
rect 16672 29044 16724 29096
rect 17040 29044 17092 29096
rect 22468 29087 22520 29096
rect 22468 29053 22477 29087
rect 22477 29053 22511 29087
rect 22511 29053 22520 29087
rect 22468 29044 22520 29053
rect 28816 29044 28868 29096
rect 34704 29087 34756 29096
rect 34704 29053 34713 29087
rect 34713 29053 34747 29087
rect 34747 29053 34756 29087
rect 34704 29044 34756 29053
rect 6920 28976 6972 29028
rect 23664 28976 23716 29028
rect 14280 28951 14332 28960
rect 14280 28917 14289 28951
rect 14289 28917 14323 28951
rect 14323 28917 14332 28951
rect 14280 28908 14332 28917
rect 18788 28951 18840 28960
rect 18788 28917 18797 28951
rect 18797 28917 18831 28951
rect 18831 28917 18840 28951
rect 18788 28908 18840 28917
rect 34244 28951 34296 28960
rect 34244 28917 34253 28951
rect 34253 28917 34287 28951
rect 34287 28917 34296 28951
rect 34244 28908 34296 28917
rect 36084 28951 36136 28960
rect 36084 28917 36093 28951
rect 36093 28917 36127 28951
rect 36127 28917 36136 28951
rect 36084 28908 36136 28917
rect 37372 28908 37424 28960
rect 39580 29112 39632 29164
rect 41512 29112 41564 29164
rect 42984 29112 43036 29164
rect 47032 29180 47084 29232
rect 49792 29248 49844 29300
rect 56600 29248 56652 29300
rect 47124 29112 47176 29164
rect 48320 29180 48372 29232
rect 51816 29180 51868 29232
rect 54116 29180 54168 29232
rect 48964 29112 49016 29164
rect 50896 29112 50948 29164
rect 57060 29112 57112 29164
rect 45652 29087 45704 29096
rect 45652 29053 45661 29087
rect 45661 29053 45695 29087
rect 45695 29053 45704 29087
rect 45652 29044 45704 29053
rect 49424 29087 49476 29096
rect 49424 29053 49433 29087
rect 49433 29053 49467 29087
rect 49467 29053 49476 29087
rect 49424 29044 49476 29053
rect 41052 29019 41104 29028
rect 41052 28985 41061 29019
rect 41061 28985 41095 29019
rect 41095 28985 41104 29019
rect 41052 28976 41104 28985
rect 46940 28976 46992 29028
rect 50712 28976 50764 29028
rect 53196 28976 53248 29028
rect 38936 28951 38988 28960
rect 38936 28917 38945 28951
rect 38945 28917 38979 28951
rect 38979 28917 38988 28951
rect 38936 28908 38988 28917
rect 45192 28951 45244 28960
rect 45192 28917 45201 28951
rect 45201 28917 45235 28951
rect 45235 28917 45244 28951
rect 45192 28908 45244 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 6368 28747 6420 28756
rect 6368 28713 6377 28747
rect 6377 28713 6411 28747
rect 6411 28713 6420 28747
rect 6368 28704 6420 28713
rect 8392 28747 8444 28756
rect 8392 28713 8401 28747
rect 8401 28713 8435 28747
rect 8435 28713 8444 28747
rect 8392 28704 8444 28713
rect 11520 28704 11572 28756
rect 18696 28747 18748 28756
rect 18696 28713 18705 28747
rect 18705 28713 18739 28747
rect 18739 28713 18748 28747
rect 18696 28704 18748 28713
rect 19984 28704 20036 28756
rect 33784 28747 33836 28756
rect 33784 28713 33793 28747
rect 33793 28713 33827 28747
rect 33827 28713 33836 28747
rect 33784 28704 33836 28713
rect 38752 28747 38804 28756
rect 38752 28713 38761 28747
rect 38761 28713 38795 28747
rect 38795 28713 38804 28747
rect 38752 28704 38804 28713
rect 41512 28747 41564 28756
rect 41512 28713 41521 28747
rect 41521 28713 41555 28747
rect 41555 28713 41564 28747
rect 41512 28704 41564 28713
rect 44364 28704 44416 28756
rect 48964 28747 49016 28756
rect 48964 28713 48973 28747
rect 48973 28713 49007 28747
rect 49007 28713 49016 28747
rect 48964 28704 49016 28713
rect 54576 28747 54628 28756
rect 54576 28713 54585 28747
rect 54585 28713 54619 28747
rect 54619 28713 54628 28747
rect 54576 28704 54628 28713
rect 4988 28611 5040 28620
rect 4988 28577 4997 28611
rect 4997 28577 5031 28611
rect 5031 28577 5040 28611
rect 4988 28568 5040 28577
rect 37372 28611 37424 28620
rect 37372 28577 37381 28611
rect 37381 28577 37415 28611
rect 37415 28577 37424 28611
rect 37372 28568 37424 28577
rect 39580 28568 39632 28620
rect 39948 28568 40000 28620
rect 42984 28568 43036 28620
rect 52736 28568 52788 28620
rect 53196 28611 53248 28620
rect 53196 28577 53205 28611
rect 53205 28577 53239 28611
rect 53239 28577 53248 28611
rect 53196 28568 53248 28577
rect 6552 28500 6604 28552
rect 8300 28500 8352 28552
rect 10692 28543 10744 28552
rect 10692 28509 10701 28543
rect 10701 28509 10735 28543
rect 10735 28509 10744 28543
rect 10692 28500 10744 28509
rect 12532 28500 12584 28552
rect 16672 28500 16724 28552
rect 18052 28500 18104 28552
rect 19248 28543 19300 28552
rect 19248 28509 19257 28543
rect 19257 28509 19291 28543
rect 19291 28509 19300 28543
rect 19248 28500 19300 28509
rect 20996 28500 21048 28552
rect 22468 28500 22520 28552
rect 25136 28543 25188 28552
rect 25136 28509 25145 28543
rect 25145 28509 25179 28543
rect 25179 28509 25188 28543
rect 25136 28500 25188 28509
rect 27620 28500 27672 28552
rect 29552 28543 29604 28552
rect 29552 28509 29561 28543
rect 29561 28509 29595 28543
rect 29595 28509 29604 28543
rect 29552 28500 29604 28509
rect 9128 28432 9180 28484
rect 16856 28407 16908 28416
rect 16856 28373 16865 28407
rect 16865 28373 16899 28407
rect 16899 28373 16908 28407
rect 16856 28364 16908 28373
rect 18052 28364 18104 28416
rect 23480 28432 23532 28484
rect 27068 28432 27120 28484
rect 28080 28432 28132 28484
rect 20536 28364 20588 28416
rect 23204 28407 23256 28416
rect 23204 28373 23213 28407
rect 23213 28373 23247 28407
rect 23247 28373 23256 28407
rect 23204 28364 23256 28373
rect 34244 28500 34296 28552
rect 34704 28500 34756 28552
rect 36084 28500 36136 28552
rect 38936 28500 38988 28552
rect 44456 28500 44508 28552
rect 33140 28432 33192 28484
rect 40684 28432 40736 28484
rect 45652 28432 45704 28484
rect 45836 28500 45888 28552
rect 48320 28500 48372 28552
rect 50160 28543 50212 28552
rect 50160 28509 50169 28543
rect 50169 28509 50203 28543
rect 50203 28509 50212 28543
rect 50160 28500 50212 28509
rect 50804 28500 50856 28552
rect 57060 28543 57112 28552
rect 57060 28509 57069 28543
rect 57069 28509 57103 28543
rect 57103 28509 57112 28543
rect 57060 28500 57112 28509
rect 49056 28432 49108 28484
rect 51448 28432 51500 28484
rect 54760 28432 54812 28484
rect 56692 28432 56744 28484
rect 28356 28407 28408 28416
rect 28356 28373 28365 28407
rect 28365 28373 28399 28407
rect 28399 28373 28408 28407
rect 28356 28364 28408 28373
rect 31484 28364 31536 28416
rect 36176 28407 36228 28416
rect 36176 28373 36185 28407
rect 36185 28373 36219 28407
rect 36219 28373 36228 28407
rect 36176 28364 36228 28373
rect 47124 28407 47176 28416
rect 47124 28373 47133 28407
rect 47133 28373 47167 28407
rect 47167 28373 47176 28407
rect 47124 28364 47176 28373
rect 50620 28364 50672 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 9128 28203 9180 28212
rect 9128 28169 9137 28203
rect 9137 28169 9171 28203
rect 9171 28169 9180 28203
rect 9128 28160 9180 28169
rect 10968 28203 11020 28212
rect 10968 28169 10977 28203
rect 10977 28169 11011 28203
rect 11011 28169 11020 28203
rect 10968 28160 11020 28169
rect 25872 28203 25924 28212
rect 25872 28169 25881 28203
rect 25881 28169 25915 28203
rect 25915 28169 25924 28203
rect 25872 28160 25924 28169
rect 27068 28160 27120 28212
rect 39948 28203 40000 28212
rect 39948 28169 39957 28203
rect 39957 28169 39991 28203
rect 39991 28169 40000 28203
rect 39948 28160 40000 28169
rect 42984 28160 43036 28212
rect 45652 28160 45704 28212
rect 47032 28203 47084 28212
rect 47032 28169 47041 28203
rect 47041 28169 47075 28203
rect 47075 28169 47084 28203
rect 47032 28160 47084 28169
rect 49056 28203 49108 28212
rect 49056 28169 49065 28203
rect 49065 28169 49099 28203
rect 49099 28169 49108 28203
rect 49056 28160 49108 28169
rect 50896 28203 50948 28212
rect 50896 28169 50905 28203
rect 50905 28169 50939 28203
rect 50939 28169 50948 28203
rect 50896 28160 50948 28169
rect 54760 28203 54812 28212
rect 54760 28169 54769 28203
rect 54769 28169 54803 28203
rect 54803 28169 54812 28203
rect 54760 28160 54812 28169
rect 9680 28092 9732 28144
rect 12440 28092 12492 28144
rect 14280 28092 14332 28144
rect 16856 28092 16908 28144
rect 18788 28092 18840 28144
rect 19432 28092 19484 28144
rect 8300 28024 8352 28076
rect 12256 28024 12308 28076
rect 14096 28024 14148 28076
rect 19248 28067 19300 28076
rect 19248 28033 19257 28067
rect 19257 28033 19291 28067
rect 19291 28033 19300 28067
rect 19248 28024 19300 28033
rect 24492 28024 24544 28076
rect 24768 28024 24820 28076
rect 27620 28092 27672 28144
rect 28172 28024 28224 28076
rect 28356 28092 28408 28144
rect 36176 28092 36228 28144
rect 38660 28135 38712 28144
rect 38660 28101 38669 28135
rect 38669 28101 38703 28135
rect 38703 28101 38712 28135
rect 38660 28092 38712 28101
rect 42064 28092 42116 28144
rect 45192 28092 45244 28144
rect 47124 28092 47176 28144
rect 28816 28067 28868 28076
rect 28816 28033 28825 28067
rect 28825 28033 28859 28067
rect 28859 28033 28868 28067
rect 28816 28024 28868 28033
rect 32680 28024 32732 28076
rect 44364 28024 44416 28076
rect 45652 28067 45704 28076
rect 45652 28033 45661 28067
rect 45661 28033 45695 28067
rect 45695 28033 45704 28067
rect 45652 28024 45704 28033
rect 48320 28092 48372 28144
rect 49424 28092 49476 28144
rect 49792 28135 49844 28144
rect 49792 28101 49826 28135
rect 49826 28101 49844 28135
rect 49792 28092 49844 28101
rect 48964 28024 49016 28076
rect 53196 28024 53248 28076
rect 54760 28024 54812 28076
rect 57060 28092 57112 28144
rect 57244 28024 57296 28076
rect 9588 27999 9640 28008
rect 9588 27965 9597 27999
rect 9597 27965 9631 27999
rect 9631 27965 9640 27999
rect 9588 27956 9640 27965
rect 16672 27956 16724 28008
rect 22468 27956 22520 28008
rect 34704 27956 34756 28008
rect 49424 27956 49476 28008
rect 28080 27888 28132 27940
rect 45100 27888 45152 27940
rect 14096 27863 14148 27872
rect 14096 27829 14105 27863
rect 14105 27829 14139 27863
rect 14139 27829 14148 27863
rect 14096 27820 14148 27829
rect 16120 27863 16172 27872
rect 16120 27829 16129 27863
rect 16129 27829 16163 27863
rect 16163 27829 16172 27863
rect 16120 27820 16172 27829
rect 18420 27863 18472 27872
rect 18420 27829 18429 27863
rect 18429 27829 18463 27863
rect 18463 27829 18472 27863
rect 18420 27820 18472 27829
rect 20628 27863 20680 27872
rect 20628 27829 20637 27863
rect 20637 27829 20671 27863
rect 20671 27829 20680 27863
rect 20628 27820 20680 27829
rect 24124 27863 24176 27872
rect 24124 27829 24133 27863
rect 24133 27829 24167 27863
rect 24167 27829 24176 27863
rect 24124 27820 24176 27829
rect 25872 27820 25924 27872
rect 29552 27820 29604 27872
rect 33508 27863 33560 27872
rect 33508 27829 33517 27863
rect 33517 27829 33551 27863
rect 33551 27829 33560 27863
rect 33508 27820 33560 27829
rect 36176 27863 36228 27872
rect 36176 27829 36185 27863
rect 36185 27829 36219 27863
rect 36219 27829 36228 27863
rect 36176 27820 36228 27829
rect 56600 27820 56652 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 8208 27591 8260 27600
rect 8208 27557 8217 27591
rect 8217 27557 8251 27591
rect 8251 27557 8260 27591
rect 8208 27548 8260 27557
rect 13544 27591 13596 27600
rect 13544 27557 13553 27591
rect 13553 27557 13587 27591
rect 13587 27557 13596 27591
rect 13544 27548 13596 27557
rect 16396 27591 16448 27600
rect 16396 27557 16405 27591
rect 16405 27557 16439 27591
rect 16439 27557 16448 27591
rect 16396 27548 16448 27557
rect 20536 27548 20588 27600
rect 28172 27548 28224 27600
rect 41880 27591 41932 27600
rect 41880 27557 41889 27591
rect 41889 27557 41923 27591
rect 41923 27557 41932 27591
rect 41880 27548 41932 27557
rect 44272 27548 44324 27600
rect 54760 27591 54812 27600
rect 54760 27557 54769 27591
rect 54769 27557 54803 27591
rect 54803 27557 54812 27591
rect 54760 27548 54812 27557
rect 19248 27523 19300 27532
rect 19248 27489 19257 27523
rect 19257 27489 19291 27523
rect 19291 27489 19300 27523
rect 19248 27480 19300 27489
rect 39948 27480 40000 27532
rect 42984 27480 43036 27532
rect 50160 27523 50212 27532
rect 50160 27489 50169 27523
rect 50169 27489 50203 27523
rect 50203 27489 50212 27523
rect 50160 27480 50212 27489
rect 6920 27412 6972 27464
rect 7104 27455 7156 27464
rect 7104 27421 7138 27455
rect 7138 27421 7156 27455
rect 7104 27412 7156 27421
rect 12256 27412 12308 27464
rect 14096 27412 14148 27464
rect 14740 27412 14792 27464
rect 16120 27412 16172 27464
rect 16672 27412 16724 27464
rect 18420 27412 18472 27464
rect 20628 27412 20680 27464
rect 22468 27455 22520 27464
rect 22468 27421 22477 27455
rect 22477 27421 22511 27455
rect 22511 27421 22520 27455
rect 22468 27412 22520 27421
rect 24124 27412 24176 27464
rect 23388 27344 23440 27396
rect 25136 27412 25188 27464
rect 27620 27412 27672 27464
rect 30104 27412 30156 27464
rect 31484 27412 31536 27464
rect 34704 27455 34756 27464
rect 34704 27421 34713 27455
rect 34713 27421 34747 27455
rect 34747 27421 34756 27455
rect 34704 27412 34756 27421
rect 36176 27412 36228 27464
rect 37280 27455 37332 27464
rect 37280 27421 37289 27455
rect 37289 27421 37323 27455
rect 37323 27421 37332 27455
rect 37280 27412 37332 27421
rect 41052 27412 41104 27464
rect 44180 27412 44232 27464
rect 44364 27412 44416 27464
rect 54116 27412 54168 27464
rect 57060 27412 57112 27464
rect 25320 27344 25372 27396
rect 29000 27344 29052 27396
rect 32588 27344 32640 27396
rect 40408 27344 40460 27396
rect 45652 27344 45704 27396
rect 48136 27344 48188 27396
rect 50804 27344 50856 27396
rect 54668 27344 54720 27396
rect 57336 27344 57388 27396
rect 18236 27319 18288 27328
rect 18236 27285 18245 27319
rect 18245 27285 18279 27319
rect 18279 27285 18288 27319
rect 18236 27276 18288 27285
rect 23848 27319 23900 27328
rect 23848 27285 23857 27319
rect 23857 27285 23891 27319
rect 23891 27285 23900 27319
rect 23848 27276 23900 27285
rect 24492 27276 24544 27328
rect 27896 27276 27948 27328
rect 32772 27319 32824 27328
rect 32772 27285 32781 27319
rect 32781 27285 32815 27319
rect 32815 27285 32824 27319
rect 32772 27276 32824 27285
rect 36084 27319 36136 27328
rect 36084 27285 36093 27319
rect 36093 27285 36127 27319
rect 36127 27285 36136 27319
rect 36084 27276 36136 27285
rect 39304 27276 39356 27328
rect 46940 27276 46992 27328
rect 48228 27319 48280 27328
rect 48228 27285 48237 27319
rect 48237 27285 48271 27319
rect 48271 27285 48280 27319
rect 48228 27276 48280 27285
rect 51540 27319 51592 27328
rect 51540 27285 51549 27319
rect 51549 27285 51583 27319
rect 51583 27285 51592 27319
rect 51540 27276 51592 27285
rect 57888 27319 57940 27328
rect 57888 27285 57897 27319
rect 57897 27285 57931 27319
rect 57931 27285 57940 27319
rect 57888 27276 57940 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 18052 27115 18104 27124
rect 18052 27081 18061 27115
rect 18061 27081 18095 27115
rect 18095 27081 18104 27115
rect 18052 27072 18104 27081
rect 23480 27115 23532 27124
rect 23480 27081 23489 27115
rect 23489 27081 23523 27115
rect 23523 27081 23532 27115
rect 23480 27072 23532 27081
rect 25320 27115 25372 27124
rect 25320 27081 25329 27115
rect 25329 27081 25363 27115
rect 25363 27081 25372 27115
rect 25320 27072 25372 27081
rect 45652 27115 45704 27124
rect 45652 27081 45661 27115
rect 45661 27081 45695 27115
rect 45695 27081 45704 27115
rect 45652 27072 45704 27081
rect 48964 27115 49016 27124
rect 48964 27081 48973 27115
rect 48973 27081 49007 27115
rect 49007 27081 49016 27115
rect 48964 27072 49016 27081
rect 50804 27115 50856 27124
rect 50804 27081 50813 27115
rect 50813 27081 50847 27115
rect 50847 27081 50856 27115
rect 50804 27072 50856 27081
rect 54668 27072 54720 27124
rect 57244 27072 57296 27124
rect 6920 26936 6972 26988
rect 8484 26936 8536 26988
rect 12256 27004 12308 27056
rect 12532 27004 12584 27056
rect 18236 27004 18288 27056
rect 23848 27004 23900 27056
rect 24768 27004 24820 27056
rect 33508 27004 33560 27056
rect 36084 27004 36136 27056
rect 37280 27004 37332 27056
rect 11796 26979 11848 26988
rect 11796 26945 11830 26979
rect 11830 26945 11848 26979
rect 11796 26936 11848 26945
rect 13636 26936 13688 26988
rect 17960 26936 18012 26988
rect 19248 26936 19300 26988
rect 16672 26911 16724 26920
rect 16672 26877 16681 26911
rect 16681 26877 16715 26911
rect 16715 26877 16724 26911
rect 16672 26868 16724 26877
rect 9036 26775 9088 26784
rect 9036 26741 9045 26775
rect 9045 26741 9079 26775
rect 9079 26741 9088 26775
rect 9036 26732 9088 26741
rect 9128 26732 9180 26784
rect 15108 26732 15160 26784
rect 23112 26936 23164 26988
rect 25780 26936 25832 26988
rect 27804 26936 27856 26988
rect 30104 26936 30156 26988
rect 33140 26936 33192 26988
rect 34704 26979 34756 26988
rect 34704 26945 34713 26979
rect 34713 26945 34747 26979
rect 34747 26945 34756 26979
rect 34704 26936 34756 26945
rect 35716 26936 35768 26988
rect 38660 26936 38712 26988
rect 39948 27004 40000 27056
rect 46296 27004 46348 27056
rect 48228 27004 48280 27056
rect 50712 27004 50764 27056
rect 57888 27004 57940 27056
rect 41236 26936 41288 26988
rect 42524 26936 42576 26988
rect 44364 26936 44416 26988
rect 46388 26936 46440 26988
rect 49424 26979 49476 26988
rect 49424 26945 49433 26979
rect 49433 26945 49467 26979
rect 49467 26945 49476 26979
rect 49424 26936 49476 26945
rect 53196 26936 53248 26988
rect 54760 26936 54812 26988
rect 57060 26936 57112 26988
rect 23388 26868 23440 26920
rect 46848 26868 46900 26920
rect 35992 26800 36044 26852
rect 21272 26775 21324 26784
rect 21272 26741 21281 26775
rect 21281 26741 21315 26775
rect 21315 26741 21324 26775
rect 21272 26732 21324 26741
rect 30196 26775 30248 26784
rect 30196 26741 30205 26775
rect 30205 26741 30239 26775
rect 30239 26741 30248 26775
rect 30196 26732 30248 26741
rect 32404 26732 32456 26784
rect 39028 26775 39080 26784
rect 39028 26741 39037 26775
rect 39037 26741 39071 26775
rect 39071 26741 39080 26775
rect 39028 26732 39080 26741
rect 41788 26732 41840 26784
rect 44456 26732 44508 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 6920 26528 6972 26580
rect 11796 26528 11848 26580
rect 16856 26528 16908 26580
rect 17316 26571 17368 26580
rect 17316 26537 17325 26571
rect 17325 26537 17359 26571
rect 17359 26537 17368 26571
rect 17316 26528 17368 26537
rect 23112 26571 23164 26580
rect 23112 26537 23121 26571
rect 23121 26537 23155 26571
rect 23155 26537 23164 26571
rect 23112 26528 23164 26537
rect 25780 26571 25832 26580
rect 25780 26537 25789 26571
rect 25789 26537 25823 26571
rect 25823 26537 25832 26571
rect 25780 26528 25832 26537
rect 29000 26571 29052 26580
rect 29000 26537 29009 26571
rect 29009 26537 29043 26571
rect 29043 26537 29052 26571
rect 29000 26528 29052 26537
rect 41236 26571 41288 26580
rect 41236 26537 41245 26571
rect 41245 26537 41279 26571
rect 41279 26537 41288 26571
rect 41236 26528 41288 26537
rect 42524 26528 42576 26580
rect 46388 26571 46440 26580
rect 46388 26537 46397 26571
rect 46397 26537 46431 26571
rect 46431 26537 46440 26571
rect 46388 26528 46440 26537
rect 48136 26528 48188 26580
rect 51448 26528 51500 26580
rect 54760 26571 54812 26580
rect 54760 26537 54769 26571
rect 54769 26537 54803 26571
rect 54803 26537 54812 26571
rect 54760 26528 54812 26537
rect 15476 26503 15528 26512
rect 15476 26469 15485 26503
rect 15485 26469 15519 26503
rect 15519 26469 15528 26503
rect 15476 26460 15528 26469
rect 31208 26460 31260 26512
rect 57060 26460 57112 26512
rect 19248 26392 19300 26444
rect 46848 26435 46900 26444
rect 46848 26401 46857 26435
rect 46857 26401 46891 26435
rect 46891 26401 46900 26435
rect 46848 26392 46900 26401
rect 50160 26435 50212 26444
rect 50160 26401 50169 26435
rect 50169 26401 50203 26435
rect 50203 26401 50212 26435
rect 50160 26392 50212 26401
rect 9128 26324 9180 26376
rect 10324 26367 10376 26376
rect 10324 26333 10333 26367
rect 10333 26333 10367 26367
rect 10367 26333 10376 26367
rect 10324 26324 10376 26333
rect 12072 26324 12124 26376
rect 12256 26324 12308 26376
rect 13636 26324 13688 26376
rect 14096 26367 14148 26376
rect 14096 26333 14105 26367
rect 14105 26333 14139 26367
rect 14139 26333 14148 26367
rect 14096 26324 14148 26333
rect 15108 26324 15160 26376
rect 15936 26367 15988 26376
rect 15936 26333 15945 26367
rect 15945 26333 15979 26367
rect 15979 26333 15988 26367
rect 15936 26324 15988 26333
rect 21272 26324 21324 26376
rect 14188 26256 14240 26308
rect 16028 26256 16080 26308
rect 17868 26256 17920 26308
rect 19984 26256 20036 26308
rect 23204 26324 23256 26376
rect 25136 26324 25188 26376
rect 27620 26367 27672 26376
rect 27620 26333 27629 26367
rect 27629 26333 27663 26367
rect 27663 26333 27672 26367
rect 27620 26324 27672 26333
rect 27896 26367 27948 26376
rect 27896 26333 27930 26367
rect 27930 26333 27948 26367
rect 27896 26324 27948 26333
rect 28908 26324 28960 26376
rect 29552 26367 29604 26376
rect 29552 26333 29561 26367
rect 29561 26333 29595 26367
rect 29595 26333 29604 26367
rect 29552 26324 29604 26333
rect 30196 26324 30248 26376
rect 32772 26324 32824 26376
rect 33968 26324 34020 26376
rect 37280 26324 37332 26376
rect 39856 26367 39908 26376
rect 39856 26333 39865 26367
rect 39865 26333 39899 26367
rect 39899 26333 39908 26367
rect 39856 26324 39908 26333
rect 42064 26367 42116 26376
rect 42064 26333 42073 26367
rect 42073 26333 42107 26367
rect 42107 26333 42116 26367
rect 42064 26324 42116 26333
rect 45008 26367 45060 26376
rect 45008 26333 45017 26367
rect 45017 26333 45051 26367
rect 45051 26333 45060 26367
rect 45008 26324 45060 26333
rect 51540 26324 51592 26376
rect 54116 26324 54168 26376
rect 56508 26367 56560 26376
rect 56508 26333 56517 26367
rect 56517 26333 56551 26367
rect 56551 26333 56560 26367
rect 56508 26324 56560 26333
rect 22468 26256 22520 26308
rect 23388 26256 23440 26308
rect 25504 26256 25556 26308
rect 26976 26256 27028 26308
rect 31300 26256 31352 26308
rect 34520 26256 34572 26308
rect 36176 26256 36228 26308
rect 41144 26256 41196 26308
rect 45928 26256 45980 26308
rect 48136 26256 48188 26308
rect 54760 26256 54812 26308
rect 8024 26231 8076 26240
rect 8024 26197 8033 26231
rect 8033 26197 8067 26231
rect 8067 26197 8076 26231
rect 8024 26188 8076 26197
rect 21272 26231 21324 26240
rect 21272 26197 21281 26231
rect 21281 26197 21315 26231
rect 21315 26197 21324 26231
rect 21272 26188 21324 26197
rect 32772 26231 32824 26240
rect 32772 26197 32781 26231
rect 32781 26197 32815 26231
rect 32815 26197 32824 26231
rect 32772 26188 32824 26197
rect 36084 26231 36136 26240
rect 36084 26197 36093 26231
rect 36093 26197 36127 26231
rect 36127 26197 36136 26231
rect 36084 26188 36136 26197
rect 37924 26231 37976 26240
rect 37924 26197 37933 26231
rect 37933 26197 37967 26231
rect 37967 26197 37976 26231
rect 37924 26188 37976 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 8484 26027 8536 26036
rect 8484 25993 8493 26027
rect 8493 25993 8527 26027
rect 8527 25993 8536 26027
rect 8484 25984 8536 25993
rect 8024 25916 8076 25968
rect 9036 25916 9088 25968
rect 16856 25984 16908 26036
rect 17868 25984 17920 26036
rect 25504 26027 25556 26036
rect 25504 25993 25513 26027
rect 25513 25993 25547 26027
rect 25547 25993 25556 26027
rect 25504 25984 25556 25993
rect 31300 25984 31352 26036
rect 38660 26027 38712 26036
rect 38660 25993 38669 26027
rect 38669 25993 38703 26027
rect 38703 25993 38712 26027
rect 38660 25984 38712 25993
rect 39304 25984 39356 26036
rect 23480 25916 23532 25968
rect 5172 25848 5224 25900
rect 6920 25848 6972 25900
rect 9588 25848 9640 25900
rect 10324 25848 10376 25900
rect 13544 25848 13596 25900
rect 14096 25848 14148 25900
rect 15476 25848 15528 25900
rect 15936 25848 15988 25900
rect 20076 25848 20128 25900
rect 20904 25848 20956 25900
rect 23112 25848 23164 25900
rect 24952 25916 25004 25968
rect 36084 25916 36136 25968
rect 44456 25984 44508 26036
rect 57336 26027 57388 26036
rect 57336 25993 57345 26027
rect 57345 25993 57379 26027
rect 57379 25993 57388 26027
rect 57336 25984 57388 25993
rect 50620 25916 50672 25968
rect 56600 25916 56652 25968
rect 25504 25848 25556 25900
rect 26976 25891 27028 25900
rect 26976 25857 26985 25891
rect 26985 25857 27019 25891
rect 27019 25857 27028 25891
rect 26976 25848 27028 25857
rect 27712 25848 27764 25900
rect 30104 25848 30156 25900
rect 30840 25848 30892 25900
rect 32956 25891 33008 25900
rect 32956 25857 32965 25891
rect 32965 25857 32999 25891
rect 32999 25857 33008 25891
rect 32956 25848 33008 25857
rect 38660 25848 38712 25900
rect 39856 25848 39908 25900
rect 43076 25848 43128 25900
rect 44364 25848 44416 25900
rect 47952 25891 48004 25900
rect 47952 25857 47961 25891
rect 47961 25857 47995 25891
rect 47995 25857 48004 25891
rect 47952 25848 48004 25857
rect 49424 25848 49476 25900
rect 50160 25891 50212 25900
rect 50160 25857 50169 25891
rect 50169 25857 50203 25891
rect 50203 25857 50212 25891
rect 50160 25848 50212 25857
rect 58164 25848 58216 25900
rect 8944 25823 8996 25832
rect 8944 25789 8953 25823
rect 8953 25789 8987 25823
rect 8987 25789 8996 25823
rect 8944 25780 8996 25789
rect 12072 25780 12124 25832
rect 4620 25644 4672 25696
rect 5816 25687 5868 25696
rect 5816 25653 5825 25687
rect 5825 25653 5859 25687
rect 5859 25653 5868 25687
rect 5816 25644 5868 25653
rect 10324 25687 10376 25696
rect 10324 25653 10333 25687
rect 10333 25653 10367 25687
rect 10367 25653 10376 25687
rect 10324 25644 10376 25653
rect 19892 25780 19944 25832
rect 21824 25823 21876 25832
rect 21824 25789 21833 25823
rect 21833 25789 21867 25823
rect 21867 25789 21876 25823
rect 21824 25780 21876 25789
rect 15384 25687 15436 25696
rect 15384 25653 15393 25687
rect 15393 25653 15427 25687
rect 15427 25653 15436 25687
rect 15384 25644 15436 25653
rect 24492 25644 24544 25696
rect 29092 25644 29144 25696
rect 33968 25644 34020 25696
rect 37280 25823 37332 25832
rect 37280 25789 37289 25823
rect 37289 25789 37323 25823
rect 37323 25789 37332 25823
rect 37280 25780 37332 25789
rect 42432 25823 42484 25832
rect 42432 25789 42441 25823
rect 42441 25789 42475 25823
rect 42475 25789 42484 25823
rect 42432 25780 42484 25789
rect 54116 25823 54168 25832
rect 54116 25789 54125 25823
rect 54125 25789 54159 25823
rect 54159 25789 54168 25823
rect 54116 25780 54168 25789
rect 35440 25644 35492 25696
rect 40500 25687 40552 25696
rect 40500 25653 40509 25687
rect 40509 25653 40543 25687
rect 40543 25653 40552 25687
rect 40500 25644 40552 25653
rect 43812 25687 43864 25696
rect 43812 25653 43821 25687
rect 43821 25653 43855 25687
rect 43855 25653 43864 25687
rect 43812 25644 43864 25653
rect 45652 25687 45704 25696
rect 45652 25653 45661 25687
rect 45661 25653 45695 25687
rect 45695 25653 45704 25687
rect 45652 25644 45704 25653
rect 49516 25644 49568 25696
rect 51540 25687 51592 25696
rect 51540 25653 51549 25687
rect 51549 25653 51583 25687
rect 51583 25653 51592 25687
rect 51540 25644 51592 25653
rect 55496 25687 55548 25696
rect 55496 25653 55505 25687
rect 55505 25653 55539 25687
rect 55539 25653 55548 25687
rect 55496 25644 55548 25653
rect 56876 25644 56928 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 13544 25483 13596 25492
rect 13544 25449 13553 25483
rect 13553 25449 13587 25483
rect 13587 25449 13596 25483
rect 13544 25440 13596 25449
rect 14188 25440 14240 25492
rect 23112 25483 23164 25492
rect 23112 25449 23121 25483
rect 23121 25449 23155 25483
rect 23155 25449 23164 25483
rect 23112 25440 23164 25449
rect 30840 25440 30892 25492
rect 32680 25440 32732 25492
rect 43076 25483 43128 25492
rect 43076 25449 43085 25483
rect 43085 25449 43119 25483
rect 43119 25449 43128 25483
rect 43076 25440 43128 25449
rect 45928 25440 45980 25492
rect 48136 25440 48188 25492
rect 54760 25483 54812 25492
rect 54760 25449 54769 25483
rect 54769 25449 54803 25483
rect 54803 25449 54812 25483
rect 54760 25440 54812 25449
rect 4528 25279 4580 25288
rect 4528 25245 4537 25279
rect 4537 25245 4571 25279
rect 4571 25245 4580 25279
rect 4528 25236 4580 25245
rect 6368 25279 6420 25288
rect 6368 25245 6377 25279
rect 6377 25245 6411 25279
rect 6411 25245 6420 25279
rect 6368 25236 6420 25245
rect 4344 25100 4396 25152
rect 6092 25168 6144 25220
rect 10324 25236 10376 25288
rect 14740 25304 14792 25356
rect 19892 25347 19944 25356
rect 12072 25168 12124 25220
rect 13452 25168 13504 25220
rect 19892 25313 19901 25347
rect 19901 25313 19935 25347
rect 19935 25313 19944 25347
rect 19892 25304 19944 25313
rect 29552 25347 29604 25356
rect 29552 25313 29561 25347
rect 29561 25313 29595 25347
rect 29595 25313 29604 25347
rect 29552 25304 29604 25313
rect 35716 25304 35768 25356
rect 45008 25347 45060 25356
rect 45008 25313 45017 25347
rect 45017 25313 45051 25347
rect 45051 25313 45060 25347
rect 45008 25304 45060 25313
rect 56600 25304 56652 25356
rect 57060 25440 57112 25492
rect 58164 25483 58216 25492
rect 58164 25449 58173 25483
rect 58173 25449 58207 25483
rect 58207 25449 58216 25483
rect 58164 25440 58216 25449
rect 15384 25279 15436 25288
rect 15384 25245 15418 25279
rect 15418 25245 15436 25279
rect 15384 25236 15436 25245
rect 16672 25236 16724 25288
rect 17316 25279 17368 25288
rect 17316 25245 17325 25279
rect 17325 25245 17359 25279
rect 17359 25245 17368 25279
rect 17316 25236 17368 25245
rect 21272 25236 21324 25288
rect 21732 25279 21784 25288
rect 21732 25245 21741 25279
rect 21741 25245 21775 25279
rect 21775 25245 21784 25279
rect 21732 25236 21784 25245
rect 24952 25236 25004 25288
rect 30104 25236 30156 25288
rect 31392 25279 31444 25288
rect 31392 25245 31401 25279
rect 31401 25245 31435 25279
rect 31435 25245 31444 25279
rect 31392 25236 31444 25245
rect 32772 25236 32824 25288
rect 19248 25168 19300 25220
rect 23204 25168 23256 25220
rect 25320 25168 25372 25220
rect 10324 25143 10376 25152
rect 10324 25109 10333 25143
rect 10333 25109 10367 25143
rect 10367 25109 10376 25143
rect 10324 25100 10376 25109
rect 18696 25143 18748 25152
rect 18696 25109 18705 25143
rect 18705 25109 18739 25143
rect 18739 25109 18748 25143
rect 18696 25100 18748 25109
rect 21272 25143 21324 25152
rect 21272 25109 21281 25143
rect 21281 25109 21315 25143
rect 21315 25109 21324 25143
rect 21272 25100 21324 25109
rect 30196 25168 30248 25220
rect 35440 25168 35492 25220
rect 37924 25236 37976 25288
rect 39856 25279 39908 25288
rect 39856 25245 39865 25279
rect 39865 25245 39899 25279
rect 39899 25245 39908 25279
rect 39856 25236 39908 25245
rect 40500 25236 40552 25288
rect 37280 25168 37332 25220
rect 41788 25236 41840 25288
rect 45652 25236 45704 25288
rect 46848 25279 46900 25288
rect 46848 25245 46857 25279
rect 46857 25245 46891 25279
rect 46891 25245 46900 25279
rect 46848 25236 46900 25245
rect 46940 25236 46992 25288
rect 49516 25236 49568 25288
rect 51540 25236 51592 25288
rect 54116 25236 54168 25288
rect 42432 25168 42484 25220
rect 44364 25168 44416 25220
rect 44916 25168 44968 25220
rect 54760 25168 54812 25220
rect 57336 25168 57388 25220
rect 27620 25143 27672 25152
rect 27620 25109 27629 25143
rect 27629 25109 27663 25143
rect 27663 25109 27672 25143
rect 27620 25100 27672 25109
rect 36084 25143 36136 25152
rect 36084 25109 36093 25143
rect 36093 25109 36127 25143
rect 36127 25109 36136 25143
rect 36084 25100 36136 25109
rect 37924 25143 37976 25152
rect 37924 25109 37933 25143
rect 37933 25109 37967 25143
rect 37967 25109 37976 25143
rect 37924 25100 37976 25109
rect 41236 25143 41288 25152
rect 41236 25109 41245 25143
rect 41245 25109 41279 25143
rect 41279 25109 41288 25143
rect 41236 25100 41288 25109
rect 51540 25143 51592 25152
rect 51540 25109 51549 25143
rect 51549 25109 51583 25143
rect 51583 25109 51592 25143
rect 51540 25100 51592 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 5172 24939 5224 24948
rect 5172 24905 5181 24939
rect 5181 24905 5215 24939
rect 5215 24905 5224 24939
rect 5172 24896 5224 24905
rect 13452 24896 13504 24948
rect 23204 24939 23256 24948
rect 23204 24905 23213 24939
rect 23213 24905 23247 24939
rect 23247 24905 23256 24939
rect 23204 24896 23256 24905
rect 25504 24939 25556 24948
rect 25504 24905 25513 24939
rect 25513 24905 25547 24939
rect 25547 24905 25556 24939
rect 25504 24896 25556 24905
rect 30196 24939 30248 24948
rect 30196 24905 30205 24939
rect 30205 24905 30239 24939
rect 30239 24905 30248 24939
rect 30196 24896 30248 24905
rect 38660 24939 38712 24948
rect 38660 24905 38669 24939
rect 38669 24905 38703 24939
rect 38703 24905 38712 24939
rect 38660 24896 38712 24905
rect 57336 24939 57388 24948
rect 57336 24905 57345 24939
rect 57345 24905 57379 24939
rect 57379 24905 57388 24939
rect 57336 24896 57388 24905
rect 1860 24692 1912 24744
rect 3332 24599 3384 24608
rect 3332 24565 3341 24599
rect 3341 24565 3375 24599
rect 3375 24565 3384 24599
rect 3332 24556 3384 24565
rect 4528 24828 4580 24880
rect 8944 24828 8996 24880
rect 4344 24760 4396 24812
rect 6368 24803 6420 24812
rect 6368 24769 6377 24803
rect 6377 24769 6411 24803
rect 6411 24769 6420 24803
rect 6368 24760 6420 24769
rect 8024 24760 8076 24812
rect 19984 24828 20036 24880
rect 37924 24828 37976 24880
rect 10324 24760 10376 24812
rect 12072 24760 12124 24812
rect 13452 24760 13504 24812
rect 14740 24803 14792 24812
rect 14740 24769 14749 24803
rect 14749 24769 14783 24803
rect 14783 24769 14792 24803
rect 14740 24760 14792 24769
rect 5816 24556 5868 24608
rect 6184 24556 6236 24608
rect 10416 24599 10468 24608
rect 10416 24565 10425 24599
rect 10425 24565 10459 24599
rect 10459 24565 10468 24599
rect 10416 24556 10468 24565
rect 16120 24599 16172 24608
rect 16120 24565 16129 24599
rect 16129 24565 16163 24599
rect 16163 24565 16172 24599
rect 16120 24556 16172 24565
rect 18696 24760 18748 24812
rect 21272 24760 21324 24812
rect 21732 24760 21784 24812
rect 23204 24760 23256 24812
rect 25504 24760 25556 24812
rect 28356 24760 28408 24812
rect 28908 24760 28960 24812
rect 30932 24760 30984 24812
rect 31392 24760 31444 24812
rect 32404 24803 32456 24812
rect 32404 24769 32438 24803
rect 32438 24769 32456 24803
rect 32404 24760 32456 24769
rect 17316 24735 17368 24744
rect 17316 24701 17325 24735
rect 17325 24701 17359 24735
rect 17359 24701 17368 24735
rect 17316 24692 17368 24701
rect 24124 24735 24176 24744
rect 24124 24701 24133 24735
rect 24133 24701 24167 24735
rect 24167 24701 24176 24735
rect 24124 24692 24176 24701
rect 26240 24692 26292 24744
rect 37280 24803 37332 24812
rect 37280 24769 37289 24803
rect 37289 24769 37323 24803
rect 37323 24769 37332 24803
rect 37280 24760 37332 24769
rect 37832 24760 37884 24812
rect 38016 24760 38068 24812
rect 43076 24760 43128 24812
rect 33968 24735 34020 24744
rect 33968 24701 33977 24735
rect 33977 24701 34011 24735
rect 34011 24701 34020 24735
rect 33968 24692 34020 24701
rect 18512 24556 18564 24608
rect 18696 24599 18748 24608
rect 18696 24565 18705 24599
rect 18705 24565 18739 24599
rect 18739 24565 18748 24599
rect 18696 24556 18748 24565
rect 21180 24599 21232 24608
rect 21180 24565 21189 24599
rect 21189 24565 21223 24599
rect 21223 24565 21232 24599
rect 21180 24556 21232 24565
rect 27896 24556 27948 24608
rect 32404 24556 32456 24608
rect 42432 24692 42484 24744
rect 40408 24624 40460 24676
rect 39856 24556 39908 24608
rect 46848 24760 46900 24812
rect 48964 24760 49016 24812
rect 49516 24760 49568 24812
rect 51540 24760 51592 24812
rect 55496 24760 55548 24812
rect 56876 24828 56928 24880
rect 57336 24760 57388 24812
rect 45008 24735 45060 24744
rect 45008 24701 45017 24735
rect 45017 24701 45051 24735
rect 45051 24701 45060 24735
rect 45008 24692 45060 24701
rect 54116 24735 54168 24744
rect 54116 24701 54125 24735
rect 54125 24701 54159 24735
rect 54159 24701 54168 24735
rect 54116 24692 54168 24701
rect 46296 24624 46348 24676
rect 45928 24556 45980 24608
rect 49700 24556 49752 24608
rect 56692 24556 56744 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 6368 24352 6420 24404
rect 11520 24352 11572 24404
rect 12440 24352 12492 24404
rect 13452 24395 13504 24404
rect 13452 24361 13461 24395
rect 13461 24361 13495 24395
rect 13495 24361 13504 24395
rect 13452 24352 13504 24361
rect 25320 24352 25372 24404
rect 30932 24395 30984 24404
rect 30932 24361 30941 24395
rect 30941 24361 30975 24395
rect 30975 24361 30984 24395
rect 30932 24352 30984 24361
rect 32588 24352 32640 24404
rect 38016 24352 38068 24404
rect 41144 24352 41196 24404
rect 1860 24259 1912 24268
rect 1860 24225 1869 24259
rect 1869 24225 1903 24259
rect 1903 24225 1912 24259
rect 1860 24216 1912 24225
rect 15476 24259 15528 24268
rect 15476 24225 15485 24259
rect 15485 24225 15519 24259
rect 15519 24225 15528 24259
rect 15476 24216 15528 24225
rect 31392 24259 31444 24268
rect 31392 24225 31401 24259
rect 31401 24225 31435 24259
rect 31435 24225 31444 24259
rect 31392 24216 31444 24225
rect 33968 24216 34020 24268
rect 3332 24148 3384 24200
rect 9220 24148 9272 24200
rect 10416 24148 10468 24200
rect 12072 24191 12124 24200
rect 5264 24123 5316 24132
rect 5264 24089 5273 24123
rect 5273 24089 5307 24123
rect 5307 24089 5316 24123
rect 5264 24080 5316 24089
rect 3240 24055 3292 24064
rect 3240 24021 3249 24055
rect 3249 24021 3283 24055
rect 3283 24021 3292 24055
rect 3240 24012 3292 24021
rect 10692 24055 10744 24064
rect 10692 24021 10701 24055
rect 10701 24021 10735 24055
rect 10735 24021 10744 24055
rect 10692 24012 10744 24021
rect 11520 24012 11572 24064
rect 12072 24157 12081 24191
rect 12081 24157 12115 24191
rect 12115 24157 12124 24191
rect 12072 24148 12124 24157
rect 16120 24148 16172 24200
rect 17316 24191 17368 24200
rect 17316 24157 17325 24191
rect 17325 24157 17359 24191
rect 17359 24157 17368 24191
rect 17316 24148 17368 24157
rect 18696 24148 18748 24200
rect 13268 24080 13320 24132
rect 19340 24080 19392 24132
rect 21180 24148 21232 24200
rect 21824 24148 21876 24200
rect 24492 24148 24544 24200
rect 26240 24191 26292 24200
rect 26240 24157 26249 24191
rect 26249 24157 26283 24191
rect 26283 24157 26292 24191
rect 26240 24148 26292 24157
rect 27620 24148 27672 24200
rect 30288 24148 30340 24200
rect 23112 24080 23164 24132
rect 30932 24080 30984 24132
rect 31208 24080 31260 24132
rect 41420 24216 41472 24268
rect 42432 24352 42484 24404
rect 43076 24395 43128 24404
rect 43076 24361 43085 24395
rect 43085 24361 43119 24395
rect 43119 24361 43128 24395
rect 43076 24352 43128 24361
rect 48964 24395 49016 24404
rect 48964 24361 48973 24395
rect 48973 24361 49007 24395
rect 49007 24361 49016 24395
rect 48964 24352 49016 24361
rect 44916 24216 44968 24268
rect 54116 24352 54168 24404
rect 56508 24352 56560 24404
rect 56784 24352 56836 24404
rect 36084 24148 36136 24200
rect 35348 24080 35400 24132
rect 39028 24148 39080 24200
rect 39856 24191 39908 24200
rect 39856 24157 39865 24191
rect 39865 24157 39899 24191
rect 39899 24157 39908 24191
rect 39856 24148 39908 24157
rect 41236 24148 41288 24200
rect 43812 24148 43864 24200
rect 47584 24191 47636 24200
rect 47584 24157 47593 24191
rect 47593 24157 47627 24191
rect 47627 24157 47636 24191
rect 47584 24148 47636 24157
rect 48320 24148 48372 24200
rect 50160 24191 50212 24200
rect 50160 24157 50169 24191
rect 50169 24157 50203 24191
rect 50203 24157 50212 24191
rect 50160 24148 50212 24157
rect 41420 24080 41472 24132
rect 46848 24080 46900 24132
rect 48872 24080 48924 24132
rect 50804 24080 50856 24132
rect 14096 24012 14148 24064
rect 16856 24055 16908 24064
rect 16856 24021 16865 24055
rect 16865 24021 16899 24055
rect 16899 24021 16908 24055
rect 16856 24012 16908 24021
rect 18696 24055 18748 24064
rect 18696 24021 18705 24055
rect 18705 24021 18739 24055
rect 18739 24021 18748 24055
rect 18696 24012 18748 24021
rect 20812 24055 20864 24064
rect 20812 24021 20821 24055
rect 20821 24021 20855 24055
rect 20855 24021 20864 24055
rect 20812 24012 20864 24021
rect 22652 24055 22704 24064
rect 22652 24021 22661 24055
rect 22661 24021 22695 24055
rect 22695 24021 22704 24055
rect 22652 24012 22704 24021
rect 27620 24055 27672 24064
rect 27620 24021 27629 24055
rect 27629 24021 27663 24055
rect 27663 24021 27672 24055
rect 27620 24012 27672 24021
rect 36084 24055 36136 24064
rect 36084 24021 36093 24055
rect 36093 24021 36127 24055
rect 36127 24021 36136 24055
rect 36084 24012 36136 24021
rect 46388 24055 46440 24064
rect 46388 24021 46397 24055
rect 46397 24021 46431 24055
rect 46431 24021 46440 24055
rect 46388 24012 46440 24021
rect 49424 24055 49476 24064
rect 49424 24021 49433 24055
rect 49433 24021 49467 24055
rect 49467 24021 49476 24055
rect 49424 24012 49476 24021
rect 49976 24012 50028 24064
rect 51540 24055 51592 24064
rect 51540 24021 51549 24055
rect 51549 24021 51583 24055
rect 51583 24021 51592 24055
rect 51540 24012 51592 24021
rect 54484 24055 54536 24064
rect 54484 24021 54493 24055
rect 54493 24021 54527 24055
rect 54527 24021 54536 24055
rect 54484 24012 54536 24021
rect 56784 24080 56836 24132
rect 57244 24080 57296 24132
rect 58532 24055 58584 24064
rect 58532 24021 58541 24055
rect 58541 24021 58575 24055
rect 58575 24021 58584 24055
rect 58532 24012 58584 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 6092 23808 6144 23860
rect 13268 23851 13320 23860
rect 13268 23817 13277 23851
rect 13277 23817 13311 23851
rect 13311 23817 13320 23851
rect 13268 23808 13320 23817
rect 14096 23808 14148 23860
rect 3240 23740 3292 23792
rect 10692 23740 10744 23792
rect 18696 23740 18748 23792
rect 19248 23808 19300 23860
rect 23204 23851 23256 23860
rect 23204 23817 23213 23851
rect 23213 23817 23247 23851
rect 23247 23817 23256 23851
rect 23204 23808 23256 23817
rect 25504 23851 25556 23860
rect 25504 23817 25513 23851
rect 25513 23817 25547 23851
rect 25547 23817 25556 23851
rect 25504 23808 25556 23817
rect 28356 23851 28408 23860
rect 28356 23817 28365 23851
rect 28365 23817 28399 23851
rect 28399 23817 28408 23851
rect 28356 23808 28408 23817
rect 34520 23808 34572 23860
rect 36176 23808 36228 23860
rect 2228 23672 2280 23724
rect 6552 23672 6604 23724
rect 9312 23672 9364 23724
rect 13084 23672 13136 23724
rect 15752 23672 15804 23724
rect 19340 23672 19392 23724
rect 20812 23740 20864 23792
rect 22652 23740 22704 23792
rect 27620 23740 27672 23792
rect 29092 23783 29144 23792
rect 29092 23749 29126 23783
rect 29126 23749 29144 23783
rect 29092 23740 29144 23749
rect 32404 23783 32456 23792
rect 32404 23749 32438 23783
rect 32438 23749 32456 23783
rect 32404 23740 32456 23749
rect 36084 23740 36136 23792
rect 48872 23808 48924 23860
rect 50804 23851 50856 23860
rect 50804 23817 50813 23851
rect 50813 23817 50847 23851
rect 50847 23817 50856 23851
rect 50804 23808 50856 23817
rect 54760 23851 54812 23860
rect 54760 23817 54769 23851
rect 54769 23817 54803 23851
rect 54803 23817 54812 23851
rect 54760 23808 54812 23817
rect 57336 23851 57388 23860
rect 57336 23817 57345 23851
rect 57345 23817 57379 23851
rect 57379 23817 57388 23851
rect 57336 23808 57388 23817
rect 45928 23783 45980 23792
rect 20996 23672 21048 23724
rect 21824 23715 21876 23724
rect 21824 23681 21833 23715
rect 21833 23681 21867 23715
rect 21867 23681 21876 23715
rect 21824 23672 21876 23681
rect 25780 23672 25832 23724
rect 31392 23672 31444 23724
rect 3700 23511 3752 23520
rect 3700 23477 3709 23511
rect 3709 23477 3743 23511
rect 3743 23477 3752 23511
rect 3700 23468 3752 23477
rect 7012 23604 7064 23656
rect 9220 23604 9272 23656
rect 5172 23468 5224 23520
rect 8944 23511 8996 23520
rect 8944 23477 8953 23511
rect 8953 23477 8987 23511
rect 8987 23477 8996 23511
rect 8944 23468 8996 23477
rect 10784 23511 10836 23520
rect 10784 23477 10793 23511
rect 10793 23477 10827 23511
rect 10827 23477 10836 23511
rect 10784 23468 10836 23477
rect 13820 23604 13872 23656
rect 14740 23647 14792 23656
rect 14740 23613 14749 23647
rect 14749 23613 14783 23647
rect 14783 23613 14792 23647
rect 14740 23604 14792 23613
rect 24124 23647 24176 23656
rect 12072 23468 12124 23520
rect 12256 23468 12308 23520
rect 15476 23468 15528 23520
rect 16028 23468 16080 23520
rect 24124 23613 24133 23647
rect 24133 23613 24167 23647
rect 24167 23613 24176 23647
rect 24124 23604 24176 23613
rect 26240 23604 26292 23656
rect 33600 23672 33652 23724
rect 45928 23749 45962 23783
rect 45962 23749 45980 23783
rect 45928 23740 45980 23749
rect 49700 23783 49752 23792
rect 49700 23749 49734 23783
rect 49734 23749 49752 23783
rect 49700 23740 49752 23749
rect 54484 23740 54536 23792
rect 58532 23740 58584 23792
rect 40040 23672 40092 23724
rect 41696 23672 41748 23724
rect 44824 23672 44876 23724
rect 47584 23715 47636 23724
rect 33968 23647 34020 23656
rect 18052 23468 18104 23520
rect 18788 23511 18840 23520
rect 18788 23477 18797 23511
rect 18797 23477 18831 23511
rect 18831 23477 18840 23511
rect 18788 23468 18840 23477
rect 27620 23468 27672 23520
rect 33968 23613 33977 23647
rect 33977 23613 34011 23647
rect 34011 23613 34020 23647
rect 33968 23604 34020 23613
rect 37648 23604 37700 23656
rect 30196 23511 30248 23520
rect 30196 23477 30205 23511
rect 30205 23477 30239 23511
rect 30239 23477 30248 23511
rect 30196 23468 30248 23477
rect 38200 23468 38252 23520
rect 43076 23604 43128 23656
rect 45560 23604 45612 23656
rect 47584 23681 47593 23715
rect 47593 23681 47627 23715
rect 47627 23681 47636 23715
rect 47584 23672 47636 23681
rect 49332 23672 49384 23724
rect 49516 23672 49568 23724
rect 50160 23672 50212 23724
rect 53380 23715 53432 23724
rect 53380 23681 53389 23715
rect 53389 23681 53423 23715
rect 53423 23681 53432 23715
rect 53380 23672 53432 23681
rect 56784 23672 56836 23724
rect 41420 23468 41472 23520
rect 45192 23511 45244 23520
rect 45192 23477 45201 23511
rect 45201 23477 45235 23511
rect 45235 23477 45244 23511
rect 45192 23468 45244 23477
rect 47032 23511 47084 23520
rect 47032 23477 47041 23511
rect 47041 23477 47075 23511
rect 47075 23477 47084 23511
rect 47032 23468 47084 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 6552 23307 6604 23316
rect 6552 23273 6561 23307
rect 6561 23273 6595 23307
rect 6595 23273 6604 23307
rect 6552 23264 6604 23273
rect 8024 23264 8076 23316
rect 15752 23264 15804 23316
rect 18512 23264 18564 23316
rect 25780 23307 25832 23316
rect 25780 23273 25789 23307
rect 25789 23273 25823 23307
rect 25823 23273 25832 23307
rect 25780 23264 25832 23273
rect 27712 23264 27764 23316
rect 40592 23264 40644 23316
rect 46848 23264 46900 23316
rect 48320 23264 48372 23316
rect 49332 23307 49384 23316
rect 49332 23273 49341 23307
rect 49341 23273 49375 23307
rect 49375 23273 49384 23307
rect 49332 23264 49384 23273
rect 5172 23171 5224 23180
rect 5172 23137 5181 23171
rect 5181 23137 5215 23171
rect 5215 23137 5224 23171
rect 5172 23128 5224 23137
rect 12256 23128 12308 23180
rect 13728 23128 13780 23180
rect 15476 23171 15528 23180
rect 15476 23137 15485 23171
rect 15485 23137 15519 23171
rect 15519 23137 15528 23171
rect 15476 23128 15528 23137
rect 17316 23171 17368 23180
rect 17316 23137 17325 23171
rect 17325 23137 17359 23171
rect 17359 23137 17368 23171
rect 17316 23128 17368 23137
rect 30380 23128 30432 23180
rect 30840 23128 30892 23180
rect 3700 23060 3752 23112
rect 6184 23060 6236 23112
rect 7012 23103 7064 23112
rect 7012 23069 7021 23103
rect 7021 23069 7055 23103
rect 7055 23069 7064 23103
rect 7012 23060 7064 23069
rect 8944 23060 8996 23112
rect 9220 23060 9272 23112
rect 10784 23060 10836 23112
rect 16856 23060 16908 23112
rect 18788 23060 18840 23112
rect 21088 23103 21140 23112
rect 2228 22992 2280 23044
rect 11520 22992 11572 23044
rect 18052 22992 18104 23044
rect 21088 23069 21097 23103
rect 21097 23069 21131 23103
rect 21131 23069 21140 23103
rect 21088 23060 21140 23069
rect 24124 23060 24176 23112
rect 21180 22992 21232 23044
rect 22836 22992 22888 23044
rect 25136 22992 25188 23044
rect 27896 23060 27948 23112
rect 47584 23128 47636 23180
rect 32772 23103 32824 23112
rect 32772 23069 32781 23103
rect 32781 23069 32815 23103
rect 32815 23069 32824 23103
rect 32772 23060 32824 23069
rect 36084 23060 36136 23112
rect 37648 23103 37700 23112
rect 37648 23069 37657 23103
rect 37657 23069 37691 23103
rect 37691 23069 37700 23103
rect 37648 23060 37700 23069
rect 40408 23060 40460 23112
rect 40592 23103 40644 23112
rect 40592 23069 40601 23103
rect 40601 23069 40635 23103
rect 40635 23069 40644 23103
rect 40592 23060 40644 23069
rect 43076 23103 43128 23112
rect 27620 22992 27672 23044
rect 31852 22992 31904 23044
rect 34796 22992 34848 23044
rect 36544 22992 36596 23044
rect 39304 22992 39356 23044
rect 40316 22992 40368 23044
rect 43076 23069 43085 23103
rect 43085 23069 43119 23103
rect 43119 23069 43128 23103
rect 43076 23060 43128 23069
rect 45560 23103 45612 23112
rect 45560 23069 45569 23103
rect 45569 23069 45603 23103
rect 45603 23069 45612 23103
rect 45560 23060 45612 23069
rect 47032 23060 47084 23112
rect 42432 22992 42484 23044
rect 44180 22992 44232 23044
rect 49608 22992 49660 23044
rect 51540 23060 51592 23112
rect 53380 23060 53432 23112
rect 56784 23060 56836 23112
rect 50620 22992 50672 23044
rect 52092 22992 52144 23044
rect 58440 22992 58492 23044
rect 3240 22967 3292 22976
rect 3240 22933 3249 22967
rect 3249 22933 3283 22967
rect 3283 22933 3292 22967
rect 3240 22924 3292 22933
rect 10692 22967 10744 22976
rect 10692 22933 10701 22967
rect 10701 22933 10735 22967
rect 10735 22933 10744 22967
rect 10692 22924 10744 22933
rect 22100 22924 22152 22976
rect 22468 22967 22520 22976
rect 22468 22933 22477 22967
rect 22477 22933 22511 22967
rect 22511 22933 22520 22967
rect 22468 22924 22520 22933
rect 32312 22967 32364 22976
rect 32312 22933 32321 22967
rect 32321 22933 32355 22967
rect 32355 22933 32364 22967
rect 32312 22924 32364 22933
rect 33508 22924 33560 22976
rect 36636 22967 36688 22976
rect 36636 22933 36645 22967
rect 36645 22933 36679 22967
rect 36679 22933 36688 22967
rect 36636 22924 36688 22933
rect 37372 22924 37424 22976
rect 40132 22924 40184 22976
rect 42064 22924 42116 22976
rect 42616 22967 42668 22976
rect 42616 22933 42625 22967
rect 42625 22933 42659 22967
rect 42659 22933 42668 22967
rect 42616 22924 42668 22933
rect 44456 22967 44508 22976
rect 44456 22933 44465 22967
rect 44465 22933 44499 22967
rect 44499 22933 44508 22967
rect 44456 22924 44508 22933
rect 51540 22967 51592 22976
rect 51540 22933 51549 22967
rect 51549 22933 51583 22967
rect 51583 22933 51592 22967
rect 51540 22924 51592 22933
rect 52736 22924 52788 22976
rect 58532 22967 58584 22976
rect 58532 22933 58541 22967
rect 58541 22933 58575 22967
rect 58575 22933 58584 22967
rect 58532 22924 58584 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 9312 22720 9364 22772
rect 13084 22763 13136 22772
rect 13084 22729 13093 22763
rect 13093 22729 13127 22763
rect 13127 22729 13136 22763
rect 13084 22720 13136 22729
rect 3240 22652 3292 22704
rect 10692 22652 10744 22704
rect 2228 22627 2280 22636
rect 2228 22593 2237 22627
rect 2237 22593 2271 22627
rect 2271 22593 2280 22627
rect 2228 22584 2280 22593
rect 9220 22627 9272 22636
rect 9220 22593 9229 22627
rect 9229 22593 9263 22627
rect 9263 22593 9272 22627
rect 12256 22652 12308 22704
rect 9220 22584 9272 22593
rect 12900 22584 12952 22636
rect 15476 22652 15528 22704
rect 15752 22584 15804 22636
rect 18052 22584 18104 22636
rect 20628 22584 20680 22636
rect 20996 22584 21048 22636
rect 22468 22652 22520 22704
rect 23112 22720 23164 22772
rect 25136 22763 25188 22772
rect 21732 22584 21784 22636
rect 24124 22652 24176 22704
rect 25136 22729 25145 22763
rect 25145 22729 25179 22763
rect 25179 22729 25188 22763
rect 25136 22720 25188 22729
rect 30932 22763 30984 22772
rect 25780 22584 25832 22636
rect 25964 22516 26016 22568
rect 27804 22652 27856 22704
rect 30196 22652 30248 22704
rect 30932 22729 30941 22763
rect 30941 22729 30975 22763
rect 30975 22729 30984 22763
rect 30932 22720 30984 22729
rect 44824 22720 44876 22772
rect 49608 22763 49660 22772
rect 49608 22729 49617 22763
rect 49617 22729 49651 22763
rect 49651 22729 49660 22763
rect 49608 22720 49660 22729
rect 31116 22652 31168 22704
rect 32772 22584 32824 22636
rect 34152 22584 34204 22636
rect 35348 22627 35400 22636
rect 35348 22593 35357 22627
rect 35357 22593 35391 22627
rect 35391 22593 35400 22627
rect 35348 22584 35400 22593
rect 37464 22584 37516 22636
rect 3608 22423 3660 22432
rect 3608 22389 3617 22423
rect 3617 22389 3651 22423
rect 3651 22389 3660 22423
rect 3608 22380 3660 22389
rect 16120 22423 16172 22432
rect 16120 22389 16129 22423
rect 16129 22389 16163 22423
rect 16163 22389 16172 22423
rect 16120 22380 16172 22389
rect 20812 22380 20864 22432
rect 20904 22423 20956 22432
rect 20904 22389 20913 22423
rect 20913 22389 20947 22423
rect 20947 22389 20956 22423
rect 20904 22380 20956 22389
rect 27620 22380 27672 22432
rect 37648 22516 37700 22568
rect 45192 22652 45244 22704
rect 50620 22720 50672 22772
rect 57244 22763 57296 22772
rect 57244 22729 57253 22763
rect 57253 22729 57287 22763
rect 57287 22729 57296 22763
rect 57244 22720 57296 22729
rect 40224 22584 40276 22636
rect 40316 22627 40368 22636
rect 40316 22593 40325 22627
rect 40325 22593 40359 22627
rect 40359 22593 40368 22627
rect 40316 22584 40368 22593
rect 41880 22584 41932 22636
rect 43076 22584 43128 22636
rect 46388 22584 46440 22636
rect 51540 22652 51592 22704
rect 58532 22652 58584 22704
rect 49700 22584 49752 22636
rect 50160 22627 50212 22636
rect 50160 22593 50169 22627
rect 50169 22593 50203 22627
rect 50203 22593 50212 22627
rect 50160 22584 50212 22593
rect 55956 22584 56008 22636
rect 34520 22380 34572 22432
rect 36728 22423 36780 22432
rect 36728 22389 36737 22423
rect 36737 22389 36771 22423
rect 36771 22389 36780 22423
rect 36728 22380 36780 22389
rect 39856 22423 39908 22432
rect 39856 22389 39865 22423
rect 39865 22389 39899 22423
rect 39899 22389 39908 22423
rect 39856 22380 39908 22389
rect 41696 22423 41748 22432
rect 41696 22389 41705 22423
rect 41705 22389 41739 22423
rect 41739 22389 41748 22423
rect 41696 22380 41748 22389
rect 42064 22380 42116 22432
rect 42800 22380 42852 22432
rect 44364 22423 44416 22432
rect 44364 22389 44373 22423
rect 44373 22389 44407 22423
rect 44407 22389 44416 22423
rect 44364 22380 44416 22389
rect 52000 22516 52052 22568
rect 55128 22448 55180 22500
rect 45560 22380 45612 22432
rect 51172 22380 51224 22432
rect 55404 22380 55456 22432
rect 56784 22380 56836 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 20628 22219 20680 22228
rect 20628 22185 20637 22219
rect 20637 22185 20671 22219
rect 20671 22185 20680 22219
rect 20628 22176 20680 22185
rect 25780 22219 25832 22228
rect 25780 22185 25789 22219
rect 25789 22185 25823 22219
rect 25823 22185 25832 22219
rect 25780 22176 25832 22185
rect 31852 22176 31904 22228
rect 34152 22219 34204 22228
rect 34152 22185 34161 22219
rect 34161 22185 34195 22219
rect 34195 22185 34204 22219
rect 34152 22176 34204 22185
rect 37464 22219 37516 22228
rect 37464 22185 37473 22219
rect 37473 22185 37507 22219
rect 37507 22185 37516 22219
rect 37464 22176 37516 22185
rect 39304 22219 39356 22228
rect 39304 22185 39313 22219
rect 39313 22185 39347 22219
rect 39347 22185 39356 22219
rect 39304 22176 39356 22185
rect 42432 22176 42484 22228
rect 44180 22176 44232 22228
rect 52092 22176 52144 22228
rect 15476 22040 15528 22092
rect 3608 21972 3660 22024
rect 4436 21972 4488 22024
rect 5172 21972 5224 22024
rect 5448 21972 5500 22024
rect 12256 21972 12308 22024
rect 30840 22040 30892 22092
rect 15844 21972 15896 22024
rect 16028 22015 16080 22024
rect 16028 21981 16062 22015
rect 16062 21981 16080 22015
rect 16028 21972 16080 21981
rect 19156 21972 19208 22024
rect 21088 22015 21140 22024
rect 21088 21981 21097 22015
rect 21097 21981 21131 22015
rect 21131 21981 21140 22015
rect 21088 21972 21140 21981
rect 21732 21972 21784 22024
rect 27620 22015 27672 22024
rect 27620 21981 27629 22015
rect 27629 21981 27663 22015
rect 27663 21981 27672 22015
rect 27620 21972 27672 21981
rect 37648 22040 37700 22092
rect 36084 22015 36136 22024
rect 36084 21981 36093 22015
rect 36093 21981 36127 22015
rect 36127 21981 36136 22015
rect 36084 21972 36136 21981
rect 37372 21972 37424 22024
rect 38200 22015 38252 22024
rect 38200 21981 38234 22015
rect 38234 21981 38252 22015
rect 38200 21972 38252 21981
rect 40316 21972 40368 22024
rect 44364 21972 44416 22024
rect 49976 21972 50028 22024
rect 50620 22015 50672 22024
rect 50620 21981 50629 22015
rect 50629 21981 50663 22015
rect 50663 21981 50672 22015
rect 50620 21972 50672 21981
rect 51172 21972 51224 22024
rect 52736 22015 52788 22024
rect 52736 21981 52770 22015
rect 52770 21981 52788 22015
rect 2228 21904 2280 21956
rect 3424 21904 3476 21956
rect 13268 21904 13320 21956
rect 20536 21904 20588 21956
rect 23204 21904 23256 21956
rect 25136 21904 25188 21956
rect 28908 21904 28960 21956
rect 3240 21879 3292 21888
rect 3240 21845 3249 21879
rect 3249 21845 3283 21879
rect 3283 21845 3292 21879
rect 3240 21836 3292 21845
rect 5172 21879 5224 21888
rect 5172 21845 5181 21879
rect 5181 21845 5215 21879
rect 5215 21845 5224 21879
rect 5172 21836 5224 21845
rect 12992 21879 13044 21888
rect 12992 21845 13001 21879
rect 13001 21845 13035 21879
rect 13035 21845 13044 21879
rect 12992 21836 13044 21845
rect 15752 21836 15804 21888
rect 21180 21836 21232 21888
rect 29000 21879 29052 21888
rect 29000 21845 29009 21879
rect 29009 21845 29043 21879
rect 29043 21845 29052 21879
rect 29000 21836 29052 21845
rect 36268 21904 36320 21956
rect 44088 21904 44140 21956
rect 50988 21904 51040 21956
rect 52736 21972 52788 21981
rect 55680 21972 55732 22024
rect 56416 21972 56468 22024
rect 33876 21836 33928 21888
rect 47584 21879 47636 21888
rect 47584 21845 47593 21879
rect 47593 21845 47627 21879
rect 47627 21845 47636 21879
rect 47584 21836 47636 21845
rect 53840 21879 53892 21888
rect 53840 21845 53849 21879
rect 53849 21845 53883 21879
rect 53883 21845 53892 21879
rect 53840 21836 53892 21845
rect 56784 21836 56836 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 3424 21675 3476 21684
rect 3424 21641 3433 21675
rect 3433 21641 3467 21675
rect 3467 21641 3476 21675
rect 3424 21632 3476 21641
rect 3240 21564 3292 21616
rect 5172 21564 5224 21616
rect 22836 21632 22888 21684
rect 25136 21675 25188 21684
rect 25136 21641 25145 21675
rect 25145 21641 25179 21675
rect 25179 21641 25188 21675
rect 25136 21632 25188 21641
rect 28908 21632 28960 21684
rect 34796 21632 34848 21684
rect 36544 21632 36596 21684
rect 40040 21675 40092 21684
rect 40040 21641 40049 21675
rect 40049 21641 40083 21675
rect 40083 21641 40092 21675
rect 40040 21632 40092 21641
rect 41880 21675 41932 21684
rect 41880 21641 41889 21675
rect 41889 21641 41923 21675
rect 41923 21641 41932 21675
rect 41880 21632 41932 21641
rect 49700 21675 49752 21684
rect 49700 21641 49709 21675
rect 49709 21641 49743 21675
rect 49743 21641 49752 21675
rect 49700 21632 49752 21641
rect 22100 21607 22152 21616
rect 22100 21573 22134 21607
rect 22134 21573 22152 21607
rect 22100 21564 22152 21573
rect 32312 21564 32364 21616
rect 34520 21564 34572 21616
rect 2136 21496 2188 21548
rect 4436 21496 4488 21548
rect 9588 21496 9640 21548
rect 12256 21539 12308 21548
rect 12256 21505 12265 21539
rect 12265 21505 12299 21539
rect 12299 21505 12308 21539
rect 12256 21496 12308 21505
rect 14464 21496 14516 21548
rect 14740 21539 14792 21548
rect 14740 21505 14749 21539
rect 14749 21505 14783 21539
rect 14783 21505 14792 21539
rect 14740 21496 14792 21505
rect 16488 21496 16540 21548
rect 18052 21496 18104 21548
rect 18420 21496 18472 21548
rect 20628 21496 20680 21548
rect 21732 21496 21784 21548
rect 25780 21496 25832 21548
rect 28816 21496 28868 21548
rect 30012 21496 30064 21548
rect 30840 21496 30892 21548
rect 36084 21564 36136 21616
rect 37556 21496 37608 21548
rect 39856 21564 39908 21616
rect 42616 21564 42668 21616
rect 42800 21607 42852 21616
rect 42800 21573 42809 21607
rect 42809 21573 42843 21607
rect 42843 21573 42852 21607
rect 42800 21564 42852 21573
rect 53840 21564 53892 21616
rect 40316 21496 40368 21548
rect 44180 21496 44232 21548
rect 50068 21496 50120 21548
rect 51540 21496 51592 21548
rect 55128 21496 55180 21548
rect 56692 21496 56744 21548
rect 7012 21471 7064 21480
rect 7012 21437 7021 21471
rect 7021 21437 7055 21471
rect 7055 21437 7064 21471
rect 7012 21428 7064 21437
rect 15844 21428 15896 21480
rect 27620 21471 27672 21480
rect 4896 21292 4948 21344
rect 8484 21292 8536 21344
rect 13636 21335 13688 21344
rect 13636 21301 13645 21335
rect 13645 21301 13679 21335
rect 13679 21301 13688 21335
rect 13636 21292 13688 21301
rect 18052 21335 18104 21344
rect 18052 21301 18061 21335
rect 18061 21301 18095 21335
rect 18095 21301 18104 21335
rect 18052 21292 18104 21301
rect 19892 21335 19944 21344
rect 19892 21301 19901 21335
rect 19901 21301 19935 21335
rect 19935 21301 19944 21335
rect 19892 21292 19944 21301
rect 27620 21437 27629 21471
rect 27629 21437 27663 21471
rect 27663 21437 27672 21471
rect 27620 21428 27672 21437
rect 24492 21292 24544 21344
rect 31576 21335 31628 21344
rect 31576 21301 31585 21335
rect 31585 21301 31619 21335
rect 31619 21301 31628 21335
rect 31576 21292 31628 21301
rect 42432 21292 42484 21344
rect 46388 21335 46440 21344
rect 46388 21301 46397 21335
rect 46397 21301 46431 21335
rect 46431 21301 46440 21335
rect 46388 21292 46440 21301
rect 52000 21292 52052 21344
rect 54576 21335 54628 21344
rect 54576 21301 54585 21335
rect 54585 21301 54619 21335
rect 54619 21301 54628 21335
rect 54576 21292 54628 21301
rect 57244 21292 57296 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 5448 21131 5500 21140
rect 5448 21097 5457 21131
rect 5457 21097 5491 21131
rect 5491 21097 5500 21131
rect 5448 21088 5500 21097
rect 4344 21020 4396 21072
rect 12256 21088 12308 21140
rect 13268 21131 13320 21140
rect 13268 21097 13277 21131
rect 13277 21097 13311 21131
rect 13311 21097 13320 21131
rect 13268 21088 13320 21097
rect 14740 20952 14792 21004
rect 15844 21088 15896 21140
rect 16488 21131 16540 21140
rect 16488 21097 16497 21131
rect 16497 21097 16531 21131
rect 16531 21097 16540 21131
rect 16488 21088 16540 21097
rect 18420 21131 18472 21140
rect 18420 21097 18429 21131
rect 18429 21097 18463 21131
rect 18463 21097 18472 21131
rect 18420 21088 18472 21097
rect 20536 21088 20588 21140
rect 25780 21131 25832 21140
rect 25780 21097 25789 21131
rect 25789 21097 25823 21131
rect 25823 21097 25832 21131
rect 25780 21088 25832 21097
rect 19248 20995 19300 21004
rect 19248 20961 19257 20995
rect 19257 20961 19291 20995
rect 19291 20961 19300 20995
rect 19248 20952 19300 20961
rect 6368 20927 6420 20936
rect 6368 20893 6377 20927
rect 6377 20893 6411 20927
rect 6411 20893 6420 20927
rect 6368 20884 6420 20893
rect 7012 20884 7064 20936
rect 8208 20884 8260 20936
rect 8944 20927 8996 20936
rect 8944 20893 8953 20927
rect 8953 20893 8987 20927
rect 8987 20893 8996 20927
rect 8944 20884 8996 20893
rect 13636 20884 13688 20936
rect 16120 20884 16172 20936
rect 19892 20884 19944 20936
rect 21088 20927 21140 20936
rect 21088 20893 21097 20927
rect 21097 20893 21131 20927
rect 21131 20893 21140 20927
rect 21088 20884 21140 20893
rect 24492 20884 24544 20936
rect 26976 20884 27028 20936
rect 27620 21088 27672 21140
rect 28816 21131 28868 21140
rect 28816 21097 28825 21131
rect 28825 21097 28859 21131
rect 28859 21097 28868 21131
rect 28816 21088 28868 21097
rect 37556 21131 37608 21140
rect 37556 21097 37565 21131
rect 37565 21097 37599 21131
rect 37599 21097 37608 21131
rect 37556 21088 37608 21097
rect 40224 21088 40276 21140
rect 44088 21131 44140 21140
rect 44088 21097 44097 21131
rect 44097 21097 44131 21131
rect 44131 21097 44140 21131
rect 44088 21088 44140 21097
rect 51540 21131 51592 21140
rect 51540 21097 51549 21131
rect 51549 21097 51583 21131
rect 51583 21097 51592 21131
rect 51540 21088 51592 21097
rect 56692 21131 56744 21140
rect 56692 21097 56701 21131
rect 56701 21097 56735 21131
rect 56735 21097 56744 21131
rect 56692 21088 56744 21097
rect 58440 21088 58492 21140
rect 30012 20995 30064 21004
rect 30012 20961 30021 20995
rect 30021 20961 30055 20995
rect 30055 20961 30064 20995
rect 30012 20952 30064 20961
rect 52000 20995 52052 21004
rect 52000 20961 52009 20995
rect 52009 20961 52043 20995
rect 52043 20961 52052 20995
rect 52000 20952 52052 20961
rect 31576 20884 31628 20936
rect 32956 20884 33008 20936
rect 34980 20884 35032 20936
rect 36084 20884 36136 20936
rect 36728 20884 36780 20936
rect 5264 20816 5316 20868
rect 5816 20816 5868 20868
rect 7656 20816 7708 20868
rect 10232 20816 10284 20868
rect 7748 20791 7800 20800
rect 7748 20757 7757 20791
rect 7757 20757 7791 20791
rect 7791 20757 7800 20791
rect 7748 20748 7800 20757
rect 9680 20748 9732 20800
rect 20812 20816 20864 20868
rect 25688 20816 25740 20868
rect 28908 20816 28960 20868
rect 41696 20884 41748 20936
rect 42432 20884 42484 20936
rect 44456 20884 44508 20936
rect 45560 20884 45612 20936
rect 47584 20884 47636 20936
rect 50160 20927 50212 20936
rect 50160 20893 50169 20927
rect 50169 20893 50203 20927
rect 50203 20893 50212 20927
rect 50160 20884 50212 20893
rect 50988 20884 51040 20936
rect 54576 20884 54628 20936
rect 55312 20927 55364 20936
rect 55312 20893 55321 20927
rect 55321 20893 55355 20927
rect 55355 20893 55364 20927
rect 55312 20884 55364 20893
rect 56784 20884 56836 20936
rect 40316 20816 40368 20868
rect 46756 20816 46808 20868
rect 48596 20816 48648 20868
rect 50804 20816 50856 20868
rect 56692 20816 56744 20868
rect 58440 20816 58492 20868
rect 20904 20748 20956 20800
rect 22468 20791 22520 20800
rect 22468 20757 22477 20791
rect 22477 20757 22511 20791
rect 22511 20757 22520 20791
rect 22468 20748 22520 20757
rect 31392 20791 31444 20800
rect 31392 20757 31401 20791
rect 31401 20757 31435 20791
rect 31435 20757 31444 20791
rect 31392 20748 31444 20757
rect 32496 20748 32548 20800
rect 47308 20748 47360 20800
rect 48872 20791 48924 20800
rect 48872 20757 48881 20791
rect 48881 20757 48915 20791
rect 48915 20757 48924 20791
rect 48872 20748 48924 20757
rect 52552 20748 52604 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 7656 20544 7708 20596
rect 9588 20587 9640 20596
rect 9588 20553 9597 20587
rect 9597 20553 9631 20587
rect 9631 20553 9640 20587
rect 9588 20544 9640 20553
rect 20628 20544 20680 20596
rect 23204 20587 23256 20596
rect 23204 20553 23213 20587
rect 23213 20553 23247 20587
rect 23247 20553 23256 20587
rect 23204 20544 23256 20553
rect 33876 20587 33928 20596
rect 33876 20553 33885 20587
rect 33885 20553 33919 20587
rect 33919 20553 33928 20587
rect 33876 20544 33928 20553
rect 4896 20408 4948 20460
rect 5540 20408 5592 20460
rect 8944 20476 8996 20528
rect 12992 20476 13044 20528
rect 18052 20476 18104 20528
rect 8300 20408 8352 20460
rect 14740 20451 14792 20460
rect 14740 20417 14749 20451
rect 14749 20417 14783 20451
rect 14783 20417 14792 20451
rect 14740 20408 14792 20417
rect 18696 20408 18748 20460
rect 19340 20408 19392 20460
rect 21088 20476 21140 20528
rect 22468 20476 22520 20528
rect 29000 20476 29052 20528
rect 20628 20408 20680 20460
rect 21732 20408 21784 20460
rect 28540 20408 28592 20460
rect 30012 20408 30064 20460
rect 32128 20408 32180 20460
rect 4068 20340 4120 20392
rect 4344 20383 4396 20392
rect 4344 20349 4353 20383
rect 4353 20349 4387 20383
rect 4387 20349 4396 20383
rect 4344 20340 4396 20349
rect 6368 20383 6420 20392
rect 6368 20349 6377 20383
rect 6377 20349 6411 20383
rect 6411 20349 6420 20383
rect 6368 20340 6420 20349
rect 11612 20383 11664 20392
rect 11612 20349 11621 20383
rect 11621 20349 11655 20383
rect 11655 20349 11664 20383
rect 11612 20340 11664 20349
rect 24492 20383 24544 20392
rect 12900 20272 12952 20324
rect 4068 20204 4120 20256
rect 5724 20247 5776 20256
rect 5724 20213 5733 20247
rect 5733 20213 5767 20247
rect 5767 20213 5776 20247
rect 5724 20204 5776 20213
rect 16120 20247 16172 20256
rect 16120 20213 16129 20247
rect 16129 20213 16163 20247
rect 16163 20213 16172 20247
rect 16120 20204 16172 20213
rect 24492 20349 24501 20383
rect 24501 20349 24535 20383
rect 24535 20349 24544 20383
rect 24492 20340 24544 20349
rect 26976 20340 27028 20392
rect 33508 20476 33560 20528
rect 34980 20519 35032 20528
rect 34980 20485 34989 20519
rect 34989 20485 35023 20519
rect 35023 20485 35032 20519
rect 40132 20544 40184 20596
rect 44180 20544 44232 20596
rect 46756 20587 46808 20596
rect 46756 20553 46765 20587
rect 46765 20553 46799 20587
rect 46799 20553 46808 20587
rect 46756 20544 46808 20553
rect 50988 20544 51040 20596
rect 55956 20587 56008 20596
rect 34980 20476 35032 20485
rect 38660 20476 38712 20528
rect 49976 20519 50028 20528
rect 49976 20485 49985 20519
rect 49985 20485 50019 20519
rect 50019 20485 50028 20519
rect 49976 20476 50028 20485
rect 55956 20553 55965 20587
rect 55965 20553 55999 20587
rect 55999 20553 56008 20587
rect 55956 20544 56008 20553
rect 38752 20408 38804 20460
rect 40316 20408 40368 20460
rect 41788 20408 41840 20460
rect 43720 20408 43772 20460
rect 32496 20383 32548 20392
rect 32496 20349 32505 20383
rect 32505 20349 32539 20383
rect 32539 20349 32548 20383
rect 32496 20340 32548 20349
rect 42432 20383 42484 20392
rect 42432 20349 42441 20383
rect 42441 20349 42475 20383
rect 42475 20349 42484 20383
rect 42432 20340 42484 20349
rect 45100 20340 45152 20392
rect 45468 20408 45520 20460
rect 46572 20408 46624 20460
rect 47584 20408 47636 20460
rect 48964 20408 49016 20460
rect 52000 20340 52052 20392
rect 53380 20408 53432 20460
rect 54576 20451 54628 20460
rect 54576 20417 54585 20451
rect 54585 20417 54619 20451
rect 54619 20417 54628 20451
rect 54576 20408 54628 20417
rect 19156 20272 19208 20324
rect 19340 20204 19392 20256
rect 25872 20247 25924 20256
rect 25872 20213 25881 20247
rect 25881 20213 25915 20247
rect 25915 20213 25924 20247
rect 25872 20204 25924 20213
rect 28724 20247 28776 20256
rect 28724 20213 28733 20247
rect 28733 20213 28767 20247
rect 28767 20213 28776 20247
rect 28724 20204 28776 20213
rect 32680 20204 32732 20256
rect 36084 20204 36136 20256
rect 38844 20204 38896 20256
rect 41420 20204 41472 20256
rect 50252 20204 50304 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 14464 20000 14516 20052
rect 18696 20043 18748 20052
rect 18696 20009 18705 20043
rect 18705 20009 18739 20043
rect 18739 20009 18748 20043
rect 18696 20000 18748 20009
rect 20628 20043 20680 20052
rect 20628 20009 20637 20043
rect 20637 20009 20671 20043
rect 20671 20009 20680 20043
rect 20628 20000 20680 20009
rect 21732 20000 21784 20052
rect 25688 20000 25740 20052
rect 28540 20043 28592 20052
rect 28540 20009 28549 20043
rect 28549 20009 28583 20043
rect 28583 20009 28592 20043
rect 28540 20000 28592 20009
rect 32128 20043 32180 20052
rect 32128 20009 32137 20043
rect 32137 20009 32171 20043
rect 32171 20009 32180 20043
rect 32128 20000 32180 20009
rect 14096 19864 14148 19916
rect 14740 19864 14792 19916
rect 30012 19864 30064 19916
rect 32128 19864 32180 19916
rect 36084 20000 36136 20052
rect 36268 20043 36320 20052
rect 36268 20009 36277 20043
rect 36277 20009 36311 20043
rect 36311 20009 36320 20043
rect 36268 20000 36320 20009
rect 43720 20043 43772 20052
rect 43720 20009 43729 20043
rect 43729 20009 43763 20043
rect 43763 20009 43772 20043
rect 43720 20000 43772 20009
rect 46572 20043 46624 20052
rect 46572 20009 46581 20043
rect 46581 20009 46615 20043
rect 46615 20009 46624 20043
rect 46572 20000 46624 20009
rect 48596 20043 48648 20052
rect 48596 20009 48605 20043
rect 48605 20009 48639 20043
rect 48639 20009 48648 20043
rect 48596 20000 48648 20009
rect 53380 20043 53432 20052
rect 53380 20009 53389 20043
rect 53389 20009 53423 20043
rect 53423 20009 53432 20043
rect 53380 20000 53432 20009
rect 56692 20043 56744 20052
rect 56692 20009 56701 20043
rect 56701 20009 56735 20043
rect 56735 20009 56744 20043
rect 56692 20000 56744 20009
rect 58440 20000 58492 20052
rect 40316 19864 40368 19916
rect 50160 19907 50212 19916
rect 5724 19796 5776 19848
rect 5816 19796 5868 19848
rect 8944 19839 8996 19848
rect 8944 19805 8953 19839
rect 8953 19805 8987 19839
rect 8987 19805 8996 19839
rect 8944 19796 8996 19805
rect 11612 19796 11664 19848
rect 16120 19796 16172 19848
rect 17316 19839 17368 19848
rect 17316 19805 17325 19839
rect 17325 19805 17359 19839
rect 17359 19805 17368 19839
rect 17316 19796 17368 19805
rect 19248 19839 19300 19848
rect 19248 19805 19257 19839
rect 19257 19805 19291 19839
rect 19291 19805 19300 19839
rect 19248 19796 19300 19805
rect 19340 19796 19392 19848
rect 23664 19796 23716 19848
rect 24492 19796 24544 19848
rect 25872 19796 25924 19848
rect 26976 19796 27028 19848
rect 31392 19796 31444 19848
rect 32680 19796 32732 19848
rect 36636 19796 36688 19848
rect 38660 19796 38712 19848
rect 50160 19873 50169 19907
rect 50169 19873 50203 19907
rect 50203 19873 50212 19907
rect 50160 19864 50212 19873
rect 52000 19907 52052 19916
rect 52000 19873 52009 19907
rect 52009 19873 52043 19907
rect 52043 19873 52052 19907
rect 52000 19864 52052 19873
rect 42432 19796 42484 19848
rect 45100 19796 45152 19848
rect 47216 19839 47268 19848
rect 47216 19805 47225 19839
rect 47225 19805 47259 19839
rect 47259 19805 47268 19839
rect 47216 19796 47268 19805
rect 47308 19796 47360 19848
rect 50252 19796 50304 19848
rect 52552 19796 52604 19848
rect 54576 19796 54628 19848
rect 55312 19839 55364 19848
rect 55312 19805 55321 19839
rect 55321 19805 55355 19839
rect 55355 19805 55364 19839
rect 55312 19796 55364 19805
rect 55404 19796 55456 19848
rect 55864 19796 55916 19848
rect 57244 19796 57296 19848
rect 8208 19771 8260 19780
rect 8208 19737 8217 19771
rect 8217 19737 8251 19771
rect 8251 19737 8260 19771
rect 8208 19728 8260 19737
rect 9588 19728 9640 19780
rect 12808 19728 12860 19780
rect 18696 19728 18748 19780
rect 20904 19728 20956 19780
rect 25964 19728 26016 19780
rect 28356 19728 28408 19780
rect 39120 19728 39172 19780
rect 4620 19660 4672 19712
rect 5724 19703 5776 19712
rect 5724 19669 5733 19703
rect 5733 19669 5767 19703
rect 5767 19669 5776 19703
rect 5724 19660 5776 19669
rect 10324 19703 10376 19712
rect 10324 19669 10333 19703
rect 10333 19669 10367 19703
rect 10367 19669 10376 19703
rect 10324 19660 10376 19669
rect 12900 19703 12952 19712
rect 12900 19669 12909 19703
rect 12909 19669 12943 19703
rect 12943 19669 12952 19703
rect 12900 19660 12952 19669
rect 31760 19660 31812 19712
rect 37832 19660 37884 19712
rect 41880 19703 41932 19712
rect 41880 19669 41889 19703
rect 41889 19669 41923 19703
rect 41923 19669 41932 19703
rect 41880 19660 41932 19669
rect 43812 19728 43864 19780
rect 46572 19728 46624 19780
rect 46388 19660 46440 19712
rect 51540 19703 51592 19712
rect 51540 19669 51549 19703
rect 51549 19669 51583 19703
rect 51583 19669 51592 19703
rect 51540 19660 51592 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 9588 19499 9640 19508
rect 5724 19388 5776 19440
rect 7748 19388 7800 19440
rect 9588 19465 9597 19499
rect 9597 19465 9631 19499
rect 9631 19465 9640 19499
rect 9588 19456 9640 19465
rect 18696 19499 18748 19508
rect 18696 19465 18705 19499
rect 18705 19465 18739 19499
rect 18739 19465 18748 19499
rect 18696 19456 18748 19465
rect 19248 19456 19300 19508
rect 9680 19388 9732 19440
rect 12900 19388 12952 19440
rect 28356 19499 28408 19508
rect 1584 19363 1636 19372
rect 1584 19329 1593 19363
rect 1593 19329 1627 19363
rect 1627 19329 1636 19363
rect 4068 19363 4120 19372
rect 1584 19320 1636 19329
rect 4068 19329 4077 19363
rect 4077 19329 4111 19363
rect 4111 19329 4120 19363
rect 4068 19320 4120 19329
rect 5540 19320 5592 19372
rect 8208 19363 8260 19372
rect 8208 19329 8217 19363
rect 8217 19329 8251 19363
rect 8251 19329 8260 19363
rect 8208 19320 8260 19329
rect 8484 19363 8536 19372
rect 8484 19329 8518 19363
rect 8518 19329 8536 19363
rect 8484 19320 8536 19329
rect 11612 19320 11664 19372
rect 12716 19320 12768 19372
rect 12808 19320 12860 19372
rect 6368 19295 6420 19304
rect 6368 19261 6377 19295
rect 6377 19261 6411 19295
rect 6411 19261 6420 19295
rect 6368 19252 6420 19261
rect 13912 19320 13964 19372
rect 17316 19363 17368 19372
rect 17316 19329 17325 19363
rect 17325 19329 17359 19363
rect 17359 19329 17368 19363
rect 17316 19320 17368 19329
rect 19248 19320 19300 19372
rect 20720 19388 20772 19440
rect 28356 19465 28365 19499
rect 28365 19465 28399 19499
rect 28399 19465 28408 19499
rect 28356 19456 28408 19465
rect 31208 19388 31260 19440
rect 34520 19456 34572 19508
rect 43812 19499 43864 19508
rect 43812 19465 43821 19499
rect 43821 19465 43855 19499
rect 43855 19465 43864 19499
rect 43812 19456 43864 19465
rect 46572 19499 46624 19508
rect 46572 19465 46581 19499
rect 46581 19465 46615 19499
rect 46615 19465 46624 19499
rect 46572 19456 46624 19465
rect 48964 19499 49016 19508
rect 48964 19465 48973 19499
rect 48973 19465 49007 19499
rect 49007 19465 49016 19499
rect 48964 19456 49016 19465
rect 50804 19499 50856 19508
rect 50804 19465 50813 19499
rect 50813 19465 50847 19499
rect 50847 19465 50856 19499
rect 50804 19456 50856 19465
rect 21272 19320 21324 19372
rect 21824 19363 21876 19372
rect 21824 19329 21833 19363
rect 21833 19329 21867 19363
rect 21867 19329 21876 19363
rect 21824 19320 21876 19329
rect 23480 19320 23532 19372
rect 26976 19363 27028 19372
rect 26976 19329 26985 19363
rect 26985 19329 27019 19363
rect 27019 19329 27028 19363
rect 26976 19320 27028 19329
rect 30012 19320 30064 19372
rect 32220 19320 32272 19372
rect 36084 19388 36136 19440
rect 36728 19320 36780 19372
rect 39856 19388 39908 19440
rect 41880 19388 41932 19440
rect 48872 19388 48924 19440
rect 51540 19388 51592 19440
rect 55680 19388 55732 19440
rect 55864 19388 55916 19440
rect 23664 19295 23716 19304
rect 23664 19261 23673 19295
rect 23673 19261 23707 19295
rect 23707 19261 23716 19295
rect 23664 19252 23716 19261
rect 32128 19295 32180 19304
rect 32128 19261 32137 19295
rect 32137 19261 32171 19295
rect 32171 19261 32180 19295
rect 32128 19252 32180 19261
rect 38292 19252 38344 19304
rect 38660 19295 38712 19304
rect 38660 19261 38669 19295
rect 38669 19261 38703 19295
rect 38703 19261 38712 19295
rect 41236 19320 41288 19372
rect 41788 19320 41840 19372
rect 42432 19363 42484 19372
rect 38660 19252 38712 19261
rect 39856 19184 39908 19236
rect 42432 19329 42441 19363
rect 42441 19329 42475 19363
rect 42475 19329 42484 19363
rect 42432 19320 42484 19329
rect 43720 19320 43772 19372
rect 46480 19320 46532 19372
rect 47216 19320 47268 19372
rect 50160 19320 50212 19372
rect 45100 19252 45152 19304
rect 2964 19159 3016 19168
rect 2964 19125 2973 19159
rect 2973 19125 3007 19159
rect 3007 19125 3016 19159
rect 2964 19116 3016 19125
rect 7748 19159 7800 19168
rect 7748 19125 7757 19159
rect 7757 19125 7791 19159
rect 7791 19125 7800 19159
rect 7748 19116 7800 19125
rect 14004 19116 14056 19168
rect 23204 19159 23256 19168
rect 23204 19125 23213 19159
rect 23213 19125 23247 19159
rect 23247 19125 23256 19159
rect 23204 19116 23256 19125
rect 25044 19159 25096 19168
rect 25044 19125 25053 19159
rect 25053 19125 25087 19159
rect 25087 19125 25096 19159
rect 25044 19116 25096 19125
rect 33508 19159 33560 19168
rect 33508 19125 33517 19159
rect 33517 19125 33551 19159
rect 33551 19125 33560 19159
rect 33508 19116 33560 19125
rect 38660 19116 38712 19168
rect 41512 19116 41564 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 10232 18912 10284 18964
rect 32220 18912 32272 18964
rect 41236 18955 41288 18964
rect 41236 18921 41245 18955
rect 41245 18921 41279 18955
rect 41279 18921 41288 18955
rect 41236 18912 41288 18921
rect 43720 18955 43772 18964
rect 43720 18921 43729 18955
rect 43729 18921 43763 18955
rect 43763 18921 43772 18955
rect 43720 18912 43772 18921
rect 46480 18955 46532 18964
rect 46480 18921 46489 18955
rect 46489 18921 46523 18955
rect 46523 18921 46532 18955
rect 46480 18912 46532 18921
rect 1584 18819 1636 18828
rect 1584 18785 1593 18819
rect 1593 18785 1627 18819
rect 1627 18785 1636 18819
rect 1584 18776 1636 18785
rect 39856 18819 39908 18828
rect 39856 18785 39865 18819
rect 39865 18785 39899 18819
rect 39899 18785 39908 18819
rect 39856 18776 39908 18785
rect 2964 18708 3016 18760
rect 6368 18751 6420 18760
rect 6368 18717 6377 18751
rect 6377 18717 6411 18751
rect 6411 18717 6420 18751
rect 6368 18708 6420 18717
rect 7748 18708 7800 18760
rect 8944 18751 8996 18760
rect 8944 18717 8953 18751
rect 8953 18717 8987 18751
rect 8987 18717 8996 18751
rect 8944 18708 8996 18717
rect 10324 18708 10376 18760
rect 11520 18751 11572 18760
rect 11520 18717 11529 18751
rect 11529 18717 11563 18751
rect 11563 18717 11572 18751
rect 11520 18708 11572 18717
rect 11612 18708 11664 18760
rect 13912 18708 13964 18760
rect 20720 18751 20772 18760
rect 20720 18717 20729 18751
rect 20729 18717 20763 18751
rect 20763 18717 20772 18751
rect 20720 18708 20772 18717
rect 21732 18708 21784 18760
rect 25964 18708 26016 18760
rect 14740 18640 14792 18692
rect 2964 18615 3016 18624
rect 2964 18581 2973 18615
rect 2973 18581 3007 18615
rect 3007 18581 3016 18615
rect 2964 18572 3016 18581
rect 7748 18615 7800 18624
rect 7748 18581 7757 18615
rect 7757 18581 7791 18615
rect 7791 18581 7800 18615
rect 7748 18572 7800 18581
rect 22284 18640 22336 18692
rect 27620 18640 27672 18692
rect 31760 18708 31812 18760
rect 36084 18751 36136 18760
rect 36084 18717 36093 18751
rect 36093 18717 36127 18751
rect 36127 18717 36136 18751
rect 36084 18708 36136 18717
rect 37832 18708 37884 18760
rect 32772 18640 32824 18692
rect 15568 18572 15620 18624
rect 20720 18572 20772 18624
rect 37464 18615 37516 18624
rect 37464 18581 37473 18615
rect 37473 18581 37507 18615
rect 37507 18581 37516 18615
rect 37464 18572 37516 18581
rect 41420 18708 41472 18760
rect 42432 18708 42484 18760
rect 45008 18708 45060 18760
rect 52000 18708 52052 18760
rect 56692 18751 56744 18760
rect 56692 18717 56701 18751
rect 56701 18717 56735 18751
rect 56735 18717 56744 18751
rect 56692 18708 56744 18717
rect 39672 18640 39724 18692
rect 43812 18640 43864 18692
rect 46388 18640 46440 18692
rect 52644 18640 52696 18692
rect 57244 18640 57296 18692
rect 38292 18572 38344 18624
rect 39304 18615 39356 18624
rect 39304 18581 39313 18615
rect 39313 18581 39347 18615
rect 39347 18581 39356 18615
rect 39304 18572 39356 18581
rect 51816 18572 51868 18624
rect 58072 18615 58124 18624
rect 58072 18581 58081 18615
rect 58081 18581 58115 18615
rect 58115 18581 58124 18615
rect 58072 18572 58124 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 2964 18300 3016 18352
rect 12716 18368 12768 18420
rect 14740 18411 14792 18420
rect 14740 18377 14749 18411
rect 14749 18377 14783 18411
rect 14783 18377 14792 18411
rect 14740 18368 14792 18377
rect 19248 18368 19300 18420
rect 21272 18411 21324 18420
rect 21272 18377 21281 18411
rect 21281 18377 21315 18411
rect 21315 18377 21324 18411
rect 21272 18368 21324 18377
rect 28908 18411 28960 18420
rect 28908 18377 28917 18411
rect 28917 18377 28951 18411
rect 28951 18377 28960 18411
rect 28908 18368 28960 18377
rect 31208 18411 31260 18420
rect 31208 18377 31217 18411
rect 31217 18377 31251 18411
rect 31251 18377 31260 18411
rect 31208 18368 31260 18377
rect 36728 18411 36780 18420
rect 36728 18377 36737 18411
rect 36737 18377 36771 18411
rect 36771 18377 36780 18411
rect 36728 18368 36780 18377
rect 39672 18411 39724 18420
rect 39672 18377 39681 18411
rect 39681 18377 39715 18411
rect 39715 18377 39724 18411
rect 39672 18368 39724 18377
rect 43812 18411 43864 18420
rect 43812 18377 43821 18411
rect 43821 18377 43855 18411
rect 43855 18377 43864 18411
rect 43812 18368 43864 18377
rect 46388 18411 46440 18420
rect 46388 18377 46397 18411
rect 46397 18377 46431 18411
rect 46431 18377 46440 18411
rect 46388 18368 46440 18377
rect 7748 18300 7800 18352
rect 14004 18300 14056 18352
rect 20536 18300 20588 18352
rect 23204 18300 23256 18352
rect 25044 18300 25096 18352
rect 28724 18300 28776 18352
rect 33508 18300 33560 18352
rect 34520 18300 34572 18352
rect 1584 18232 1636 18284
rect 4620 18232 4672 18284
rect 6368 18275 6420 18284
rect 6368 18241 6377 18275
rect 6377 18241 6411 18275
rect 6411 18241 6420 18275
rect 6368 18232 6420 18241
rect 8300 18232 8352 18284
rect 9404 18232 9456 18284
rect 11612 18232 11664 18284
rect 12900 18232 12952 18284
rect 14096 18232 14148 18284
rect 21272 18232 21324 18284
rect 21732 18232 21784 18284
rect 23664 18275 23716 18284
rect 23664 18241 23673 18275
rect 23673 18241 23707 18275
rect 23707 18241 23716 18275
rect 23664 18232 23716 18241
rect 27620 18232 27672 18284
rect 29920 18232 29972 18284
rect 36084 18300 36136 18352
rect 38660 18300 38712 18352
rect 40132 18343 40184 18352
rect 40132 18309 40141 18343
rect 40141 18309 40175 18343
rect 40175 18309 40184 18343
rect 40132 18300 40184 18309
rect 17316 18164 17368 18216
rect 4988 18071 5040 18080
rect 4988 18037 4997 18071
rect 4997 18037 5031 18071
rect 5031 18037 5040 18071
rect 4988 18028 5040 18037
rect 9588 18071 9640 18080
rect 9588 18037 9597 18071
rect 9597 18037 9631 18071
rect 9631 18037 9640 18071
rect 9588 18028 9640 18037
rect 32772 18164 32824 18216
rect 37096 18232 37148 18284
rect 38292 18275 38344 18284
rect 38292 18241 38301 18275
rect 38301 18241 38335 18275
rect 38335 18241 38344 18275
rect 38292 18232 38344 18241
rect 41512 18232 41564 18284
rect 43536 18232 43588 18284
rect 45100 18232 45152 18284
rect 46388 18232 46440 18284
rect 51264 18300 51316 18352
rect 52000 18300 52052 18352
rect 58072 18300 58124 18352
rect 52184 18232 52236 18284
rect 54760 18232 54812 18284
rect 56692 18232 56744 18284
rect 53840 18164 53892 18216
rect 23480 18096 23532 18148
rect 20904 18028 20956 18080
rect 25228 18028 25280 18080
rect 36360 18028 36412 18080
rect 50620 18028 50672 18080
rect 54300 18028 54352 18080
rect 55864 18028 55916 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 22284 17867 22336 17876
rect 22284 17833 22293 17867
rect 22293 17833 22327 17867
rect 22327 17833 22336 17867
rect 22284 17824 22336 17833
rect 37096 17824 37148 17876
rect 1584 17688 1636 17740
rect 2504 17688 2556 17740
rect 14096 17731 14148 17740
rect 14096 17697 14105 17731
rect 14105 17697 14139 17731
rect 14139 17697 14148 17731
rect 14096 17688 14148 17697
rect 29920 17688 29972 17740
rect 32772 17731 32824 17740
rect 32772 17697 32781 17731
rect 32781 17697 32815 17731
rect 32815 17697 32824 17731
rect 32772 17688 32824 17697
rect 37372 17688 37424 17740
rect 38292 17824 38344 17876
rect 39120 17824 39172 17876
rect 42432 17824 42484 17876
rect 43536 17867 43588 17876
rect 43536 17833 43545 17867
rect 43545 17833 43579 17867
rect 43579 17833 43588 17867
rect 43536 17824 43588 17833
rect 46388 17867 46440 17876
rect 46388 17833 46397 17867
rect 46397 17833 46431 17867
rect 46431 17833 46440 17867
rect 46388 17824 46440 17833
rect 52644 17867 52696 17876
rect 52644 17833 52653 17867
rect 52653 17833 52687 17867
rect 52687 17833 52696 17867
rect 52644 17824 52696 17833
rect 45008 17731 45060 17740
rect 45008 17697 45017 17731
rect 45017 17697 45051 17731
rect 45051 17697 45060 17731
rect 45008 17688 45060 17697
rect 47216 17688 47268 17740
rect 51264 17731 51316 17740
rect 51264 17697 51273 17731
rect 51273 17697 51307 17731
rect 51307 17697 51316 17731
rect 51264 17688 51316 17697
rect 4528 17620 4580 17672
rect 5448 17620 5500 17672
rect 8944 17663 8996 17672
rect 8944 17629 8953 17663
rect 8953 17629 8987 17663
rect 8987 17629 8996 17663
rect 8944 17620 8996 17629
rect 11612 17620 11664 17672
rect 15568 17620 15620 17672
rect 17316 17620 17368 17672
rect 20904 17663 20956 17672
rect 20904 17629 20913 17663
rect 20913 17629 20947 17663
rect 20947 17629 20956 17663
rect 20904 17620 20956 17629
rect 21732 17620 21784 17672
rect 24400 17620 24452 17672
rect 3884 17552 3936 17604
rect 7748 17552 7800 17604
rect 10232 17552 10284 17604
rect 4620 17484 4672 17536
rect 8392 17484 8444 17536
rect 15844 17552 15896 17604
rect 23204 17552 23256 17604
rect 25228 17620 25280 17672
rect 27620 17663 27672 17672
rect 27620 17629 27629 17663
rect 27629 17629 27663 17663
rect 27663 17629 27672 17663
rect 27620 17620 27672 17629
rect 39304 17620 39356 17672
rect 53840 17824 53892 17876
rect 54300 17620 54352 17672
rect 55956 17620 56008 17672
rect 29736 17552 29788 17604
rect 31576 17552 31628 17604
rect 35348 17552 35400 17604
rect 38844 17552 38896 17604
rect 43812 17552 43864 17604
rect 46296 17552 46348 17604
rect 48780 17552 48832 17604
rect 11336 17484 11388 17536
rect 15476 17527 15528 17536
rect 15476 17493 15485 17527
rect 15485 17493 15519 17527
rect 15519 17493 15528 17527
rect 15476 17484 15528 17493
rect 15752 17484 15804 17536
rect 26516 17527 26568 17536
rect 26516 17493 26525 17527
rect 26525 17493 26559 17527
rect 26559 17493 26568 17527
rect 26516 17484 26568 17493
rect 29000 17527 29052 17536
rect 29000 17493 29009 17527
rect 29009 17493 29043 17527
rect 29043 17493 29052 17527
rect 29000 17484 29052 17493
rect 30472 17484 30524 17536
rect 34796 17484 34848 17536
rect 49056 17527 49108 17536
rect 49056 17493 49065 17527
rect 49065 17493 49099 17527
rect 49099 17493 49108 17527
rect 49056 17484 49108 17493
rect 57336 17552 57388 17604
rect 58164 17527 58216 17536
rect 58164 17493 58173 17527
rect 58173 17493 58207 17527
rect 58207 17493 58216 17527
rect 58164 17484 58216 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 3884 17323 3936 17332
rect 3884 17289 3893 17323
rect 3893 17289 3927 17323
rect 3927 17289 3936 17323
rect 3884 17280 3936 17289
rect 7748 17323 7800 17332
rect 7748 17289 7757 17323
rect 7757 17289 7791 17323
rect 7791 17289 7800 17323
rect 7748 17280 7800 17289
rect 9404 17280 9456 17332
rect 12900 17323 12952 17332
rect 12900 17289 12909 17323
rect 12909 17289 12943 17323
rect 12943 17289 12952 17323
rect 12900 17280 12952 17289
rect 21272 17323 21324 17332
rect 21272 17289 21281 17323
rect 21281 17289 21315 17323
rect 21315 17289 21324 17323
rect 21272 17280 21324 17289
rect 23204 17323 23256 17332
rect 23204 17289 23213 17323
rect 23213 17289 23247 17323
rect 23247 17289 23256 17323
rect 23204 17280 23256 17289
rect 29000 17280 29052 17332
rect 35348 17323 35400 17332
rect 4988 17212 5040 17264
rect 2504 17187 2556 17196
rect 2504 17153 2513 17187
rect 2513 17153 2547 17187
rect 2547 17153 2556 17187
rect 2504 17144 2556 17153
rect 4436 17144 4488 17196
rect 5172 17144 5224 17196
rect 5448 17144 5500 17196
rect 7012 17144 7064 17196
rect 8944 17212 8996 17264
rect 15476 17212 15528 17264
rect 20720 17212 20772 17264
rect 26516 17212 26568 17264
rect 30472 17255 30524 17264
rect 30472 17221 30506 17255
rect 30506 17221 30524 17255
rect 30472 17212 30524 17221
rect 35348 17289 35357 17323
rect 35357 17289 35391 17323
rect 35391 17289 35400 17323
rect 35348 17280 35400 17289
rect 37004 17280 37056 17332
rect 38752 17323 38804 17332
rect 32772 17212 32824 17264
rect 9404 17144 9456 17196
rect 11612 17144 11664 17196
rect 12164 17144 12216 17196
rect 14096 17187 14148 17196
rect 14096 17153 14105 17187
rect 14105 17153 14139 17187
rect 14139 17153 14148 17187
rect 14096 17144 14148 17153
rect 17316 17144 17368 17196
rect 18512 17144 18564 17196
rect 20904 17144 20956 17196
rect 21824 17187 21876 17196
rect 21824 17153 21833 17187
rect 21833 17153 21867 17187
rect 21867 17153 21876 17187
rect 21824 17144 21876 17153
rect 23204 17144 23256 17196
rect 23664 17144 23716 17196
rect 24400 17187 24452 17196
rect 24400 17153 24409 17187
rect 24409 17153 24443 17187
rect 24443 17153 24452 17187
rect 24400 17144 24452 17153
rect 33508 17144 33560 17196
rect 37464 17212 37516 17264
rect 38752 17289 38761 17323
rect 38761 17289 38795 17323
rect 38795 17289 38804 17323
rect 38752 17280 38804 17289
rect 40684 17280 40736 17332
rect 43812 17323 43864 17332
rect 43812 17289 43821 17323
rect 43821 17289 43855 17323
rect 43855 17289 43864 17323
rect 43812 17280 43864 17289
rect 46296 17280 46348 17332
rect 52184 17323 52236 17332
rect 52184 17289 52193 17323
rect 52193 17289 52227 17323
rect 52227 17289 52236 17323
rect 52184 17280 52236 17289
rect 57244 17280 57296 17332
rect 37280 17144 37332 17196
rect 37372 17187 37424 17196
rect 37372 17153 37381 17187
rect 37381 17153 37415 17187
rect 37415 17153 37424 17187
rect 37372 17144 37424 17153
rect 37924 17144 37976 17196
rect 43904 17144 43956 17196
rect 45008 17187 45060 17196
rect 45008 17153 45017 17187
rect 45017 17153 45051 17187
rect 45051 17153 45060 17187
rect 45008 17144 45060 17153
rect 46388 17144 46440 17196
rect 47216 17144 47268 17196
rect 50804 17212 50856 17264
rect 55864 17212 55916 17264
rect 58164 17212 58216 17264
rect 50896 17144 50948 17196
rect 52920 17144 52972 17196
rect 53840 17144 53892 17196
rect 55956 17187 56008 17196
rect 55956 17153 55965 17187
rect 55965 17153 55999 17187
rect 55999 17153 56008 17187
rect 55956 17144 56008 17153
rect 27620 17076 27672 17128
rect 4712 16940 4764 16992
rect 15476 16983 15528 16992
rect 15476 16949 15485 16983
rect 15485 16949 15519 16983
rect 15519 16949 15528 16983
rect 15476 16940 15528 16949
rect 19340 16940 19392 16992
rect 25780 16983 25832 16992
rect 25780 16949 25789 16983
rect 25789 16949 25823 16983
rect 25823 16949 25832 16983
rect 25780 16940 25832 16949
rect 29920 17076 29972 17128
rect 42432 17119 42484 17128
rect 29736 17051 29788 17060
rect 29736 17017 29745 17051
rect 29745 17017 29779 17051
rect 29779 17017 29788 17051
rect 29736 17008 29788 17017
rect 42432 17085 42441 17119
rect 42441 17085 42475 17119
rect 42475 17085 42484 17119
rect 42432 17076 42484 17085
rect 50804 17119 50856 17128
rect 50804 17085 50813 17119
rect 50813 17085 50847 17119
rect 50847 17085 50856 17119
rect 50804 17076 50856 17085
rect 32312 16940 32364 16992
rect 33232 16940 33284 16992
rect 49332 16940 49384 16992
rect 55496 16983 55548 16992
rect 55496 16949 55505 16983
rect 55505 16949 55539 16983
rect 55539 16949 55548 16983
rect 55496 16940 55548 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 5172 16779 5224 16788
rect 5172 16745 5181 16779
rect 5181 16745 5215 16779
rect 5215 16745 5224 16779
rect 5172 16736 5224 16745
rect 7012 16779 7064 16788
rect 7012 16745 7021 16779
rect 7021 16745 7055 16779
rect 7055 16745 7064 16779
rect 7012 16736 7064 16745
rect 9312 16736 9364 16788
rect 10232 16736 10284 16788
rect 12164 16779 12216 16788
rect 12164 16745 12173 16779
rect 12173 16745 12207 16779
rect 12207 16745 12216 16779
rect 12164 16736 12216 16745
rect 15844 16736 15896 16788
rect 18512 16779 18564 16788
rect 18512 16745 18521 16779
rect 18521 16745 18555 16779
rect 18555 16745 18564 16779
rect 18512 16736 18564 16745
rect 37280 16736 37332 16788
rect 43904 16779 43956 16788
rect 43904 16745 43913 16779
rect 43913 16745 43947 16779
rect 43947 16745 43956 16779
rect 43904 16736 43956 16745
rect 46388 16779 46440 16788
rect 46388 16745 46397 16779
rect 46397 16745 46431 16779
rect 46431 16745 46440 16779
rect 46388 16736 46440 16745
rect 48780 16779 48832 16788
rect 48780 16745 48789 16779
rect 48789 16745 48823 16779
rect 48823 16745 48832 16779
rect 48780 16736 48832 16745
rect 52920 16779 52972 16788
rect 52920 16745 52929 16779
rect 52929 16745 52963 16779
rect 52963 16745 52972 16779
rect 52920 16736 52972 16745
rect 14004 16600 14056 16652
rect 24400 16643 24452 16652
rect 24400 16609 24409 16643
rect 24409 16609 24443 16643
rect 24443 16609 24452 16643
rect 24400 16600 24452 16609
rect 36084 16643 36136 16652
rect 36084 16609 36093 16643
rect 36093 16609 36127 16643
rect 36127 16609 36136 16643
rect 36084 16600 36136 16609
rect 37832 16600 37884 16652
rect 39764 16600 39816 16652
rect 42432 16600 42484 16652
rect 47400 16643 47452 16652
rect 2688 16532 2740 16584
rect 4620 16532 4672 16584
rect 5540 16532 5592 16584
rect 9588 16532 9640 16584
rect 10416 16532 10468 16584
rect 11336 16532 11388 16584
rect 15476 16532 15528 16584
rect 16672 16532 16724 16584
rect 19156 16532 19208 16584
rect 20904 16575 20956 16584
rect 20904 16541 20913 16575
rect 20913 16541 20947 16575
rect 20947 16541 20956 16575
rect 20904 16532 20956 16541
rect 25780 16532 25832 16584
rect 26240 16575 26292 16584
rect 26240 16541 26249 16575
rect 26249 16541 26283 16575
rect 26283 16541 26292 16575
rect 26240 16532 26292 16541
rect 31760 16532 31812 16584
rect 36360 16575 36412 16584
rect 36360 16541 36394 16575
rect 36394 16541 36412 16575
rect 45008 16575 45060 16584
rect 36360 16532 36412 16541
rect 45008 16541 45017 16575
rect 45017 16541 45051 16575
rect 45051 16541 45060 16575
rect 47400 16609 47409 16643
rect 47409 16609 47443 16643
rect 47443 16609 47452 16643
rect 47400 16600 47452 16609
rect 45008 16532 45060 16541
rect 49332 16532 49384 16584
rect 51540 16575 51592 16584
rect 51540 16541 51549 16575
rect 51549 16541 51583 16575
rect 51583 16541 51592 16575
rect 51540 16532 51592 16541
rect 51816 16575 51868 16584
rect 51816 16541 51850 16575
rect 51850 16541 51868 16575
rect 51816 16532 51868 16541
rect 7748 16464 7800 16516
rect 9312 16464 9364 16516
rect 19248 16464 19300 16516
rect 23480 16464 23532 16516
rect 25872 16464 25924 16516
rect 31852 16464 31904 16516
rect 39856 16464 39908 16516
rect 42616 16464 42668 16516
rect 43812 16464 43864 16516
rect 46388 16464 46440 16516
rect 55956 16532 56008 16584
rect 55404 16464 55456 16516
rect 57796 16464 57848 16516
rect 22284 16439 22336 16448
rect 22284 16405 22293 16439
rect 22293 16405 22327 16439
rect 22327 16405 22336 16439
rect 22284 16396 22336 16405
rect 25780 16439 25832 16448
rect 25780 16405 25789 16439
rect 25789 16405 25823 16439
rect 25823 16405 25832 16439
rect 25780 16396 25832 16405
rect 27068 16396 27120 16448
rect 32220 16396 32272 16448
rect 39948 16396 40000 16448
rect 42064 16439 42116 16448
rect 42064 16405 42073 16439
rect 42073 16405 42107 16439
rect 42107 16405 42116 16439
rect 42064 16396 42116 16405
rect 54760 16439 54812 16448
rect 54760 16405 54769 16439
rect 54769 16405 54803 16439
rect 54803 16405 54812 16439
rect 54760 16396 54812 16405
rect 57888 16439 57940 16448
rect 57888 16405 57897 16439
rect 57897 16405 57931 16439
rect 57931 16405 57940 16439
rect 57888 16396 57940 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 7748 16235 7800 16244
rect 7748 16201 7757 16235
rect 7757 16201 7791 16235
rect 7791 16201 7800 16235
rect 7748 16192 7800 16201
rect 8392 16192 8444 16244
rect 4712 16124 4764 16176
rect 9404 16192 9456 16244
rect 19340 16192 19392 16244
rect 20536 16235 20588 16244
rect 2688 15988 2740 16040
rect 1768 15852 1820 15904
rect 5540 15988 5592 16040
rect 6920 16056 6972 16108
rect 15752 16124 15804 16176
rect 20536 16201 20545 16235
rect 20545 16201 20579 16235
rect 20579 16201 20588 16235
rect 20536 16192 20588 16201
rect 23204 16235 23256 16244
rect 23204 16201 23213 16235
rect 23213 16201 23247 16235
rect 23247 16201 23256 16235
rect 23204 16192 23256 16201
rect 22284 16124 22336 16176
rect 26240 16192 26292 16244
rect 26792 16192 26844 16244
rect 31576 16235 31628 16244
rect 31576 16201 31585 16235
rect 31585 16201 31619 16235
rect 31619 16201 31628 16235
rect 31576 16192 31628 16201
rect 32312 16192 32364 16244
rect 33508 16235 33560 16244
rect 25780 16124 25832 16176
rect 32220 16124 32272 16176
rect 33508 16201 33517 16235
rect 33517 16201 33551 16235
rect 33551 16201 33560 16235
rect 33508 16192 33560 16201
rect 43812 16235 43864 16244
rect 43812 16201 43821 16235
rect 43821 16201 43855 16235
rect 43855 16201 43864 16235
rect 43812 16192 43864 16201
rect 46388 16235 46440 16244
rect 46388 16201 46397 16235
rect 46397 16201 46431 16235
rect 46431 16201 46440 16235
rect 46388 16192 46440 16201
rect 50896 16192 50948 16244
rect 57336 16235 57388 16244
rect 57336 16201 57345 16235
rect 57345 16201 57379 16235
rect 57379 16201 57388 16235
rect 57336 16192 57388 16201
rect 34796 16124 34848 16176
rect 14280 16056 14332 16108
rect 16672 16056 16724 16108
rect 17316 16099 17368 16108
rect 17316 16065 17325 16099
rect 17325 16065 17359 16099
rect 17359 16065 17368 16099
rect 17316 16056 17368 16065
rect 18696 16056 18748 16108
rect 19156 16099 19208 16108
rect 19156 16065 19165 16099
rect 19165 16065 19199 16099
rect 19199 16065 19208 16099
rect 19156 16056 19208 16065
rect 24400 16099 24452 16108
rect 24400 16065 24409 16099
rect 24409 16065 24443 16099
rect 24443 16065 24452 16099
rect 24400 16056 24452 16065
rect 26332 16056 26384 16108
rect 31760 16056 31812 16108
rect 32864 16056 32916 16108
rect 20904 15988 20956 16040
rect 26792 15988 26844 16040
rect 34704 16031 34756 16040
rect 34704 15997 34713 16031
rect 34713 15997 34747 16031
rect 34747 15997 34756 16031
rect 34704 15988 34756 15997
rect 37832 16031 37884 16040
rect 37832 15997 37841 16031
rect 37841 15997 37875 16031
rect 37875 15997 37884 16031
rect 39764 16124 39816 16176
rect 39028 16056 39080 16108
rect 37832 15988 37884 15997
rect 40040 15988 40092 16040
rect 41236 16056 41288 16108
rect 42064 16124 42116 16176
rect 49056 16124 49108 16176
rect 50620 16167 50672 16176
rect 50620 16133 50654 16167
rect 50654 16133 50672 16167
rect 50620 16124 50672 16133
rect 55496 16124 55548 16176
rect 57888 16124 57940 16176
rect 42432 16099 42484 16108
rect 42432 16065 42441 16099
rect 42441 16065 42475 16099
rect 42475 16065 42484 16099
rect 42432 16056 42484 16065
rect 45008 16099 45060 16108
rect 45008 16065 45017 16099
rect 45017 16065 45051 16099
rect 45051 16065 45060 16099
rect 45008 16056 45060 16065
rect 46388 16056 46440 16108
rect 51540 16056 51592 16108
rect 52000 16056 52052 16108
rect 47584 15988 47636 16040
rect 55956 16031 56008 16040
rect 2872 15895 2924 15904
rect 2872 15861 2881 15895
rect 2881 15861 2915 15895
rect 2915 15861 2924 15895
rect 2872 15852 2924 15861
rect 15752 15895 15804 15904
rect 15752 15861 15761 15895
rect 15761 15861 15795 15895
rect 15795 15861 15804 15895
rect 15752 15852 15804 15861
rect 19340 15852 19392 15904
rect 25780 15895 25832 15904
rect 25780 15861 25789 15895
rect 25789 15861 25823 15895
rect 25823 15861 25832 15895
rect 25780 15852 25832 15861
rect 28356 15895 28408 15904
rect 28356 15861 28365 15895
rect 28365 15861 28399 15895
rect 28399 15861 28408 15895
rect 28356 15852 28408 15861
rect 36084 15895 36136 15904
rect 36084 15861 36093 15895
rect 36093 15861 36127 15895
rect 36127 15861 36136 15895
rect 36084 15852 36136 15861
rect 39212 15895 39264 15904
rect 39212 15861 39221 15895
rect 39221 15861 39255 15895
rect 39255 15861 39264 15895
rect 39212 15852 39264 15861
rect 41512 15895 41564 15904
rect 41512 15861 41521 15895
rect 41521 15861 41555 15895
rect 41555 15861 41564 15895
rect 41512 15852 41564 15861
rect 49056 15895 49108 15904
rect 49056 15861 49065 15895
rect 49065 15861 49099 15895
rect 49099 15861 49108 15895
rect 49056 15852 49108 15861
rect 55956 15997 55965 16031
rect 55965 15997 55999 16031
rect 55999 15997 56008 16031
rect 55956 15988 56008 15997
rect 55404 15920 55456 15972
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 6920 15691 6972 15700
rect 6920 15657 6929 15691
rect 6929 15657 6963 15691
rect 6963 15657 6972 15691
rect 18696 15691 18748 15700
rect 6920 15648 6972 15657
rect 18696 15657 18705 15691
rect 18705 15657 18739 15691
rect 18739 15657 18748 15691
rect 18696 15648 18748 15657
rect 20904 15648 20956 15700
rect 23480 15691 23532 15700
rect 14004 15512 14056 15564
rect 23480 15657 23489 15691
rect 23489 15657 23523 15691
rect 23523 15657 23532 15691
rect 23480 15648 23532 15657
rect 25872 15648 25924 15700
rect 39028 15691 39080 15700
rect 39028 15657 39037 15691
rect 39037 15657 39071 15691
rect 39071 15657 39080 15691
rect 39028 15648 39080 15657
rect 41236 15691 41288 15700
rect 41236 15657 41245 15691
rect 41245 15657 41279 15691
rect 41279 15657 41288 15691
rect 41236 15648 41288 15657
rect 42616 15648 42668 15700
rect 46388 15691 46440 15700
rect 46388 15657 46397 15691
rect 46397 15657 46431 15691
rect 46431 15657 46440 15691
rect 46388 15648 46440 15657
rect 57796 15691 57848 15700
rect 57796 15657 57805 15691
rect 57805 15657 57839 15691
rect 57839 15657 57848 15691
rect 57796 15648 57848 15657
rect 24400 15555 24452 15564
rect 24400 15521 24409 15555
rect 24409 15521 24443 15555
rect 24443 15521 24452 15555
rect 24400 15512 24452 15521
rect 39764 15512 39816 15564
rect 1768 15444 1820 15496
rect 2872 15444 2924 15496
rect 5540 15487 5592 15496
rect 5540 15453 5549 15487
rect 5549 15453 5583 15487
rect 5583 15453 5592 15487
rect 5540 15444 5592 15453
rect 9772 15444 9824 15496
rect 10416 15487 10468 15496
rect 10416 15453 10425 15487
rect 10425 15453 10459 15487
rect 10459 15453 10468 15487
rect 10416 15444 10468 15453
rect 15752 15444 15804 15496
rect 17316 15487 17368 15496
rect 17316 15453 17325 15487
rect 17325 15453 17359 15487
rect 17359 15453 17368 15487
rect 17316 15444 17368 15453
rect 25780 15444 25832 15496
rect 26792 15487 26844 15496
rect 26792 15453 26801 15487
rect 26801 15453 26835 15487
rect 26835 15453 26844 15487
rect 26792 15444 26844 15453
rect 28356 15444 28408 15496
rect 32864 15444 32916 15496
rect 34612 15444 34664 15496
rect 36084 15444 36136 15496
rect 37740 15444 37792 15496
rect 39948 15444 40000 15496
rect 45008 15487 45060 15496
rect 45008 15453 45017 15487
rect 45017 15453 45051 15487
rect 45051 15453 45060 15487
rect 45008 15444 45060 15453
rect 48136 15512 48188 15564
rect 7932 15376 7984 15428
rect 12164 15376 12216 15428
rect 18788 15376 18840 15428
rect 19432 15376 19484 15428
rect 23664 15376 23716 15428
rect 3240 15351 3292 15360
rect 3240 15317 3249 15351
rect 3249 15317 3283 15351
rect 3283 15317 3292 15351
rect 3240 15308 3292 15317
rect 11796 15351 11848 15360
rect 11796 15317 11805 15351
rect 11805 15317 11839 15351
rect 11839 15317 11848 15351
rect 11796 15308 11848 15317
rect 15752 15351 15804 15360
rect 15752 15317 15761 15351
rect 15761 15317 15795 15351
rect 15795 15317 15804 15351
rect 15752 15308 15804 15317
rect 28172 15351 28224 15360
rect 28172 15317 28181 15351
rect 28181 15317 28215 15351
rect 28215 15317 28224 15351
rect 28172 15308 28224 15317
rect 32128 15351 32180 15360
rect 32128 15317 32137 15351
rect 32137 15317 32171 15351
rect 32171 15317 32180 15351
rect 32128 15308 32180 15317
rect 33968 15376 34020 15428
rect 38936 15376 38988 15428
rect 41604 15376 41656 15428
rect 46388 15376 46440 15428
rect 52000 15487 52052 15496
rect 51448 15376 51500 15428
rect 52000 15453 52009 15487
rect 52009 15453 52043 15487
rect 52043 15453 52052 15487
rect 52000 15444 52052 15453
rect 55956 15444 56008 15496
rect 56416 15487 56468 15496
rect 56416 15453 56425 15487
rect 56425 15453 56459 15487
rect 56459 15453 56468 15487
rect 56416 15444 56468 15453
rect 33692 15308 33744 15360
rect 34152 15351 34204 15360
rect 34152 15317 34161 15351
rect 34161 15317 34195 15351
rect 34195 15317 34204 15351
rect 34152 15308 34204 15317
rect 36084 15351 36136 15360
rect 36084 15317 36093 15351
rect 36093 15317 36127 15351
rect 36127 15317 36136 15351
rect 36084 15308 36136 15317
rect 47584 15308 47636 15360
rect 49516 15308 49568 15360
rect 52092 15308 52144 15360
rect 53288 15376 53340 15428
rect 57336 15376 57388 15428
rect 53104 15308 53156 15360
rect 53748 15308 53800 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 7932 15147 7984 15156
rect 7932 15113 7941 15147
rect 7941 15113 7975 15147
rect 7975 15113 7984 15147
rect 7932 15104 7984 15113
rect 18788 15147 18840 15156
rect 18788 15113 18797 15147
rect 18797 15113 18831 15147
rect 18831 15113 18840 15147
rect 18788 15104 18840 15113
rect 19248 15104 19300 15156
rect 26332 15147 26384 15156
rect 26332 15113 26341 15147
rect 26341 15113 26375 15147
rect 26375 15113 26384 15147
rect 26332 15104 26384 15113
rect 38936 15147 38988 15156
rect 38936 15113 38945 15147
rect 38945 15113 38979 15147
rect 38979 15113 38988 15147
rect 38936 15104 38988 15113
rect 39856 15104 39908 15156
rect 46388 15147 46440 15156
rect 46388 15113 46397 15147
rect 46397 15113 46431 15147
rect 46431 15113 46440 15147
rect 46388 15104 46440 15113
rect 57336 15147 57388 15156
rect 57336 15113 57345 15147
rect 57345 15113 57379 15147
rect 57379 15113 57388 15147
rect 57336 15104 57388 15113
rect 3240 15036 3292 15088
rect 1768 14968 1820 15020
rect 8116 14968 8168 15020
rect 9772 15036 9824 15088
rect 10968 14968 11020 15020
rect 14280 15011 14332 15020
rect 14280 14977 14289 15011
rect 14289 14977 14323 15011
rect 14323 14977 14332 15011
rect 14280 14968 14332 14977
rect 15752 15036 15804 15088
rect 15384 14968 15436 15020
rect 18512 14968 18564 15020
rect 19156 14968 19208 15020
rect 19340 14968 19392 15020
rect 24400 14968 24452 15020
rect 6276 14900 6328 14952
rect 12256 14943 12308 14952
rect 12256 14909 12265 14943
rect 12265 14909 12299 14943
rect 12299 14909 12308 14943
rect 12256 14900 12308 14909
rect 16672 14900 16724 14952
rect 17316 14900 17368 14952
rect 27068 15036 27120 15088
rect 28172 15036 28224 15088
rect 33232 15036 33284 15088
rect 36084 15036 36136 15088
rect 37740 15036 37792 15088
rect 39212 15036 39264 15088
rect 26792 14968 26844 15020
rect 34520 14968 34572 15020
rect 34612 14968 34664 15020
rect 37556 15011 37608 15020
rect 37556 14977 37565 15011
rect 37565 14977 37599 15011
rect 37599 14977 37608 15011
rect 37556 14968 37608 14977
rect 38936 14968 38988 15020
rect 40040 14968 40092 15020
rect 45560 15036 45612 15088
rect 49056 15036 49108 15088
rect 46664 14968 46716 15020
rect 49148 14968 49200 15020
rect 52000 14968 52052 15020
rect 54852 14968 54904 15020
rect 57336 14968 57388 15020
rect 28816 14943 28868 14952
rect 3056 14807 3108 14816
rect 3056 14773 3065 14807
rect 3065 14773 3099 14807
rect 3099 14773 3108 14807
rect 3056 14764 3108 14773
rect 9680 14764 9732 14816
rect 13636 14807 13688 14816
rect 13636 14773 13645 14807
rect 13645 14773 13679 14807
rect 13679 14773 13688 14807
rect 13636 14764 13688 14773
rect 15660 14807 15712 14816
rect 15660 14773 15669 14807
rect 15669 14773 15703 14807
rect 15703 14773 15712 14807
rect 15660 14764 15712 14773
rect 24492 14807 24544 14816
rect 24492 14773 24501 14807
rect 24501 14773 24535 14807
rect 24535 14773 24544 14807
rect 24492 14764 24544 14773
rect 28816 14909 28825 14943
rect 28825 14909 28859 14943
rect 28859 14909 28868 14943
rect 28816 14900 28868 14909
rect 32864 14943 32916 14952
rect 32864 14909 32873 14943
rect 32873 14909 32907 14943
rect 32907 14909 32916 14943
rect 32864 14900 32916 14909
rect 47584 14900 47636 14952
rect 49516 14943 49568 14952
rect 49516 14909 49525 14943
rect 49525 14909 49559 14943
rect 49559 14909 49568 14943
rect 49516 14900 49568 14909
rect 54944 14900 54996 14952
rect 26700 14764 26752 14816
rect 28356 14807 28408 14816
rect 28356 14773 28365 14807
rect 28365 14773 28399 14807
rect 28399 14773 28408 14807
rect 28356 14764 28408 14773
rect 30196 14807 30248 14816
rect 30196 14773 30205 14807
rect 30205 14773 30239 14807
rect 30239 14773 30248 14807
rect 30196 14764 30248 14773
rect 34704 14764 34756 14816
rect 36084 14807 36136 14816
rect 36084 14773 36093 14807
rect 36093 14773 36127 14807
rect 36127 14773 36136 14807
rect 36084 14764 36136 14773
rect 49056 14807 49108 14816
rect 49056 14773 49065 14807
rect 49065 14773 49099 14807
rect 49099 14773 49108 14807
rect 49056 14764 49108 14773
rect 49792 14764 49844 14816
rect 53656 14764 53708 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 8116 14603 8168 14612
rect 8116 14569 8125 14603
rect 8125 14569 8159 14603
rect 8159 14569 8168 14603
rect 8116 14560 8168 14569
rect 18512 14603 18564 14612
rect 18512 14569 18521 14603
rect 18521 14569 18555 14603
rect 18555 14569 18564 14603
rect 18512 14560 18564 14569
rect 23664 14603 23716 14612
rect 23664 14569 23673 14603
rect 23673 14569 23707 14603
rect 23707 14569 23716 14603
rect 23664 14560 23716 14569
rect 31852 14603 31904 14612
rect 31852 14569 31861 14603
rect 31861 14569 31895 14603
rect 31895 14569 31904 14603
rect 31852 14560 31904 14569
rect 41604 14560 41656 14612
rect 46664 14603 46716 14612
rect 46664 14569 46673 14603
rect 46673 14569 46707 14603
rect 46707 14569 46716 14603
rect 46664 14560 46716 14569
rect 19156 14424 19208 14476
rect 32864 14424 32916 14476
rect 34612 14424 34664 14476
rect 34796 14424 34848 14476
rect 39764 14424 39816 14476
rect 45008 14424 45060 14476
rect 52000 14467 52052 14476
rect 52000 14433 52009 14467
rect 52009 14433 52043 14467
rect 52043 14433 52052 14467
rect 52000 14424 52052 14433
rect 1768 14356 1820 14408
rect 3056 14356 3108 14408
rect 6276 14356 6328 14408
rect 11060 14356 11112 14408
rect 7932 14288 7984 14340
rect 3056 14263 3108 14272
rect 3056 14229 3065 14263
rect 3065 14229 3099 14263
rect 3099 14229 3108 14263
rect 3056 14220 3108 14229
rect 5540 14220 5592 14272
rect 10784 14220 10836 14272
rect 12256 14356 12308 14408
rect 14188 14356 14240 14408
rect 15660 14356 15712 14408
rect 16764 14356 16816 14408
rect 14556 14288 14608 14340
rect 21272 14288 21324 14340
rect 24400 14356 24452 14408
rect 28816 14356 28868 14408
rect 22376 14288 22428 14340
rect 23204 14288 23256 14340
rect 26240 14288 26292 14340
rect 27528 14331 27580 14340
rect 27528 14297 27537 14331
rect 27537 14297 27571 14331
rect 27571 14297 27580 14331
rect 27528 14288 27580 14297
rect 14188 14220 14240 14272
rect 15476 14263 15528 14272
rect 15476 14229 15485 14263
rect 15485 14229 15519 14263
rect 15519 14229 15528 14263
rect 15476 14220 15528 14229
rect 21824 14263 21876 14272
rect 21824 14229 21833 14263
rect 21833 14229 21867 14263
rect 21867 14229 21876 14263
rect 21824 14220 21876 14229
rect 32128 14356 32180 14408
rect 36084 14356 36136 14408
rect 41512 14356 41564 14408
rect 47584 14399 47636 14408
rect 47584 14365 47593 14399
rect 47593 14365 47627 14399
rect 47627 14365 47636 14399
rect 47584 14356 47636 14365
rect 49056 14356 49108 14408
rect 52092 14356 52144 14408
rect 55956 14356 56008 14408
rect 56416 14356 56468 14408
rect 32312 14331 32364 14340
rect 32312 14297 32321 14331
rect 32321 14297 32355 14331
rect 32355 14297 32364 14331
rect 32312 14288 32364 14297
rect 39856 14288 39908 14340
rect 46388 14288 46440 14340
rect 49700 14288 49752 14340
rect 55588 14288 55640 14340
rect 32864 14220 32916 14272
rect 36268 14263 36320 14272
rect 36268 14229 36277 14263
rect 36277 14229 36311 14263
rect 36311 14229 36320 14263
rect 36268 14220 36320 14229
rect 48964 14263 49016 14272
rect 48964 14229 48973 14263
rect 48973 14229 49007 14263
rect 49007 14229 49016 14263
rect 48964 14220 49016 14229
rect 51540 14263 51592 14272
rect 51540 14229 51549 14263
rect 51549 14229 51583 14263
rect 51583 14229 51592 14263
rect 51540 14220 51592 14229
rect 53380 14263 53432 14272
rect 53380 14229 53389 14263
rect 53389 14229 53423 14263
rect 53423 14229 53432 14263
rect 53380 14220 53432 14229
rect 58072 14263 58124 14272
rect 58072 14229 58081 14263
rect 58081 14229 58115 14263
rect 58115 14229 58124 14263
rect 58072 14220 58124 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 7932 14059 7984 14068
rect 7932 14025 7941 14059
rect 7941 14025 7975 14059
rect 7975 14025 7984 14059
rect 7932 14016 7984 14025
rect 23204 14059 23256 14068
rect 3056 13948 3108 14000
rect 15476 13948 15528 14000
rect 1768 13880 1820 13932
rect 8208 13880 8260 13932
rect 13636 13880 13688 13932
rect 14096 13923 14148 13932
rect 14096 13889 14105 13923
rect 14105 13889 14139 13923
rect 14139 13889 14148 13923
rect 14096 13880 14148 13889
rect 16764 13880 16816 13932
rect 21824 13948 21876 14000
rect 23204 14025 23213 14059
rect 23213 14025 23247 14059
rect 23247 14025 23256 14059
rect 23204 14016 23256 14025
rect 22192 13948 22244 14000
rect 30196 14016 30248 14068
rect 33968 14016 34020 14068
rect 38936 14059 38988 14068
rect 38936 14025 38945 14059
rect 38945 14025 38979 14059
rect 38979 14025 38988 14059
rect 38936 14016 38988 14025
rect 44548 14016 44600 14068
rect 49148 14016 49200 14068
rect 28356 13948 28408 14000
rect 6276 13812 6328 13864
rect 3056 13719 3108 13728
rect 3056 13685 3065 13719
rect 3065 13685 3099 13719
rect 3099 13685 3108 13719
rect 3056 13676 3108 13685
rect 10784 13812 10836 13864
rect 24400 13880 24452 13932
rect 27068 13880 27120 13932
rect 27528 13880 27580 13932
rect 29092 13923 29144 13932
rect 29092 13889 29126 13923
rect 29126 13889 29144 13923
rect 29092 13880 29144 13889
rect 32864 13880 32916 13932
rect 34796 13880 34848 13932
rect 36268 13948 36320 14000
rect 36084 13880 36136 13932
rect 37556 13923 37608 13932
rect 37556 13889 37565 13923
rect 37565 13889 37599 13923
rect 37599 13889 37608 13923
rect 37556 13880 37608 13889
rect 38936 13880 38988 13932
rect 18236 13812 18288 13864
rect 19156 13812 19208 13864
rect 42984 13880 43036 13932
rect 44916 13948 44968 14000
rect 48964 13948 49016 14000
rect 51540 13948 51592 14000
rect 54944 13948 54996 14000
rect 46756 13880 46808 13932
rect 49516 13880 49568 13932
rect 53104 13923 53156 13932
rect 53104 13889 53113 13923
rect 53113 13889 53147 13923
rect 53147 13889 53156 13923
rect 56692 14016 56744 14068
rect 57336 14059 57388 14068
rect 57336 14025 57345 14059
rect 57345 14025 57379 14059
rect 57379 14025 57388 14059
rect 57336 14016 57388 14025
rect 58072 13948 58124 14000
rect 53104 13880 53156 13889
rect 9772 13676 9824 13728
rect 11060 13676 11112 13728
rect 15476 13719 15528 13728
rect 15476 13685 15485 13719
rect 15485 13685 15519 13719
rect 15519 13685 15528 13719
rect 15476 13676 15528 13685
rect 47584 13812 47636 13864
rect 55956 13855 56008 13864
rect 20812 13676 20864 13728
rect 26424 13719 26476 13728
rect 26424 13685 26433 13719
rect 26433 13685 26467 13719
rect 26467 13685 26476 13719
rect 26424 13676 26476 13685
rect 28356 13719 28408 13728
rect 28356 13685 28365 13719
rect 28365 13685 28399 13719
rect 28399 13685 28408 13719
rect 28356 13676 28408 13685
rect 30196 13719 30248 13728
rect 30196 13685 30205 13719
rect 30205 13685 30239 13719
rect 30239 13685 30248 13719
rect 30196 13676 30248 13685
rect 36360 13719 36412 13728
rect 36360 13685 36369 13719
rect 36369 13685 36403 13719
rect 36403 13685 36412 13719
rect 36360 13676 36412 13685
rect 44272 13719 44324 13728
rect 44272 13685 44281 13719
rect 44281 13685 44315 13719
rect 44315 13685 44324 13719
rect 44272 13676 44324 13685
rect 55956 13821 55965 13855
rect 55965 13821 55999 13855
rect 55999 13821 56008 13855
rect 55956 13812 56008 13821
rect 47952 13676 48004 13728
rect 51172 13719 51224 13728
rect 51172 13685 51181 13719
rect 51181 13685 51215 13719
rect 51215 13685 51224 13719
rect 51172 13676 51224 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 8208 13515 8260 13524
rect 8208 13481 8217 13515
rect 8217 13481 8251 13515
rect 8251 13481 8260 13515
rect 8208 13472 8260 13481
rect 12164 13515 12216 13524
rect 12164 13481 12173 13515
rect 12173 13481 12207 13515
rect 12207 13481 12216 13515
rect 12164 13472 12216 13481
rect 26700 13515 26752 13524
rect 26700 13481 26709 13515
rect 26709 13481 26743 13515
rect 26743 13481 26752 13515
rect 26700 13472 26752 13481
rect 34520 13472 34572 13524
rect 38936 13515 38988 13524
rect 38936 13481 38945 13515
rect 38945 13481 38979 13515
rect 38979 13481 38988 13515
rect 38936 13472 38988 13481
rect 42984 13472 43036 13524
rect 46388 13515 46440 13524
rect 46388 13481 46397 13515
rect 46397 13481 46431 13515
rect 46431 13481 46440 13515
rect 46388 13472 46440 13481
rect 49700 13472 49752 13524
rect 51448 13472 51500 13524
rect 53288 13472 53340 13524
rect 24400 13336 24452 13388
rect 27068 13336 27120 13388
rect 34796 13336 34848 13388
rect 37556 13379 37608 13388
rect 1860 13311 1912 13320
rect 1860 13277 1869 13311
rect 1869 13277 1903 13311
rect 1903 13277 1912 13311
rect 1860 13268 1912 13277
rect 3056 13268 3108 13320
rect 5540 13268 5592 13320
rect 6276 13268 6328 13320
rect 9772 13268 9824 13320
rect 10784 13311 10836 13320
rect 10784 13277 10793 13311
rect 10793 13277 10827 13311
rect 10827 13277 10836 13311
rect 10784 13268 10836 13277
rect 11060 13311 11112 13320
rect 11060 13277 11094 13311
rect 11094 13277 11112 13311
rect 11060 13268 11112 13277
rect 20812 13268 20864 13320
rect 26424 13268 26476 13320
rect 28356 13268 28408 13320
rect 32864 13268 32916 13320
rect 5816 13200 5868 13252
rect 7748 13200 7800 13252
rect 11796 13200 11848 13252
rect 15292 13200 15344 13252
rect 22284 13200 22336 13252
rect 31944 13200 31996 13252
rect 33784 13200 33836 13252
rect 37556 13345 37565 13379
rect 37565 13345 37599 13379
rect 37599 13345 37608 13379
rect 37556 13336 37608 13345
rect 52000 13379 52052 13388
rect 52000 13345 52009 13379
rect 52009 13345 52043 13379
rect 52043 13345 52052 13379
rect 52000 13336 52052 13345
rect 36360 13268 36412 13320
rect 42524 13268 42576 13320
rect 45560 13268 45612 13320
rect 47952 13311 48004 13320
rect 47952 13277 47961 13311
rect 47961 13277 47995 13311
rect 47995 13277 48004 13311
rect 47952 13268 48004 13277
rect 49792 13268 49844 13320
rect 37556 13200 37608 13252
rect 38844 13200 38896 13252
rect 43904 13200 43956 13252
rect 45744 13200 45796 13252
rect 51172 13268 51224 13320
rect 53380 13268 53432 13320
rect 56692 13311 56744 13320
rect 56692 13277 56701 13311
rect 56701 13277 56735 13311
rect 56735 13277 56744 13311
rect 56692 13268 56744 13277
rect 3240 13175 3292 13184
rect 3240 13141 3249 13175
rect 3249 13141 3283 13175
rect 3283 13141 3292 13175
rect 3240 13132 3292 13141
rect 6368 13175 6420 13184
rect 6368 13141 6377 13175
rect 6377 13141 6411 13175
rect 6411 13141 6420 13175
rect 6368 13132 6420 13141
rect 10324 13175 10376 13184
rect 10324 13141 10333 13175
rect 10333 13141 10367 13175
rect 10367 13141 10376 13175
rect 10324 13132 10376 13141
rect 16672 13132 16724 13184
rect 22100 13175 22152 13184
rect 22100 13141 22109 13175
rect 22109 13141 22143 13175
rect 22143 13141 22152 13175
rect 22100 13132 22152 13141
rect 28540 13175 28592 13184
rect 28540 13141 28549 13175
rect 28549 13141 28583 13175
rect 28583 13141 28592 13175
rect 28540 13132 28592 13141
rect 32404 13132 32456 13184
rect 34244 13132 34296 13184
rect 51172 13132 51224 13184
rect 57244 13132 57296 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 7748 12971 7800 12980
rect 3240 12860 3292 12912
rect 7748 12937 7757 12971
rect 7757 12937 7791 12971
rect 7791 12937 7800 12971
rect 7748 12928 7800 12937
rect 9772 12928 9824 12980
rect 10968 12971 11020 12980
rect 10968 12937 10977 12971
rect 10977 12937 11011 12971
rect 11011 12937 11020 12971
rect 10968 12928 11020 12937
rect 14556 12928 14608 12980
rect 21272 12971 21324 12980
rect 21272 12937 21281 12971
rect 21281 12937 21315 12971
rect 21315 12937 21324 12971
rect 21272 12928 21324 12937
rect 36084 12971 36136 12980
rect 36084 12937 36093 12971
rect 36093 12937 36127 12971
rect 36127 12937 36136 12971
rect 36084 12928 36136 12937
rect 38844 12928 38896 12980
rect 46756 12971 46808 12980
rect 46756 12937 46765 12971
rect 46765 12937 46799 12971
rect 46799 12937 46808 12971
rect 46756 12928 46808 12937
rect 54852 12971 54904 12980
rect 1860 12792 1912 12844
rect 7748 12792 7800 12844
rect 10324 12860 10376 12912
rect 15476 12860 15528 12912
rect 22100 12860 22152 12912
rect 24492 12860 24544 12912
rect 28540 12860 28592 12912
rect 32864 12860 32916 12912
rect 34704 12860 34756 12912
rect 44916 12903 44968 12912
rect 44916 12869 44925 12903
rect 44925 12869 44959 12903
rect 44959 12869 44968 12903
rect 44916 12860 44968 12869
rect 16764 12792 16816 12844
rect 17960 12792 18012 12844
rect 20720 12792 20772 12844
rect 24400 12792 24452 12844
rect 27344 12792 27396 12844
rect 29000 12792 29052 12844
rect 32128 12835 32180 12844
rect 32128 12801 32137 12835
rect 32137 12801 32171 12835
rect 32171 12801 32180 12835
rect 32128 12792 32180 12801
rect 33416 12792 33468 12844
rect 3884 12724 3936 12776
rect 5632 12724 5684 12776
rect 6276 12724 6328 12776
rect 13820 12767 13872 12776
rect 13820 12733 13829 12767
rect 13829 12733 13863 12767
rect 13863 12733 13872 12767
rect 13820 12724 13872 12733
rect 34796 12792 34848 12844
rect 37556 12835 37608 12844
rect 37556 12801 37565 12835
rect 37565 12801 37599 12835
rect 37599 12801 37608 12835
rect 37556 12792 37608 12801
rect 38936 12792 38988 12844
rect 43168 12835 43220 12844
rect 43168 12801 43177 12835
rect 43177 12801 43211 12835
rect 43211 12801 43220 12835
rect 43168 12792 43220 12801
rect 54852 12937 54861 12971
rect 54861 12937 54895 12971
rect 54895 12937 54904 12971
rect 54852 12928 54904 12937
rect 53748 12903 53800 12912
rect 53748 12869 53782 12903
rect 53782 12869 53800 12903
rect 53748 12860 53800 12869
rect 45652 12835 45704 12844
rect 45652 12801 45686 12835
rect 45686 12801 45704 12835
rect 45652 12792 45704 12801
rect 48228 12792 48280 12844
rect 50620 12792 50672 12844
rect 52000 12792 52052 12844
rect 52368 12792 52420 12844
rect 55496 12792 55548 12844
rect 5356 12631 5408 12640
rect 5356 12597 5365 12631
rect 5365 12597 5399 12631
rect 5399 12597 5408 12631
rect 5356 12588 5408 12597
rect 18144 12588 18196 12640
rect 25136 12631 25188 12640
rect 25136 12597 25145 12631
rect 25145 12597 25179 12631
rect 25179 12597 25188 12631
rect 25136 12588 25188 12597
rect 28632 12631 28684 12640
rect 28632 12597 28641 12631
rect 28641 12597 28675 12631
rect 28675 12597 28684 12631
rect 28632 12588 28684 12597
rect 29276 12588 29328 12640
rect 29368 12588 29420 12640
rect 33508 12631 33560 12640
rect 33508 12597 33517 12631
rect 33517 12597 33551 12631
rect 33551 12597 33560 12631
rect 33508 12588 33560 12597
rect 50068 12631 50120 12640
rect 50068 12597 50077 12631
rect 50077 12597 50111 12631
rect 50111 12597 50120 12631
rect 50068 12588 50120 12597
rect 55404 12724 55456 12776
rect 55956 12767 56008 12776
rect 55956 12733 55965 12767
rect 55965 12733 55999 12767
rect 55999 12733 56008 12767
rect 55956 12724 56008 12733
rect 51172 12588 51224 12640
rect 56600 12588 56652 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 5632 12291 5684 12300
rect 5632 12257 5641 12291
rect 5641 12257 5675 12291
rect 5675 12257 5684 12291
rect 5632 12248 5684 12257
rect 9772 12384 9824 12436
rect 11152 12384 11204 12436
rect 15292 12384 15344 12436
rect 15384 12384 15436 12436
rect 22284 12427 22336 12436
rect 22284 12393 22293 12427
rect 22293 12393 22327 12427
rect 22327 12393 22336 12427
rect 22284 12384 22336 12393
rect 29000 12384 29052 12436
rect 38936 12427 38988 12436
rect 38936 12393 38945 12427
rect 38945 12393 38979 12427
rect 38979 12393 38988 12427
rect 38936 12384 38988 12393
rect 39856 12384 39908 12436
rect 41696 12384 41748 12436
rect 43168 12384 43220 12436
rect 43904 12427 43956 12436
rect 43904 12393 43913 12427
rect 43913 12393 43947 12427
rect 43947 12393 43956 12427
rect 43904 12384 43956 12393
rect 24124 12248 24176 12300
rect 24400 12291 24452 12300
rect 24400 12257 24409 12291
rect 24409 12257 24443 12291
rect 24443 12257 24452 12291
rect 24400 12248 24452 12257
rect 37556 12291 37608 12300
rect 37556 12257 37565 12291
rect 37565 12257 37599 12291
rect 37599 12257 37608 12291
rect 37556 12248 37608 12257
rect 45560 12248 45612 12300
rect 45836 12248 45888 12300
rect 48228 12291 48280 12300
rect 48228 12257 48237 12291
rect 48237 12257 48271 12291
rect 48271 12257 48280 12291
rect 48228 12248 48280 12257
rect 52368 12248 52420 12300
rect 56876 12248 56928 12300
rect 57244 12291 57296 12300
rect 57244 12257 57253 12291
rect 57253 12257 57287 12291
rect 57287 12257 57296 12291
rect 57244 12248 57296 12257
rect 3884 12180 3936 12232
rect 5540 12180 5592 12232
rect 9680 12223 9732 12232
rect 9680 12189 9714 12223
rect 9714 12189 9732 12223
rect 9680 12180 9732 12189
rect 13820 12180 13872 12232
rect 4252 12112 4304 12164
rect 6092 12112 6144 12164
rect 14188 12180 14240 12232
rect 16672 12180 16724 12232
rect 25136 12180 25188 12232
rect 27436 12223 27488 12232
rect 27436 12189 27445 12223
rect 27445 12189 27479 12223
rect 27479 12189 27488 12223
rect 27436 12180 27488 12189
rect 28632 12180 28684 12232
rect 29276 12180 29328 12232
rect 17224 12112 17276 12164
rect 23480 12112 23532 12164
rect 30196 12180 30248 12232
rect 32128 12180 32180 12232
rect 34796 12180 34848 12232
rect 40500 12180 40552 12232
rect 42524 12223 42576 12232
rect 42524 12189 42533 12223
rect 42533 12189 42567 12223
rect 42567 12189 42576 12223
rect 42524 12180 42576 12189
rect 51172 12223 51224 12232
rect 51172 12189 51181 12223
rect 51181 12189 51215 12223
rect 51215 12189 51224 12223
rect 51172 12180 51224 12189
rect 53656 12180 53708 12232
rect 55404 12223 55456 12232
rect 55404 12189 55413 12223
rect 55413 12189 55447 12223
rect 55447 12189 55456 12223
rect 55404 12180 55456 12189
rect 56600 12180 56652 12232
rect 57520 12223 57572 12232
rect 57520 12189 57554 12223
rect 57554 12189 57572 12223
rect 57520 12180 57572 12189
rect 31116 12112 31168 12164
rect 35992 12112 36044 12164
rect 38844 12112 38896 12164
rect 41880 12112 41932 12164
rect 7012 12087 7064 12096
rect 7012 12053 7021 12087
rect 7021 12053 7055 12087
rect 7055 12053 7064 12087
rect 7012 12044 7064 12053
rect 10784 12087 10836 12096
rect 10784 12053 10793 12087
rect 10793 12053 10827 12087
rect 10827 12053 10836 12087
rect 10784 12044 10836 12053
rect 17316 12087 17368 12096
rect 17316 12053 17325 12087
rect 17325 12053 17359 12087
rect 17359 12053 17368 12087
rect 17316 12044 17368 12053
rect 25780 12087 25832 12096
rect 25780 12053 25789 12087
rect 25789 12053 25823 12087
rect 25823 12053 25832 12087
rect 25780 12044 25832 12053
rect 30932 12087 30984 12096
rect 30932 12053 30941 12087
rect 30941 12053 30975 12087
rect 30975 12053 30984 12087
rect 30932 12044 30984 12053
rect 31208 12044 31260 12096
rect 36084 12087 36136 12096
rect 36084 12053 36093 12087
rect 36093 12053 36127 12087
rect 36127 12053 36136 12087
rect 36084 12044 36136 12053
rect 47768 12087 47820 12096
rect 47768 12053 47777 12087
rect 47777 12053 47811 12087
rect 47811 12053 47820 12087
rect 47768 12044 47820 12053
rect 50160 12112 50212 12164
rect 52920 12112 52972 12164
rect 53656 12044 53708 12096
rect 54392 12087 54444 12096
rect 54392 12053 54401 12087
rect 54401 12053 54435 12087
rect 54435 12053 54444 12087
rect 54392 12044 54444 12053
rect 56784 12087 56836 12096
rect 56784 12053 56793 12087
rect 56793 12053 56827 12087
rect 56827 12053 56836 12087
rect 56784 12044 56836 12053
rect 58440 12044 58492 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 4252 11883 4304 11892
rect 4252 11849 4261 11883
rect 4261 11849 4295 11883
rect 4295 11849 4304 11883
rect 4252 11840 4304 11849
rect 7748 11883 7800 11892
rect 7748 11849 7757 11883
rect 7757 11849 7791 11883
rect 7791 11849 7800 11883
rect 7748 11840 7800 11849
rect 5356 11772 5408 11824
rect 6368 11772 6420 11824
rect 3884 11704 3936 11756
rect 9772 11840 9824 11892
rect 10784 11772 10836 11824
rect 22376 11840 22428 11892
rect 29092 11840 29144 11892
rect 31116 11883 31168 11892
rect 31116 11849 31125 11883
rect 31125 11849 31159 11883
rect 31159 11849 31168 11883
rect 31116 11840 31168 11849
rect 33416 11840 33468 11892
rect 38844 11883 38896 11892
rect 38844 11849 38853 11883
rect 38853 11849 38887 11883
rect 38887 11849 38896 11883
rect 38844 11840 38896 11849
rect 41880 11883 41932 11892
rect 41880 11849 41889 11883
rect 41889 11849 41923 11883
rect 41923 11849 41932 11883
rect 41880 11840 41932 11849
rect 45468 11840 45520 11892
rect 45744 11840 45796 11892
rect 50160 11840 50212 11892
rect 55588 11840 55640 11892
rect 17316 11772 17368 11824
rect 15476 11704 15528 11756
rect 21272 11704 21324 11756
rect 22192 11772 22244 11824
rect 25780 11772 25832 11824
rect 29368 11772 29420 11824
rect 30932 11772 30984 11824
rect 44272 11772 44324 11824
rect 44548 11815 44600 11824
rect 44548 11781 44582 11815
rect 44582 11781 44600 11815
rect 44548 11772 44600 11781
rect 24124 11747 24176 11756
rect 24124 11713 24133 11747
rect 24133 11713 24167 11747
rect 24167 11713 24176 11747
rect 24124 11704 24176 11713
rect 27436 11704 27488 11756
rect 32128 11747 32180 11756
rect 32128 11713 32137 11747
rect 32137 11713 32171 11747
rect 32171 11713 32180 11747
rect 32128 11704 32180 11713
rect 32404 11747 32456 11756
rect 32404 11713 32438 11747
rect 32438 11713 32456 11747
rect 32404 11704 32456 11713
rect 34244 11747 34296 11756
rect 34244 11713 34278 11747
rect 34278 11713 34296 11747
rect 34244 11704 34296 11713
rect 37556 11704 37608 11756
rect 38752 11704 38804 11756
rect 40500 11747 40552 11756
rect 40500 11713 40509 11747
rect 40509 11713 40543 11747
rect 40543 11713 40552 11747
rect 40500 11704 40552 11713
rect 41880 11704 41932 11756
rect 42524 11704 42576 11756
rect 6092 11636 6144 11688
rect 12164 11679 12216 11688
rect 12164 11645 12173 11679
rect 12173 11645 12207 11679
rect 12207 11645 12216 11679
rect 12164 11636 12216 11645
rect 14004 11679 14056 11688
rect 14004 11645 14013 11679
rect 14013 11645 14047 11679
rect 14047 11645 14056 11679
rect 14004 11636 14056 11645
rect 16672 11679 16724 11688
rect 16672 11645 16681 11679
rect 16681 11645 16715 11679
rect 16715 11645 16724 11679
rect 16672 11636 16724 11645
rect 19892 11679 19944 11688
rect 19892 11645 19901 11679
rect 19901 11645 19935 11679
rect 19935 11645 19944 11679
rect 19892 11636 19944 11645
rect 29552 11636 29604 11688
rect 33968 11679 34020 11688
rect 33968 11645 33977 11679
rect 33977 11645 34011 11679
rect 34011 11645 34020 11679
rect 33968 11636 34020 11645
rect 44916 11704 44968 11756
rect 49608 11704 49660 11756
rect 51172 11772 51224 11824
rect 56784 11772 56836 11824
rect 58440 11815 58492 11824
rect 58440 11781 58449 11815
rect 58449 11781 58483 11815
rect 58483 11781 58492 11815
rect 58440 11772 58492 11781
rect 52092 11704 52144 11756
rect 48596 11636 48648 11688
rect 53288 11636 53340 11688
rect 55404 11704 55456 11756
rect 57244 11704 57296 11756
rect 58624 11747 58676 11756
rect 58624 11713 58633 11747
rect 58633 11713 58667 11747
rect 58667 11713 58676 11747
rect 58624 11704 58676 11713
rect 10784 11543 10836 11552
rect 10784 11509 10793 11543
rect 10793 11509 10827 11543
rect 10827 11509 10836 11543
rect 10784 11500 10836 11509
rect 15384 11543 15436 11552
rect 15384 11509 15393 11543
rect 15393 11509 15427 11543
rect 15427 11509 15436 11543
rect 15384 11500 15436 11509
rect 18052 11543 18104 11552
rect 18052 11509 18061 11543
rect 18061 11509 18095 11543
rect 18095 11509 18104 11543
rect 18052 11500 18104 11509
rect 22100 11500 22152 11552
rect 25504 11543 25556 11552
rect 25504 11509 25513 11543
rect 25513 11509 25547 11543
rect 25547 11509 25556 11543
rect 25504 11500 25556 11509
rect 35348 11543 35400 11552
rect 35348 11509 35357 11543
rect 35357 11509 35391 11543
rect 35391 11509 35400 11543
rect 35348 11500 35400 11509
rect 40408 11500 40460 11552
rect 48412 11500 48464 11552
rect 51172 11500 51224 11552
rect 55956 11500 56008 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 5816 11339 5868 11348
rect 5816 11305 5825 11339
rect 5825 11305 5859 11339
rect 5859 11305 5868 11339
rect 5816 11296 5868 11305
rect 11152 11296 11204 11348
rect 12164 11296 12216 11348
rect 14004 11296 14056 11348
rect 15476 11339 15528 11348
rect 15476 11305 15485 11339
rect 15485 11305 15519 11339
rect 15519 11305 15528 11339
rect 15476 11296 15528 11305
rect 12072 11228 12124 11280
rect 10968 11160 11020 11212
rect 14096 11228 14148 11280
rect 13820 11160 13872 11212
rect 16672 11296 16724 11348
rect 17224 11296 17276 11348
rect 21272 11339 21324 11348
rect 21272 11305 21281 11339
rect 21281 11305 21315 11339
rect 21315 11305 21324 11339
rect 21272 11296 21324 11305
rect 23480 11339 23532 11348
rect 23480 11305 23489 11339
rect 23489 11305 23523 11339
rect 23523 11305 23532 11339
rect 23480 11296 23532 11305
rect 31944 11339 31996 11348
rect 31944 11305 31953 11339
rect 31953 11305 31987 11339
rect 31987 11305 31996 11339
rect 31944 11296 31996 11305
rect 33784 11339 33836 11348
rect 33784 11305 33793 11339
rect 33793 11305 33827 11339
rect 33827 11305 33836 11339
rect 33784 11296 33836 11305
rect 35992 11296 36044 11348
rect 38752 11339 38804 11348
rect 38752 11305 38761 11339
rect 38761 11305 38795 11339
rect 38795 11305 38804 11339
rect 38752 11296 38804 11305
rect 39856 11339 39908 11348
rect 39856 11305 39865 11339
rect 39865 11305 39899 11339
rect 39899 11305 39908 11339
rect 39856 11296 39908 11305
rect 41880 11339 41932 11348
rect 41880 11305 41889 11339
rect 41889 11305 41923 11339
rect 41923 11305 41932 11339
rect 41880 11296 41932 11305
rect 7012 11092 7064 11144
rect 6092 11024 6144 11076
rect 10784 11092 10836 11144
rect 40500 11203 40552 11212
rect 40500 11169 40509 11203
rect 40509 11169 40543 11203
rect 40543 11169 40552 11203
rect 40500 11160 40552 11169
rect 47952 11296 48004 11348
rect 49608 11339 49660 11348
rect 49608 11305 49617 11339
rect 49617 11305 49651 11339
rect 49651 11305 49660 11339
rect 49608 11296 49660 11305
rect 52460 11296 52512 11348
rect 52920 11339 52972 11348
rect 52920 11305 52929 11339
rect 52929 11305 52963 11339
rect 52963 11305 52972 11339
rect 52920 11296 52972 11305
rect 56876 11203 56928 11212
rect 56876 11169 56885 11203
rect 56885 11169 56919 11203
rect 56919 11169 56928 11203
rect 56876 11160 56928 11169
rect 9864 11024 9916 11076
rect 10968 11024 11020 11076
rect 13912 11024 13964 11076
rect 15200 11024 15252 11076
rect 15384 11092 15436 11144
rect 19340 11092 19392 11144
rect 19892 11135 19944 11144
rect 19892 11101 19901 11135
rect 19901 11101 19935 11135
rect 19935 11101 19944 11135
rect 19892 11092 19944 11101
rect 24124 11092 24176 11144
rect 24400 11135 24452 11144
rect 24400 11101 24409 11135
rect 24409 11101 24443 11135
rect 24443 11101 24452 11135
rect 24400 11092 24452 11101
rect 25504 11092 25556 11144
rect 19248 11024 19300 11076
rect 20996 11024 21048 11076
rect 23204 11024 23256 11076
rect 31208 11092 31260 11144
rect 32128 11024 32180 11076
rect 33508 11092 33560 11144
rect 33416 11024 33468 11076
rect 33968 11024 34020 11076
rect 35348 11092 35400 11144
rect 37464 11092 37516 11144
rect 40408 11092 40460 11144
rect 47768 11092 47820 11144
rect 38660 11024 38712 11076
rect 41788 11024 41840 11076
rect 45836 11024 45888 11076
rect 50068 11092 50120 11144
rect 53288 11092 53340 11144
rect 54392 11092 54444 11144
rect 48596 11024 48648 11076
rect 53748 11024 53800 11076
rect 57336 11024 57388 11076
rect 10784 10999 10836 11008
rect 10784 10965 10793 10999
rect 10793 10965 10827 10999
rect 10827 10965 10836 10999
rect 10784 10956 10836 10965
rect 25780 10999 25832 11008
rect 25780 10965 25789 10999
rect 25789 10965 25823 10999
rect 25823 10965 25832 10999
rect 25780 10956 25832 10965
rect 47768 10999 47820 11008
rect 47768 10965 47777 10999
rect 47777 10965 47811 10999
rect 47811 10965 47820 10999
rect 47768 10956 47820 10965
rect 54760 10999 54812 11008
rect 54760 10965 54769 10999
rect 54769 10965 54803 10999
rect 54803 10965 54812 10999
rect 54760 10956 54812 10965
rect 58256 10999 58308 11008
rect 58256 10965 58265 10999
rect 58265 10965 58299 10999
rect 58299 10965 58308 10999
rect 58256 10956 58308 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 15200 10752 15252 10804
rect 20996 10795 21048 10804
rect 20996 10761 21005 10795
rect 21005 10761 21039 10795
rect 21039 10761 21048 10795
rect 20996 10752 21048 10761
rect 23204 10795 23256 10804
rect 23204 10761 23213 10795
rect 23213 10761 23247 10795
rect 23247 10761 23256 10795
rect 23204 10752 23256 10761
rect 33692 10752 33744 10804
rect 38660 10795 38712 10804
rect 38660 10761 38669 10795
rect 38669 10761 38703 10795
rect 38703 10761 38712 10795
rect 38660 10752 38712 10761
rect 41788 10752 41840 10804
rect 10784 10684 10836 10736
rect 14096 10684 14148 10736
rect 18052 10684 18104 10736
rect 19248 10684 19300 10736
rect 20904 10684 20956 10736
rect 22100 10727 22152 10736
rect 22100 10693 22134 10727
rect 22134 10693 22152 10727
rect 22100 10684 22152 10693
rect 25780 10684 25832 10736
rect 9864 10616 9916 10668
rect 11796 10659 11848 10668
rect 11796 10625 11830 10659
rect 11830 10625 11848 10659
rect 11796 10616 11848 10625
rect 16764 10616 16816 10668
rect 20720 10616 20772 10668
rect 24124 10616 24176 10668
rect 27528 10616 27580 10668
rect 29552 10684 29604 10736
rect 34152 10684 34204 10736
rect 36084 10684 36136 10736
rect 48136 10752 48188 10804
rect 50620 10752 50672 10804
rect 51080 10752 51132 10804
rect 55496 10795 55548 10804
rect 55496 10761 55505 10795
rect 55505 10761 55539 10795
rect 55539 10761 55548 10795
rect 55496 10752 55548 10761
rect 57244 10752 57296 10804
rect 47768 10684 47820 10736
rect 30196 10616 30248 10668
rect 32128 10616 32180 10668
rect 38568 10616 38620 10668
rect 40500 10659 40552 10668
rect 40500 10625 40509 10659
rect 40509 10625 40543 10659
rect 40543 10625 40552 10659
rect 40500 10616 40552 10625
rect 41880 10616 41932 10668
rect 45744 10616 45796 10668
rect 48412 10659 48464 10668
rect 48412 10625 48421 10659
rect 48421 10625 48455 10659
rect 48455 10625 48464 10659
rect 48412 10616 48464 10625
rect 50160 10616 50212 10668
rect 55956 10684 56008 10736
rect 58256 10684 58308 10736
rect 52920 10616 52972 10668
rect 53288 10616 53340 10668
rect 10784 10548 10836 10600
rect 13820 10548 13872 10600
rect 19340 10548 19392 10600
rect 20628 10548 20680 10600
rect 33416 10548 33468 10600
rect 37280 10591 37332 10600
rect 37280 10557 37289 10591
rect 37289 10557 37323 10591
rect 37323 10557 37332 10591
rect 37280 10548 37332 10557
rect 48964 10591 49016 10600
rect 48964 10557 48973 10591
rect 48973 10557 49007 10591
rect 49007 10557 49016 10591
rect 48964 10548 49016 10557
rect 10692 10455 10744 10464
rect 10692 10421 10701 10455
rect 10701 10421 10735 10455
rect 10735 10421 10744 10455
rect 10692 10412 10744 10421
rect 14372 10412 14424 10464
rect 18052 10455 18104 10464
rect 18052 10421 18061 10455
rect 18061 10421 18095 10455
rect 18095 10421 18104 10455
rect 18052 10412 18104 10421
rect 18604 10412 18656 10464
rect 25412 10455 25464 10464
rect 25412 10421 25421 10455
rect 25421 10421 25455 10455
rect 25455 10421 25464 10455
rect 25412 10412 25464 10421
rect 29828 10412 29880 10464
rect 35624 10455 35676 10464
rect 35624 10421 35633 10455
rect 35633 10421 35667 10455
rect 35667 10421 35676 10455
rect 35624 10412 35676 10421
rect 43352 10412 43404 10464
rect 52184 10455 52236 10464
rect 52184 10421 52193 10455
rect 52193 10421 52227 10455
rect 52227 10421 52236 10455
rect 52184 10412 52236 10421
rect 56876 10412 56928 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 6092 10115 6144 10124
rect 6092 10081 6101 10115
rect 6101 10081 6135 10115
rect 6135 10081 6144 10115
rect 6092 10072 6144 10081
rect 9036 10072 9088 10124
rect 9864 10208 9916 10260
rect 13912 10208 13964 10260
rect 17960 10251 18012 10260
rect 17960 10217 17969 10251
rect 17969 10217 18003 10251
rect 18003 10217 18012 10251
rect 17960 10208 18012 10217
rect 19340 10208 19392 10260
rect 20628 10208 20680 10260
rect 26240 10208 26292 10260
rect 10968 10115 11020 10124
rect 10968 10081 10977 10115
rect 10977 10081 11011 10115
rect 11011 10081 11020 10115
rect 10968 10072 11020 10081
rect 10692 10004 10744 10056
rect 14096 10004 14148 10056
rect 16672 10004 16724 10056
rect 18052 10004 18104 10056
rect 18604 10004 18656 10056
rect 19432 10004 19484 10056
rect 29552 10115 29604 10124
rect 29552 10081 29561 10115
rect 29561 10081 29595 10115
rect 29595 10081 29604 10115
rect 29552 10072 29604 10081
rect 37464 10208 37516 10260
rect 38568 10251 38620 10260
rect 38568 10217 38577 10251
rect 38577 10217 38611 10251
rect 38611 10217 38620 10251
rect 38568 10208 38620 10217
rect 47860 10208 47912 10260
rect 48596 10251 48648 10260
rect 48596 10217 48605 10251
rect 48605 10217 48639 10251
rect 48639 10217 48648 10251
rect 48596 10208 48648 10217
rect 52920 10251 52972 10260
rect 52920 10217 52929 10251
rect 52929 10217 52963 10251
rect 52963 10217 52972 10251
rect 52920 10208 52972 10217
rect 53748 10208 53800 10260
rect 53288 10072 53340 10124
rect 56876 10115 56928 10124
rect 56876 10081 56885 10115
rect 56885 10081 56919 10115
rect 56919 10081 56928 10115
rect 56876 10072 56928 10081
rect 24400 10047 24452 10056
rect 24400 10013 24409 10047
rect 24409 10013 24443 10047
rect 24443 10013 24452 10047
rect 24400 10004 24452 10013
rect 25412 10004 25464 10056
rect 26240 10004 26292 10056
rect 33416 10004 33468 10056
rect 45744 10004 45796 10056
rect 48136 10004 48188 10056
rect 51540 10047 51592 10056
rect 51540 10013 51549 10047
rect 51549 10013 51583 10047
rect 51583 10013 51592 10047
rect 51540 10004 51592 10013
rect 54760 10004 54812 10056
rect 7288 9936 7340 9988
rect 11060 9936 11112 9988
rect 15476 9936 15528 9988
rect 30840 9936 30892 9988
rect 34060 9936 34112 9988
rect 38660 9936 38712 9988
rect 43352 9979 43404 9988
rect 43352 9945 43386 9979
rect 43386 9945 43404 9979
rect 43352 9936 43404 9945
rect 45652 9936 45704 9988
rect 53748 9936 53800 9988
rect 7472 9911 7524 9920
rect 7472 9877 7481 9911
rect 7481 9877 7515 9911
rect 7515 9877 7524 9911
rect 7472 9868 7524 9877
rect 10508 9911 10560 9920
rect 10508 9877 10517 9911
rect 10517 9877 10551 9911
rect 10551 9877 10560 9911
rect 10508 9868 10560 9877
rect 10600 9868 10652 9920
rect 25136 9868 25188 9920
rect 32220 9868 32272 9920
rect 34152 9911 34204 9920
rect 34152 9877 34161 9911
rect 34161 9877 34195 9911
rect 34195 9877 34204 9911
rect 34152 9868 34204 9877
rect 45376 9868 45428 9920
rect 58256 9911 58308 9920
rect 58256 9877 58265 9911
rect 58265 9877 58299 9911
rect 58299 9877 58308 9911
rect 58256 9868 58308 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 20720 9707 20772 9716
rect 20720 9673 20729 9707
rect 20729 9673 20763 9707
rect 20763 9673 20772 9707
rect 20720 9664 20772 9673
rect 30196 9707 30248 9716
rect 30196 9673 30205 9707
rect 30205 9673 30239 9707
rect 30239 9673 30248 9707
rect 30196 9664 30248 9673
rect 38660 9707 38712 9716
rect 38660 9673 38669 9707
rect 38669 9673 38703 9707
rect 38703 9673 38712 9707
rect 38660 9664 38712 9673
rect 41880 9707 41932 9716
rect 41880 9673 41889 9707
rect 41889 9673 41923 9707
rect 41923 9673 41932 9707
rect 41880 9664 41932 9673
rect 45652 9707 45704 9716
rect 45652 9673 45661 9707
rect 45661 9673 45695 9707
rect 45695 9673 45704 9707
rect 45652 9664 45704 9673
rect 50160 9664 50212 9716
rect 10508 9596 10560 9648
rect 12440 9596 12492 9648
rect 18144 9596 18196 9648
rect 12808 9528 12860 9580
rect 16672 9571 16724 9580
rect 16672 9537 16681 9571
rect 16681 9537 16715 9571
rect 16715 9537 16724 9571
rect 16672 9528 16724 9537
rect 20536 9528 20588 9580
rect 24400 9596 24452 9648
rect 24952 9528 25004 9580
rect 26240 9596 26292 9648
rect 25780 9528 25832 9580
rect 27528 9596 27580 9648
rect 35624 9596 35676 9648
rect 27620 9528 27672 9580
rect 29092 9571 29144 9580
rect 29092 9537 29126 9571
rect 29126 9537 29144 9571
rect 37280 9571 37332 9580
rect 29092 9528 29144 9537
rect 37280 9537 37289 9571
rect 37289 9537 37323 9571
rect 37323 9537 37332 9571
rect 37280 9528 37332 9537
rect 37372 9528 37424 9580
rect 40500 9571 40552 9580
rect 40500 9537 40509 9571
rect 40509 9537 40543 9571
rect 40543 9537 40552 9571
rect 40500 9528 40552 9537
rect 42064 9528 42116 9580
rect 43904 9528 43956 9580
rect 51172 9596 51224 9648
rect 53656 9639 53708 9648
rect 53656 9605 53690 9639
rect 53690 9605 53708 9639
rect 53656 9596 53708 9605
rect 58256 9596 58308 9648
rect 45652 9528 45704 9580
rect 48964 9571 49016 9580
rect 48964 9537 48973 9571
rect 48973 9537 49007 9571
rect 49007 9537 49016 9571
rect 48964 9528 49016 9537
rect 5908 9460 5960 9512
rect 9036 9503 9088 9512
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 19340 9503 19392 9512
rect 19340 9469 19349 9503
rect 19349 9469 19383 9503
rect 19383 9469 19392 9503
rect 19340 9460 19392 9469
rect 18236 9392 18288 9444
rect 7748 9367 7800 9376
rect 7748 9333 7757 9367
rect 7757 9333 7791 9367
rect 7791 9333 7800 9367
rect 7748 9324 7800 9333
rect 9220 9324 9272 9376
rect 14096 9324 14148 9376
rect 24584 9367 24636 9376
rect 24584 9333 24593 9367
rect 24593 9333 24627 9367
rect 24627 9333 24636 9367
rect 24584 9324 24636 9333
rect 26516 9324 26568 9376
rect 28356 9367 28408 9376
rect 28356 9333 28365 9367
rect 28365 9333 28399 9367
rect 28399 9333 28408 9367
rect 28356 9324 28408 9333
rect 33416 9460 33468 9512
rect 29000 9324 29052 9376
rect 34060 9324 34112 9376
rect 43812 9367 43864 9376
rect 43812 9333 43821 9367
rect 43821 9333 43855 9367
rect 43855 9333 43864 9367
rect 43812 9324 43864 9333
rect 52552 9528 52604 9580
rect 53012 9460 53064 9512
rect 55312 9460 55364 9512
rect 52092 9392 52144 9444
rect 57336 9435 57388 9444
rect 57336 9401 57345 9435
rect 57345 9401 57379 9435
rect 57379 9401 57388 9435
rect 57336 9392 57388 9401
rect 51172 9324 51224 9376
rect 51540 9324 51592 9376
rect 53748 9324 53800 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 7288 9163 7340 9172
rect 7288 9129 7297 9163
rect 7297 9129 7331 9163
rect 7331 9129 7340 9163
rect 7288 9120 7340 9129
rect 11060 9120 11112 9172
rect 15476 9163 15528 9172
rect 15476 9129 15485 9163
rect 15485 9129 15519 9163
rect 15519 9129 15528 9163
rect 15476 9120 15528 9129
rect 25780 9163 25832 9172
rect 25780 9129 25789 9163
rect 25789 9129 25823 9163
rect 25823 9129 25832 9163
rect 25780 9120 25832 9129
rect 27620 9163 27672 9172
rect 27620 9129 27629 9163
rect 27629 9129 27663 9163
rect 27663 9129 27672 9163
rect 27620 9120 27672 9129
rect 42064 9163 42116 9172
rect 42064 9129 42073 9163
rect 42073 9129 42107 9163
rect 42107 9129 42116 9163
rect 42064 9120 42116 9129
rect 43904 9163 43956 9172
rect 43904 9129 43913 9163
rect 43913 9129 43947 9163
rect 43947 9129 43956 9163
rect 43904 9120 43956 9129
rect 52552 9163 52604 9172
rect 52552 9129 52561 9163
rect 52561 9129 52595 9163
rect 52595 9129 52604 9163
rect 52552 9120 52604 9129
rect 5356 8984 5408 9036
rect 5908 9027 5960 9036
rect 5908 8993 5917 9027
rect 5917 8993 5951 9027
rect 5951 8993 5960 9027
rect 5908 8984 5960 8993
rect 19340 8984 19392 9036
rect 7748 8916 7800 8968
rect 8668 8916 8720 8968
rect 9220 8959 9272 8968
rect 9220 8925 9254 8959
rect 9254 8925 9272 8959
rect 9220 8916 9272 8925
rect 10876 8916 10928 8968
rect 14096 8959 14148 8968
rect 14096 8925 14105 8959
rect 14105 8925 14139 8959
rect 14139 8925 14148 8959
rect 14096 8916 14148 8925
rect 14372 8959 14424 8968
rect 14372 8925 14406 8959
rect 14406 8925 14424 8959
rect 14372 8916 14424 8925
rect 26240 9027 26292 9036
rect 26240 8993 26249 9027
rect 26249 8993 26283 9027
rect 26283 8993 26292 9027
rect 26240 8984 26292 8993
rect 40500 8984 40552 9036
rect 51172 9027 51224 9036
rect 23848 8916 23900 8968
rect 24400 8959 24452 8968
rect 24400 8925 24409 8959
rect 24409 8925 24443 8959
rect 24443 8925 24452 8959
rect 24400 8916 24452 8925
rect 25136 8916 25188 8968
rect 26516 8959 26568 8968
rect 26516 8925 26550 8959
rect 26550 8925 26568 8959
rect 26516 8916 26568 8925
rect 29644 8916 29696 8968
rect 32312 8916 32364 8968
rect 5632 8848 5684 8900
rect 10416 8848 10468 8900
rect 22008 8848 22060 8900
rect 23388 8848 23440 8900
rect 30472 8848 30524 8900
rect 5448 8823 5500 8832
rect 5448 8789 5457 8823
rect 5457 8789 5491 8823
rect 5491 8789 5500 8823
rect 5448 8780 5500 8789
rect 12164 8823 12216 8832
rect 12164 8789 12173 8823
rect 12173 8789 12207 8823
rect 12207 8789 12216 8823
rect 12164 8780 12216 8789
rect 21732 8823 21784 8832
rect 21732 8789 21741 8823
rect 21741 8789 21775 8823
rect 21775 8789 21784 8823
rect 21732 8780 21784 8789
rect 22192 8780 22244 8832
rect 30932 8823 30984 8832
rect 30932 8789 30941 8823
rect 30941 8789 30975 8823
rect 30975 8789 30984 8823
rect 30932 8780 30984 8789
rect 33416 8780 33468 8832
rect 34428 8916 34480 8968
rect 35808 8916 35860 8968
rect 51172 8993 51181 9027
rect 51181 8993 51215 9027
rect 51215 8993 51224 9027
rect 51172 8984 51224 8993
rect 45744 8916 45796 8968
rect 46848 8959 46900 8968
rect 46848 8925 46857 8959
rect 46857 8925 46891 8959
rect 46891 8925 46900 8959
rect 46848 8916 46900 8925
rect 34796 8848 34848 8900
rect 36636 8848 36688 8900
rect 41880 8848 41932 8900
rect 41972 8848 42024 8900
rect 44180 8848 44232 8900
rect 47124 8891 47176 8900
rect 47124 8857 47158 8891
rect 47158 8857 47176 8891
rect 52184 8916 52236 8968
rect 53012 8959 53064 8968
rect 53012 8925 53021 8959
rect 53021 8925 53055 8959
rect 53055 8925 53064 8959
rect 53012 8916 53064 8925
rect 55312 8959 55364 8968
rect 55312 8925 55321 8959
rect 55321 8925 55355 8959
rect 55355 8925 55364 8959
rect 55312 8916 55364 8925
rect 47124 8848 47176 8857
rect 52644 8848 52696 8900
rect 54116 8848 54168 8900
rect 56600 8848 56652 8900
rect 58440 8848 58492 8900
rect 36084 8823 36136 8832
rect 36084 8789 36093 8823
rect 36093 8789 36127 8823
rect 36127 8789 36136 8823
rect 36084 8780 36136 8789
rect 37924 8823 37976 8832
rect 37924 8789 37933 8823
rect 37933 8789 37967 8823
rect 37967 8789 37976 8823
rect 37924 8780 37976 8789
rect 46388 8823 46440 8832
rect 46388 8789 46397 8823
rect 46397 8789 46431 8823
rect 46431 8789 46440 8823
rect 46388 8780 46440 8789
rect 47400 8780 47452 8832
rect 54392 8823 54444 8832
rect 54392 8789 54401 8823
rect 54401 8789 54435 8823
rect 54435 8789 54444 8823
rect 54392 8780 54444 8789
rect 55864 8780 55916 8832
rect 58532 8823 58584 8832
rect 58532 8789 58541 8823
rect 58541 8789 58575 8823
rect 58575 8789 58584 8823
rect 58532 8780 58584 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 10416 8619 10468 8628
rect 10416 8585 10425 8619
rect 10425 8585 10459 8619
rect 10459 8585 10468 8619
rect 10416 8576 10468 8585
rect 12808 8576 12860 8628
rect 5448 8508 5500 8560
rect 7472 8508 7524 8560
rect 10600 8508 10652 8560
rect 12164 8508 12216 8560
rect 5264 8440 5316 8492
rect 16028 8440 16080 8492
rect 5908 8372 5960 8424
rect 8668 8372 8720 8424
rect 12164 8372 12216 8424
rect 14096 8372 14148 8424
rect 17316 8372 17368 8424
rect 19340 8576 19392 8628
rect 20536 8619 20588 8628
rect 20536 8585 20545 8619
rect 20545 8585 20579 8619
rect 20579 8585 20588 8619
rect 20536 8576 20588 8585
rect 23388 8619 23440 8628
rect 23388 8585 23397 8619
rect 23397 8585 23431 8619
rect 23431 8585 23440 8619
rect 23388 8576 23440 8585
rect 24952 8576 25004 8628
rect 21732 8508 21784 8560
rect 24584 8508 24636 8560
rect 28540 8576 28592 8628
rect 34796 8619 34848 8628
rect 34796 8585 34805 8619
rect 34805 8585 34839 8619
rect 34839 8585 34848 8619
rect 34796 8576 34848 8585
rect 36636 8619 36688 8628
rect 36636 8585 36645 8619
rect 36645 8585 36679 8619
rect 36679 8585 36688 8619
rect 36636 8576 36688 8585
rect 45652 8619 45704 8628
rect 45652 8585 45661 8619
rect 45661 8585 45695 8619
rect 45695 8585 45704 8619
rect 45652 8576 45704 8585
rect 54116 8619 54168 8628
rect 34152 8508 34204 8560
rect 37924 8508 37976 8560
rect 46388 8508 46440 8560
rect 54116 8585 54125 8619
rect 54125 8585 54159 8619
rect 54159 8585 54168 8619
rect 54116 8576 54168 8585
rect 53840 8508 53892 8560
rect 25780 8440 25832 8492
rect 26240 8440 26292 8492
rect 27620 8440 27672 8492
rect 34428 8440 34480 8492
rect 35992 8440 36044 8492
rect 37280 8483 37332 8492
rect 37280 8449 37289 8483
rect 37289 8449 37323 8483
rect 37323 8449 37332 8483
rect 37280 8440 37332 8449
rect 21640 8372 21692 8424
rect 23848 8415 23900 8424
rect 23848 8381 23857 8415
rect 23857 8381 23891 8415
rect 23891 8381 23900 8415
rect 23848 8372 23900 8381
rect 28724 8372 28776 8424
rect 33416 8415 33468 8424
rect 33416 8381 33425 8415
rect 33425 8381 33459 8415
rect 33459 8381 33468 8415
rect 33416 8372 33468 8381
rect 38844 8440 38896 8492
rect 41420 8440 41472 8492
rect 45744 8440 45796 8492
rect 46848 8440 46900 8492
rect 48228 8440 48280 8492
rect 50160 8440 50212 8492
rect 52736 8483 52788 8492
rect 52736 8449 52745 8483
rect 52745 8449 52779 8483
rect 52779 8449 52788 8483
rect 52736 8440 52788 8449
rect 54116 8440 54168 8492
rect 40500 8372 40552 8424
rect 5448 8304 5500 8356
rect 7748 8279 7800 8288
rect 7748 8245 7757 8279
rect 7757 8245 7791 8279
rect 7791 8245 7800 8279
rect 7748 8236 7800 8245
rect 13820 8236 13872 8288
rect 38660 8279 38712 8288
rect 38660 8245 38669 8279
rect 38669 8245 38703 8279
rect 38703 8245 38712 8279
rect 38660 8236 38712 8245
rect 40500 8279 40552 8288
rect 40500 8245 40509 8279
rect 40509 8245 40543 8279
rect 40543 8245 40552 8279
rect 40500 8236 40552 8245
rect 43628 8304 43680 8356
rect 42800 8236 42852 8288
rect 50804 8279 50856 8288
rect 50804 8245 50813 8279
rect 50813 8245 50847 8279
rect 50847 8245 50856 8279
rect 50804 8236 50856 8245
rect 55312 8236 55364 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 5632 8032 5684 8084
rect 11796 8032 11848 8084
rect 22008 8032 22060 8084
rect 25780 8075 25832 8084
rect 25780 8041 25789 8075
rect 25789 8041 25823 8075
rect 25823 8041 25832 8075
rect 25780 8032 25832 8041
rect 27620 8075 27672 8084
rect 27620 8041 27629 8075
rect 27629 8041 27663 8075
rect 27663 8041 27672 8075
rect 27620 8032 27672 8041
rect 30472 8032 30524 8084
rect 35992 8032 36044 8084
rect 38844 8075 38896 8084
rect 38844 8041 38853 8075
rect 38853 8041 38887 8075
rect 38887 8041 38896 8075
rect 38844 8032 38896 8041
rect 42800 8032 42852 8084
rect 47124 8032 47176 8084
rect 48228 8075 48280 8084
rect 48228 8041 48237 8075
rect 48237 8041 48271 8075
rect 48271 8041 48280 8075
rect 48228 8032 48280 8041
rect 54116 8075 54168 8084
rect 54116 8041 54125 8075
rect 54125 8041 54159 8075
rect 54159 8041 54168 8075
rect 54116 8032 54168 8041
rect 56600 8032 56652 8084
rect 58440 8032 58492 8084
rect 26240 7939 26292 7948
rect 26240 7905 26249 7939
rect 26249 7905 26283 7939
rect 26283 7905 26292 7939
rect 46848 7939 46900 7948
rect 26240 7896 26292 7905
rect 46848 7905 46857 7939
rect 46857 7905 46891 7939
rect 46891 7905 46900 7939
rect 46848 7896 46900 7905
rect 50160 7939 50212 7948
rect 50160 7905 50169 7939
rect 50169 7905 50203 7939
rect 50203 7905 50212 7939
rect 50160 7896 50212 7905
rect 52644 7896 52696 7948
rect 1860 7871 1912 7880
rect 1860 7837 1869 7871
rect 1869 7837 1903 7871
rect 1903 7837 1912 7871
rect 1860 7828 1912 7837
rect 4160 7828 4212 7880
rect 5356 7828 5408 7880
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 7748 7828 7800 7880
rect 12164 7871 12216 7880
rect 12164 7837 12173 7871
rect 12173 7837 12207 7871
rect 12207 7837 12216 7871
rect 12164 7828 12216 7837
rect 16856 7828 16908 7880
rect 17316 7828 17368 7880
rect 21640 7871 21692 7880
rect 21640 7837 21649 7871
rect 21649 7837 21683 7871
rect 21683 7837 21692 7871
rect 21640 7828 21692 7837
rect 22192 7828 22244 7880
rect 24308 7828 24360 7880
rect 3240 7735 3292 7744
rect 3240 7701 3249 7735
rect 3249 7701 3283 7735
rect 3283 7701 3292 7735
rect 3240 7692 3292 7701
rect 6552 7760 6604 7812
rect 12256 7760 12308 7812
rect 13084 7760 13136 7812
rect 13544 7735 13596 7744
rect 13544 7701 13553 7735
rect 13553 7701 13587 7735
rect 13587 7701 13596 7735
rect 13544 7692 13596 7701
rect 14832 7760 14884 7812
rect 16212 7760 16264 7812
rect 18328 7760 18380 7812
rect 21088 7760 21140 7812
rect 22008 7760 22060 7812
rect 25228 7760 25280 7812
rect 28356 7828 28408 7880
rect 29828 7871 29880 7880
rect 29828 7837 29862 7871
rect 29862 7837 29880 7871
rect 26976 7760 27028 7812
rect 29828 7828 29880 7837
rect 32128 7871 32180 7880
rect 32128 7837 32137 7871
rect 32137 7837 32171 7871
rect 32171 7837 32180 7871
rect 32128 7828 32180 7837
rect 32220 7828 32272 7880
rect 33416 7760 33468 7812
rect 36084 7828 36136 7880
rect 35808 7760 35860 7812
rect 38660 7828 38712 7880
rect 41696 7828 41748 7880
rect 45744 7828 45796 7880
rect 47400 7828 47452 7880
rect 55312 7871 55364 7880
rect 55312 7837 55321 7871
rect 55321 7837 55355 7871
rect 55355 7837 55364 7871
rect 55312 7828 55364 7837
rect 45376 7760 45428 7812
rect 50620 7760 50672 7812
rect 54024 7760 54076 7812
rect 55956 7760 56008 7812
rect 56784 7760 56836 7812
rect 15844 7735 15896 7744
rect 15844 7701 15853 7735
rect 15853 7701 15887 7735
rect 15887 7701 15896 7735
rect 15844 7692 15896 7701
rect 17684 7735 17736 7744
rect 17684 7701 17693 7735
rect 17693 7701 17727 7735
rect 17727 7701 17736 7735
rect 17684 7692 17736 7701
rect 20720 7735 20772 7744
rect 20720 7701 20729 7735
rect 20729 7701 20763 7735
rect 20763 7701 20772 7735
rect 20720 7692 20772 7701
rect 33508 7735 33560 7744
rect 33508 7701 33517 7735
rect 33517 7701 33551 7735
rect 33551 7701 33560 7735
rect 33508 7692 33560 7701
rect 51172 7692 51224 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 5356 7531 5408 7540
rect 5356 7497 5365 7531
rect 5365 7497 5399 7531
rect 5399 7497 5408 7531
rect 5356 7488 5408 7497
rect 21088 7531 21140 7540
rect 21088 7497 21097 7531
rect 21097 7497 21131 7531
rect 21131 7497 21140 7531
rect 21088 7488 21140 7497
rect 25228 7531 25280 7540
rect 25228 7497 25237 7531
rect 25237 7497 25271 7531
rect 25271 7497 25280 7531
rect 25228 7488 25280 7497
rect 29092 7488 29144 7540
rect 37372 7488 37424 7540
rect 41420 7488 41472 7540
rect 41880 7531 41932 7540
rect 41880 7497 41889 7531
rect 41889 7497 41923 7531
rect 41923 7497 41932 7531
rect 41880 7488 41932 7497
rect 44180 7531 44232 7540
rect 44180 7497 44189 7531
rect 44189 7497 44223 7531
rect 44223 7497 44232 7531
rect 44180 7488 44232 7497
rect 50620 7488 50672 7540
rect 54024 7488 54076 7540
rect 55956 7531 56008 7540
rect 55956 7497 55965 7531
rect 55965 7497 55999 7531
rect 55999 7497 56008 7531
rect 55956 7488 56008 7497
rect 3240 7420 3292 7472
rect 7196 7420 7248 7472
rect 13820 7420 13872 7472
rect 17684 7420 17736 7472
rect 20720 7420 20772 7472
rect 1860 7352 1912 7404
rect 8392 7352 8444 7404
rect 8668 7352 8720 7404
rect 10784 7352 10836 7404
rect 14832 7352 14884 7404
rect 17316 7352 17368 7404
rect 21180 7352 21232 7404
rect 24400 7420 24452 7472
rect 28540 7420 28592 7472
rect 30932 7420 30984 7472
rect 33508 7420 33560 7472
rect 35808 7420 35860 7472
rect 40500 7420 40552 7472
rect 43812 7420 43864 7472
rect 50804 7420 50856 7472
rect 52644 7420 52696 7472
rect 5908 7284 5960 7336
rect 6736 7327 6788 7336
rect 6736 7293 6745 7327
rect 6745 7293 6779 7327
rect 6779 7293 6788 7327
rect 6736 7284 6788 7293
rect 19708 7327 19760 7336
rect 4068 7148 4120 7200
rect 8852 7148 8904 7200
rect 9956 7191 10008 7200
rect 9956 7157 9965 7191
rect 9965 7157 9999 7191
rect 9999 7157 10008 7191
rect 9956 7148 10008 7157
rect 12164 7148 12216 7200
rect 19708 7293 19717 7327
rect 19717 7293 19751 7327
rect 19751 7293 19760 7327
rect 19708 7284 19760 7293
rect 23848 7327 23900 7336
rect 23848 7293 23857 7327
rect 23857 7293 23891 7327
rect 23891 7293 23900 7327
rect 25780 7352 25832 7404
rect 26976 7395 27028 7404
rect 26976 7361 26985 7395
rect 26985 7361 27019 7395
rect 27019 7361 27028 7395
rect 26976 7352 27028 7361
rect 35348 7395 35400 7404
rect 35348 7361 35357 7395
rect 35357 7361 35391 7395
rect 35391 7361 35400 7395
rect 35348 7352 35400 7361
rect 39212 7352 39264 7404
rect 43536 7352 43588 7404
rect 47124 7352 47176 7404
rect 51540 7352 51592 7404
rect 52736 7395 52788 7404
rect 52736 7361 52745 7395
rect 52745 7361 52779 7395
rect 52779 7361 52788 7395
rect 52736 7352 52788 7361
rect 54208 7352 54260 7404
rect 54392 7420 54444 7472
rect 55312 7352 55364 7404
rect 23848 7284 23900 7293
rect 29184 7284 29236 7336
rect 32128 7327 32180 7336
rect 32128 7293 32137 7327
rect 32137 7293 32171 7327
rect 32171 7293 32180 7327
rect 32128 7284 32180 7293
rect 38660 7327 38712 7336
rect 38660 7293 38669 7327
rect 38669 7293 38703 7327
rect 38703 7293 38712 7327
rect 38660 7284 38712 7293
rect 40408 7284 40460 7336
rect 42800 7327 42852 7336
rect 42800 7293 42809 7327
rect 42809 7293 42843 7327
rect 42843 7293 42852 7327
rect 42800 7284 42852 7293
rect 45652 7327 45704 7336
rect 45652 7293 45661 7327
rect 45661 7293 45695 7327
rect 45695 7293 45704 7327
rect 45652 7284 45704 7293
rect 46848 7284 46900 7336
rect 47492 7284 47544 7336
rect 50160 7284 50212 7336
rect 30840 7216 30892 7268
rect 14096 7148 14148 7200
rect 14280 7191 14332 7200
rect 14280 7157 14289 7191
rect 14289 7157 14323 7191
rect 14323 7157 14332 7191
rect 14280 7148 14332 7157
rect 16120 7191 16172 7200
rect 16120 7157 16129 7191
rect 16129 7157 16163 7191
rect 16163 7157 16172 7191
rect 16120 7148 16172 7157
rect 19248 7191 19300 7200
rect 19248 7157 19257 7191
rect 19257 7157 19291 7191
rect 19291 7157 19300 7191
rect 19248 7148 19300 7157
rect 32312 7148 32364 7200
rect 47676 7148 47728 7200
rect 52184 7191 52236 7200
rect 52184 7157 52193 7191
rect 52193 7157 52227 7191
rect 52227 7157 52236 7191
rect 52184 7148 52236 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 6552 6987 6604 6996
rect 6552 6953 6561 6987
rect 6561 6953 6595 6987
rect 6595 6953 6604 6987
rect 6552 6944 6604 6953
rect 8392 6987 8444 6996
rect 8392 6953 8401 6987
rect 8401 6953 8435 6987
rect 8435 6953 8444 6987
rect 8392 6944 8444 6953
rect 13084 6944 13136 6996
rect 21180 6987 21232 6996
rect 21180 6953 21189 6987
rect 21189 6953 21223 6987
rect 21223 6953 21232 6987
rect 21180 6944 21232 6953
rect 25780 6987 25832 6996
rect 25780 6953 25789 6987
rect 25789 6953 25823 6987
rect 25823 6953 25832 6987
rect 25780 6944 25832 6953
rect 39212 6987 39264 6996
rect 39212 6953 39221 6987
rect 39221 6953 39255 6987
rect 39255 6953 39264 6987
rect 39212 6944 39264 6953
rect 47124 6987 47176 6996
rect 47124 6953 47133 6987
rect 47133 6953 47167 6987
rect 47167 6953 47176 6987
rect 47124 6944 47176 6953
rect 51540 6987 51592 6996
rect 51540 6953 51549 6987
rect 51549 6953 51583 6987
rect 51583 6953 51592 6987
rect 51540 6944 51592 6953
rect 54208 6987 54260 6996
rect 54208 6953 54217 6987
rect 54217 6953 54251 6987
rect 54251 6953 54260 6987
rect 54208 6944 54260 6953
rect 56784 6944 56836 6996
rect 14096 6808 14148 6860
rect 14740 6808 14792 6860
rect 17316 6851 17368 6860
rect 17316 6817 17325 6851
rect 17325 6817 17359 6851
rect 17359 6817 17368 6851
rect 17316 6808 17368 6817
rect 24400 6851 24452 6860
rect 24400 6817 24409 6851
rect 24409 6817 24443 6851
rect 24443 6817 24452 6851
rect 24400 6808 24452 6817
rect 28724 6808 28776 6860
rect 29644 6808 29696 6860
rect 32128 6808 32180 6860
rect 40592 6851 40644 6860
rect 40592 6817 40601 6851
rect 40601 6817 40635 6851
rect 40635 6817 40644 6851
rect 40592 6808 40644 6817
rect 52736 6808 52788 6860
rect 1952 6740 2004 6792
rect 5264 6672 5316 6724
rect 5448 6783 5500 6792
rect 5448 6749 5482 6783
rect 5482 6749 5500 6783
rect 5448 6740 5500 6749
rect 6736 6740 6788 6792
rect 8668 6740 8720 6792
rect 8944 6783 8996 6792
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 8944 6740 8996 6749
rect 10692 6740 10744 6792
rect 11888 6740 11940 6792
rect 12164 6783 12216 6792
rect 12164 6749 12173 6783
rect 12173 6749 12207 6783
rect 12207 6749 12216 6783
rect 12164 6740 12216 6749
rect 14280 6740 14332 6792
rect 16120 6740 16172 6792
rect 19248 6740 19300 6792
rect 19708 6740 19760 6792
rect 22008 6740 22060 6792
rect 24308 6740 24360 6792
rect 28816 6740 28868 6792
rect 29184 6740 29236 6792
rect 30288 6740 30340 6792
rect 32312 6740 32364 6792
rect 35808 6740 35860 6792
rect 37740 6740 37792 6792
rect 38660 6740 38712 6792
rect 43076 6783 43128 6792
rect 43076 6749 43085 6783
rect 43085 6749 43119 6783
rect 43119 6749 43128 6783
rect 43076 6740 43128 6749
rect 5816 6672 5868 6724
rect 7748 6672 7800 6724
rect 10232 6672 10284 6724
rect 20904 6672 20956 6724
rect 23480 6672 23532 6724
rect 25780 6672 25832 6724
rect 31024 6672 31076 6724
rect 3240 6647 3292 6656
rect 3240 6613 3249 6647
rect 3249 6613 3283 6647
rect 3283 6613 3292 6647
rect 3240 6604 3292 6613
rect 10324 6647 10376 6656
rect 10324 6613 10333 6647
rect 10333 6613 10367 6647
rect 10367 6613 10376 6647
rect 10324 6604 10376 6613
rect 16580 6604 16632 6656
rect 18696 6647 18748 6656
rect 18696 6613 18705 6647
rect 18705 6613 18739 6647
rect 18739 6613 18748 6647
rect 18696 6604 18748 6613
rect 23848 6647 23900 6656
rect 23848 6613 23857 6647
rect 23857 6613 23891 6647
rect 23891 6613 23900 6647
rect 23848 6604 23900 6613
rect 29000 6647 29052 6656
rect 29000 6613 29009 6647
rect 29009 6613 29043 6647
rect 29043 6613 29052 6647
rect 29000 6604 29052 6613
rect 36728 6672 36780 6724
rect 34060 6647 34112 6656
rect 34060 6613 34069 6647
rect 34069 6613 34103 6647
rect 34103 6613 34112 6647
rect 34060 6604 34112 6613
rect 43628 6740 43680 6792
rect 43904 6740 43956 6792
rect 45652 6740 45704 6792
rect 47492 6740 47544 6792
rect 47860 6783 47912 6792
rect 47860 6749 47894 6783
rect 47894 6749 47912 6783
rect 47860 6740 47912 6749
rect 49792 6740 49844 6792
rect 50160 6783 50212 6792
rect 50160 6749 50169 6783
rect 50169 6749 50203 6783
rect 50203 6749 50212 6783
rect 50160 6740 50212 6749
rect 51172 6740 51224 6792
rect 55312 6783 55364 6792
rect 55312 6749 55321 6783
rect 55321 6749 55355 6783
rect 55355 6749 55364 6783
rect 55312 6740 55364 6749
rect 55864 6740 55916 6792
rect 45284 6672 45336 6724
rect 49332 6672 49384 6724
rect 54668 6672 54720 6724
rect 58532 6740 58584 6792
rect 41972 6647 42024 6656
rect 41972 6613 41981 6647
rect 41981 6613 42015 6647
rect 42015 6613 42024 6647
rect 41972 6604 42024 6613
rect 44456 6647 44508 6656
rect 44456 6613 44465 6647
rect 44465 6613 44499 6647
rect 44499 6613 44508 6647
rect 44456 6604 44508 6613
rect 48964 6647 49016 6656
rect 48964 6613 48973 6647
rect 48973 6613 49007 6647
rect 49007 6613 49016 6647
rect 48964 6604 49016 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 5264 6443 5316 6452
rect 5264 6409 5273 6443
rect 5273 6409 5307 6443
rect 5307 6409 5316 6443
rect 5264 6400 5316 6409
rect 8668 6443 8720 6452
rect 8668 6409 8677 6443
rect 8677 6409 8711 6443
rect 8711 6409 8720 6443
rect 8668 6400 8720 6409
rect 10784 6443 10836 6452
rect 10784 6409 10793 6443
rect 10793 6409 10827 6443
rect 10827 6409 10836 6443
rect 10784 6400 10836 6409
rect 12256 6400 12308 6452
rect 16028 6400 16080 6452
rect 18328 6443 18380 6452
rect 18328 6409 18337 6443
rect 18337 6409 18371 6443
rect 18371 6409 18380 6443
rect 18328 6400 18380 6409
rect 20904 6443 20956 6452
rect 20904 6409 20913 6443
rect 20913 6409 20947 6443
rect 20947 6409 20956 6443
rect 20904 6400 20956 6409
rect 23480 6443 23532 6452
rect 23480 6409 23489 6443
rect 23489 6409 23523 6443
rect 23523 6409 23532 6443
rect 23480 6400 23532 6409
rect 25780 6443 25832 6452
rect 25780 6409 25789 6443
rect 25789 6409 25823 6443
rect 25823 6409 25832 6443
rect 25780 6400 25832 6409
rect 36728 6443 36780 6452
rect 36728 6409 36737 6443
rect 36737 6409 36771 6443
rect 36771 6409 36780 6443
rect 36728 6400 36780 6409
rect 49332 6443 49384 6452
rect 3240 6332 3292 6384
rect 4160 6375 4212 6384
rect 4160 6341 4194 6375
rect 4194 6341 4212 6375
rect 4160 6332 4212 6341
rect 8852 6332 8904 6384
rect 1952 6264 2004 6316
rect 3976 6264 4028 6316
rect 7196 6307 7248 6316
rect 7196 6273 7205 6307
rect 7205 6273 7239 6307
rect 7239 6273 7248 6307
rect 11888 6307 11940 6316
rect 7196 6264 7248 6273
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 11888 6264 11940 6273
rect 13544 6332 13596 6384
rect 15844 6332 15896 6384
rect 18696 6332 18748 6384
rect 23848 6332 23900 6384
rect 30288 6332 30340 6384
rect 12440 6264 12492 6316
rect 14740 6307 14792 6316
rect 14740 6273 14749 6307
rect 14749 6273 14783 6307
rect 14783 6273 14792 6307
rect 14740 6264 14792 6273
rect 20628 6264 20680 6316
rect 22008 6264 22060 6316
rect 23204 6264 23256 6316
rect 28908 6264 28960 6316
rect 29644 6264 29696 6316
rect 30932 6264 30984 6316
rect 8944 6196 8996 6248
rect 16304 6196 16356 6248
rect 19432 6196 19484 6248
rect 24308 6196 24360 6248
rect 26976 6239 27028 6248
rect 4068 6060 4120 6112
rect 26976 6205 26985 6239
rect 26985 6205 27019 6239
rect 27019 6205 27028 6239
rect 26976 6196 27028 6205
rect 34060 6332 34112 6384
rect 49332 6409 49341 6443
rect 49341 6409 49375 6443
rect 49375 6409 49384 6443
rect 49332 6400 49384 6409
rect 54668 6443 54720 6452
rect 54668 6409 54677 6443
rect 54677 6409 54711 6443
rect 54711 6409 54720 6443
rect 54668 6400 54720 6409
rect 48964 6332 49016 6384
rect 52184 6332 52236 6384
rect 36728 6264 36780 6316
rect 41696 6264 41748 6316
rect 43076 6264 43128 6316
rect 43904 6264 43956 6316
rect 45376 6264 45428 6316
rect 47400 6264 47452 6316
rect 47492 6264 47544 6316
rect 49792 6307 49844 6316
rect 32128 6239 32180 6248
rect 32128 6205 32137 6239
rect 32137 6205 32171 6239
rect 32171 6205 32180 6239
rect 32128 6196 32180 6205
rect 35348 6239 35400 6248
rect 35348 6205 35357 6239
rect 35357 6205 35391 6239
rect 35391 6205 35400 6239
rect 35348 6196 35400 6205
rect 37740 6196 37792 6248
rect 49792 6273 49801 6307
rect 49801 6273 49835 6307
rect 49835 6273 49844 6307
rect 49792 6264 49844 6273
rect 54116 6264 54168 6316
rect 24676 6060 24728 6112
rect 26056 6060 26108 6112
rect 31116 6103 31168 6112
rect 31116 6069 31125 6103
rect 31125 6069 31159 6103
rect 31159 6069 31168 6103
rect 31116 6060 31168 6069
rect 33508 6103 33560 6112
rect 33508 6069 33517 6103
rect 33517 6069 33551 6103
rect 33551 6069 33560 6103
rect 33508 6060 33560 6069
rect 39396 6103 39448 6112
rect 39396 6069 39405 6103
rect 39405 6069 39439 6103
rect 39439 6069 39448 6103
rect 39396 6060 39448 6069
rect 40224 6060 40276 6112
rect 40592 6060 40644 6112
rect 43352 6060 43404 6112
rect 52736 6196 52788 6248
rect 46848 6060 46900 6112
rect 47032 6103 47084 6112
rect 47032 6069 47041 6103
rect 47041 6069 47075 6103
rect 47075 6069 47084 6103
rect 47032 6060 47084 6069
rect 51172 6103 51224 6112
rect 51172 6069 51181 6103
rect 51181 6069 51215 6103
rect 51215 6069 51224 6103
rect 51172 6060 51224 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 10232 5856 10284 5908
rect 16212 5856 16264 5908
rect 20628 5899 20680 5908
rect 20628 5865 20637 5899
rect 20637 5865 20671 5899
rect 20671 5865 20680 5899
rect 20628 5856 20680 5865
rect 23204 5899 23256 5908
rect 23204 5865 23213 5899
rect 23213 5865 23247 5899
rect 23247 5865 23256 5899
rect 23204 5856 23256 5865
rect 26976 5856 27028 5908
rect 3976 5763 4028 5772
rect 3976 5729 3985 5763
rect 3985 5729 4019 5763
rect 4019 5729 4028 5763
rect 3976 5720 4028 5729
rect 5816 5763 5868 5772
rect 5816 5729 5825 5763
rect 5825 5729 5859 5763
rect 5859 5729 5868 5763
rect 5816 5720 5868 5729
rect 8944 5763 8996 5772
rect 8944 5729 8953 5763
rect 8953 5729 8987 5763
rect 8987 5729 8996 5763
rect 8944 5720 8996 5729
rect 10692 5720 10744 5772
rect 16304 5763 16356 5772
rect 16304 5729 16313 5763
rect 16313 5729 16347 5763
rect 16347 5729 16356 5763
rect 16304 5720 16356 5729
rect 28908 5856 28960 5908
rect 29736 5856 29788 5908
rect 30932 5899 30984 5908
rect 30932 5865 30941 5899
rect 30941 5865 30975 5899
rect 30975 5865 30984 5899
rect 30932 5856 30984 5865
rect 35348 5856 35400 5908
rect 35808 5856 35860 5908
rect 39396 5856 39448 5908
rect 41512 5856 41564 5908
rect 41696 5899 41748 5908
rect 41696 5865 41705 5899
rect 41705 5865 41739 5899
rect 41739 5865 41748 5899
rect 41696 5856 41748 5865
rect 52736 5899 52788 5908
rect 52736 5865 52745 5899
rect 52745 5865 52779 5899
rect 52779 5865 52788 5899
rect 52736 5856 52788 5865
rect 29184 5720 29236 5772
rect 32128 5720 32180 5772
rect 40224 5720 40276 5772
rect 48044 5720 48096 5772
rect 4068 5652 4120 5704
rect 9956 5652 10008 5704
rect 13728 5652 13780 5704
rect 16580 5695 16632 5704
rect 16580 5661 16614 5695
rect 16614 5661 16632 5695
rect 16580 5652 16632 5661
rect 21916 5652 21968 5704
rect 24676 5652 24728 5704
rect 26056 5695 26108 5704
rect 26056 5661 26090 5695
rect 26090 5661 26108 5695
rect 26056 5652 26108 5661
rect 29000 5652 29052 5704
rect 33508 5652 33560 5704
rect 37740 5652 37792 5704
rect 6092 5627 6144 5636
rect 6092 5593 6126 5627
rect 6126 5593 6144 5627
rect 6092 5584 6144 5593
rect 11060 5627 11112 5636
rect 11060 5593 11094 5627
rect 11094 5593 11112 5627
rect 11060 5584 11112 5593
rect 15476 5584 15528 5636
rect 5356 5559 5408 5568
rect 5356 5525 5365 5559
rect 5365 5525 5399 5559
rect 5399 5525 5408 5559
rect 5356 5516 5408 5525
rect 7196 5559 7248 5568
rect 7196 5525 7205 5559
rect 7205 5525 7239 5559
rect 7239 5525 7248 5559
rect 7196 5516 7248 5525
rect 11152 5516 11204 5568
rect 16764 5516 16816 5568
rect 23296 5584 23348 5636
rect 29644 5584 29696 5636
rect 27252 5516 27304 5568
rect 34060 5559 34112 5568
rect 34060 5525 34069 5559
rect 34069 5525 34103 5559
rect 34103 5525 34112 5559
rect 34060 5516 34112 5525
rect 35992 5516 36044 5568
rect 41236 5584 41288 5636
rect 42800 5652 42852 5704
rect 43352 5695 43404 5704
rect 43352 5661 43386 5695
rect 43386 5661 43404 5695
rect 43352 5652 43404 5661
rect 43904 5652 43956 5704
rect 43812 5584 43864 5636
rect 49608 5652 49660 5704
rect 53840 5652 53892 5704
rect 39212 5516 39264 5568
rect 42708 5516 42760 5568
rect 44272 5516 44324 5568
rect 46388 5559 46440 5568
rect 46388 5525 46397 5559
rect 46397 5525 46431 5559
rect 46431 5525 46440 5559
rect 46388 5516 46440 5525
rect 48044 5584 48096 5636
rect 48228 5516 48280 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 11060 5312 11112 5364
rect 7196 5244 7248 5296
rect 10324 5244 10376 5296
rect 12440 5244 12492 5296
rect 25780 5244 25832 5296
rect 29736 5287 29788 5296
rect 29736 5253 29745 5287
rect 29745 5253 29779 5287
rect 29779 5253 29788 5287
rect 29736 5244 29788 5253
rect 34060 5244 34112 5296
rect 44456 5312 44508 5364
rect 45376 5355 45428 5364
rect 45376 5321 45385 5355
rect 45385 5321 45419 5355
rect 45419 5321 45428 5355
rect 45376 5312 45428 5321
rect 39212 5244 39264 5296
rect 39856 5244 39908 5296
rect 46388 5244 46440 5296
rect 54116 5312 54168 5364
rect 51172 5244 51224 5296
rect 1952 5176 2004 5228
rect 5356 5176 5408 5228
rect 5816 5176 5868 5228
rect 8944 5176 8996 5228
rect 9772 5176 9824 5228
rect 14740 5176 14792 5228
rect 18604 5176 18656 5228
rect 32588 5176 32640 5228
rect 39488 5176 39540 5228
rect 43904 5176 43956 5228
rect 52644 5176 52696 5228
rect 54024 5176 54076 5228
rect 3976 5108 4028 5160
rect 4068 4972 4120 5024
rect 7380 4972 7432 5024
rect 10692 4972 10744 5024
rect 13728 5108 13780 5160
rect 13820 4972 13872 5024
rect 34612 5108 34664 5160
rect 37740 5151 37792 5160
rect 37740 5117 37749 5151
rect 37749 5117 37783 5151
rect 37783 5117 37792 5151
rect 37740 5108 37792 5117
rect 41696 5108 41748 5160
rect 50160 5151 50212 5160
rect 50160 5117 50169 5151
rect 50169 5117 50203 5151
rect 50203 5117 50212 5151
rect 50160 5108 50212 5117
rect 22008 5040 22060 5092
rect 22744 4972 22796 5024
rect 24032 4972 24084 5024
rect 24676 5015 24728 5024
rect 24676 4981 24685 5015
rect 24685 4981 24719 5015
rect 24719 4981 24728 5015
rect 24676 4972 24728 4981
rect 33876 5015 33928 5024
rect 33876 4981 33885 5015
rect 33885 4981 33919 5015
rect 33919 4981 33928 5015
rect 33876 4972 33928 4981
rect 36544 5015 36596 5024
rect 36544 4981 36553 5015
rect 36553 4981 36587 5015
rect 36587 4981 36596 5015
rect 36544 4972 36596 4981
rect 39948 4972 40000 5024
rect 50436 4972 50488 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 15476 4811 15528 4820
rect 15476 4777 15485 4811
rect 15485 4777 15519 4811
rect 15519 4777 15528 4811
rect 15476 4768 15528 4777
rect 9772 4675 9824 4684
rect 9772 4641 9781 4675
rect 9781 4641 9815 4675
rect 9815 4641 9824 4675
rect 9772 4632 9824 4641
rect 10784 4632 10836 4684
rect 16304 4768 16356 4820
rect 22100 4768 22152 4820
rect 23296 4811 23348 4820
rect 23296 4777 23305 4811
rect 23305 4777 23339 4811
rect 23339 4777 23348 4811
rect 23296 4768 23348 4777
rect 36728 4811 36780 4820
rect 36728 4777 36737 4811
rect 36737 4777 36771 4811
rect 36771 4777 36780 4811
rect 36728 4768 36780 4777
rect 41236 4811 41288 4820
rect 41236 4777 41245 4811
rect 41245 4777 41279 4811
rect 41279 4777 41288 4811
rect 41236 4768 41288 4777
rect 47400 4768 47452 4820
rect 26976 4675 27028 4684
rect 26976 4641 26985 4675
rect 26985 4641 27019 4675
rect 27019 4641 27028 4675
rect 26976 4632 27028 4641
rect 29184 4632 29236 4684
rect 4068 4607 4120 4616
rect 4068 4573 4102 4607
rect 4102 4573 4120 4607
rect 4068 4564 4120 4573
rect 5724 4564 5776 4616
rect 11152 4564 11204 4616
rect 13360 4564 13412 4616
rect 19432 4564 19484 4616
rect 20628 4564 20680 4616
rect 22008 4564 22060 4616
rect 27252 4607 27304 4616
rect 27252 4573 27286 4607
rect 27286 4573 27304 4607
rect 27252 4564 27304 4573
rect 31116 4564 31168 4616
rect 32588 4564 32640 4616
rect 33876 4564 33928 4616
rect 34612 4564 34664 4616
rect 5540 4496 5592 4548
rect 5172 4471 5224 4480
rect 5172 4437 5181 4471
rect 5181 4437 5215 4471
rect 5215 4437 5224 4471
rect 5172 4428 5224 4437
rect 6000 4428 6052 4480
rect 15476 4496 15528 4548
rect 17132 4496 17184 4548
rect 21824 4496 21876 4548
rect 23204 4496 23256 4548
rect 36544 4564 36596 4616
rect 39856 4607 39908 4616
rect 11244 4428 11296 4480
rect 17316 4471 17368 4480
rect 17316 4437 17325 4471
rect 17325 4437 17359 4471
rect 17359 4437 17368 4471
rect 17316 4428 17368 4437
rect 26516 4471 26568 4480
rect 26516 4437 26525 4471
rect 26525 4437 26559 4471
rect 26559 4437 26568 4471
rect 26516 4428 26568 4437
rect 35808 4496 35860 4548
rect 38844 4496 38896 4548
rect 39856 4573 39865 4607
rect 39865 4573 39899 4607
rect 39899 4573 39908 4607
rect 39856 4564 39908 4573
rect 39948 4564 40000 4616
rect 41696 4607 41748 4616
rect 41696 4573 41705 4607
rect 41705 4573 41739 4607
rect 41739 4573 41748 4607
rect 41696 4564 41748 4573
rect 42432 4564 42484 4616
rect 41512 4496 41564 4548
rect 47676 4564 47728 4616
rect 50160 4607 50212 4616
rect 50160 4573 50169 4607
rect 50169 4573 50203 4607
rect 50203 4573 50212 4607
rect 50160 4564 50212 4573
rect 50436 4607 50488 4616
rect 50436 4573 50470 4607
rect 50470 4573 50488 4607
rect 50436 4564 50488 4573
rect 52736 4564 52788 4616
rect 48228 4496 48280 4548
rect 53564 4496 53616 4548
rect 31392 4471 31444 4480
rect 31392 4437 31401 4471
rect 31401 4437 31435 4471
rect 31435 4437 31444 4471
rect 31392 4428 31444 4437
rect 34152 4471 34204 4480
rect 34152 4437 34161 4471
rect 34161 4437 34195 4471
rect 34195 4437 34204 4471
rect 34152 4428 34204 4437
rect 38568 4471 38620 4480
rect 38568 4437 38577 4471
rect 38577 4437 38611 4471
rect 38611 4437 38620 4471
rect 38568 4428 38620 4437
rect 43076 4471 43128 4480
rect 43076 4437 43085 4471
rect 43085 4437 43119 4471
rect 43119 4437 43128 4471
rect 43076 4428 43128 4437
rect 51540 4471 51592 4480
rect 51540 4437 51549 4471
rect 51549 4437 51583 4471
rect 51583 4437 51592 4471
rect 51540 4428 51592 4437
rect 53380 4471 53432 4480
rect 53380 4437 53389 4471
rect 53389 4437 53423 4471
rect 53423 4437 53432 4471
rect 53380 4428 53432 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 3976 4224 4028 4276
rect 14740 4267 14792 4276
rect 14740 4233 14749 4267
rect 14749 4233 14783 4267
rect 14783 4233 14792 4267
rect 14740 4224 14792 4233
rect 23204 4267 23256 4276
rect 23204 4233 23213 4267
rect 23213 4233 23247 4267
rect 23247 4233 23256 4267
rect 23204 4224 23256 4233
rect 18604 4199 18656 4208
rect 18604 4165 18613 4199
rect 18613 4165 18647 4199
rect 18647 4165 18656 4199
rect 18604 4156 18656 4165
rect 5172 4088 5224 4140
rect 5724 4088 5776 4140
rect 7380 4088 7432 4140
rect 10784 4088 10836 4140
rect 11796 4131 11848 4140
rect 11796 4097 11830 4131
rect 11830 4097 11848 4131
rect 11796 4088 11848 4097
rect 13084 4088 13136 4140
rect 16304 4088 16356 4140
rect 16764 4088 16816 4140
rect 22008 4156 22060 4208
rect 26516 4156 26568 4208
rect 37740 4156 37792 4208
rect 22100 4131 22152 4140
rect 22100 4097 22134 4131
rect 22134 4097 22152 4131
rect 22100 4088 22152 4097
rect 25688 4088 25740 4140
rect 26976 4131 27028 4140
rect 26976 4097 26985 4131
rect 26985 4097 27019 4131
rect 27019 4097 27028 4131
rect 26976 4088 27028 4097
rect 31392 4088 31444 4140
rect 34152 4088 34204 4140
rect 13360 4063 13412 4072
rect 13360 4029 13369 4063
rect 13369 4029 13403 4063
rect 13403 4029 13412 4063
rect 13360 4020 13412 4029
rect 20628 4020 20680 4072
rect 24032 4063 24084 4072
rect 24032 4029 24041 4063
rect 24041 4029 24075 4063
rect 24075 4029 24084 4063
rect 24032 4020 24084 4029
rect 5540 3952 5592 4004
rect 7748 3995 7800 4004
rect 7748 3961 7757 3995
rect 7757 3961 7791 3995
rect 7791 3961 7800 3995
rect 7748 3952 7800 3961
rect 12900 3927 12952 3936
rect 12900 3893 12909 3927
rect 12909 3893 12943 3927
rect 12943 3893 12952 3927
rect 12900 3884 12952 3893
rect 18052 3927 18104 3936
rect 18052 3893 18061 3927
rect 18061 3893 18095 3927
rect 18095 3893 18104 3927
rect 18052 3884 18104 3893
rect 25412 3927 25464 3936
rect 25412 3893 25421 3927
rect 25421 3893 25455 3927
rect 25455 3893 25464 3927
rect 25412 3884 25464 3893
rect 28356 3927 28408 3936
rect 28356 3893 28365 3927
rect 28365 3893 28399 3927
rect 28399 3893 28408 3927
rect 28356 3884 28408 3893
rect 32588 4020 32640 4072
rect 37280 4131 37332 4140
rect 37280 4097 37289 4131
rect 37289 4097 37323 4131
rect 37323 4097 37332 4131
rect 37280 4088 37332 4097
rect 38752 4088 38804 4140
rect 39856 4156 39908 4208
rect 53380 4156 53432 4208
rect 40408 4088 40460 4140
rect 44272 4131 44324 4140
rect 44272 4097 44306 4131
rect 44306 4097 44324 4131
rect 44272 4088 44324 4097
rect 47032 4088 47084 4140
rect 49976 4088 50028 4140
rect 51540 4088 51592 4140
rect 52736 4131 52788 4140
rect 52736 4097 52745 4131
rect 52745 4097 52779 4131
rect 52779 4097 52788 4131
rect 52736 4088 52788 4097
rect 34612 4063 34664 4072
rect 34612 4029 34621 4063
rect 34621 4029 34655 4063
rect 34655 4029 34664 4063
rect 34612 4020 34664 4029
rect 42432 4020 42484 4072
rect 46940 4020 46992 4072
rect 35992 3995 36044 4004
rect 35992 3961 36001 3995
rect 36001 3961 36035 3995
rect 36035 3961 36044 3995
rect 35992 3952 36044 3961
rect 45284 3952 45336 4004
rect 31116 3927 31168 3936
rect 31116 3893 31125 3927
rect 31125 3893 31159 3927
rect 31159 3893 31168 3927
rect 31116 3884 31168 3893
rect 38660 3927 38712 3936
rect 38660 3893 38669 3927
rect 38669 3893 38703 3927
rect 38703 3893 38712 3927
rect 38660 3884 38712 3893
rect 40500 3927 40552 3936
rect 40500 3893 40509 3927
rect 40509 3893 40543 3927
rect 40543 3893 40552 3927
rect 40500 3884 40552 3893
rect 48964 3927 49016 3936
rect 48964 3893 48973 3927
rect 48973 3893 49007 3927
rect 49007 3893 49016 3927
rect 48964 3884 49016 3893
rect 50620 3884 50672 3936
rect 54116 3927 54168 3936
rect 54116 3893 54125 3927
rect 54125 3893 54159 3927
rect 54159 3893 54168 3927
rect 54116 3884 54168 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 5724 3680 5776 3732
rect 6092 3680 6144 3732
rect 10784 3680 10836 3732
rect 11796 3723 11848 3732
rect 11796 3689 11805 3723
rect 11805 3689 11839 3723
rect 11839 3689 11848 3723
rect 11796 3680 11848 3689
rect 15476 3723 15528 3732
rect 15476 3689 15485 3723
rect 15485 3689 15519 3723
rect 15519 3689 15528 3723
rect 15476 3680 15528 3689
rect 13360 3544 13412 3596
rect 16304 3680 16356 3732
rect 17132 3680 17184 3732
rect 21824 3680 21876 3732
rect 26976 3680 27028 3732
rect 31024 3723 31076 3732
rect 31024 3689 31033 3723
rect 31033 3689 31067 3723
rect 31067 3689 31076 3723
rect 31024 3680 31076 3689
rect 39488 3680 39540 3732
rect 32588 3587 32640 3596
rect 6000 3476 6052 3528
rect 11244 3476 11296 3528
rect 18052 3476 18104 3528
rect 19340 3476 19392 3528
rect 20628 3476 20680 3528
rect 32588 3553 32597 3587
rect 32597 3553 32631 3587
rect 32631 3553 32640 3587
rect 32588 3544 32640 3553
rect 34612 3544 34664 3596
rect 39856 3587 39908 3596
rect 28356 3476 28408 3528
rect 29736 3476 29788 3528
rect 31116 3476 31168 3528
rect 39856 3553 39865 3587
rect 39865 3553 39899 3587
rect 39899 3553 39908 3587
rect 39856 3544 39908 3553
rect 42800 3680 42852 3732
rect 43812 3723 43864 3732
rect 43812 3689 43821 3723
rect 43821 3689 43855 3723
rect 43855 3689 43864 3723
rect 43812 3680 43864 3689
rect 49608 3723 49660 3732
rect 49608 3689 49617 3723
rect 49617 3689 49651 3723
rect 49651 3689 49660 3723
rect 49608 3680 49660 3689
rect 53564 3723 53616 3732
rect 53564 3689 53573 3723
rect 53573 3689 53607 3723
rect 53607 3689 53616 3723
rect 53564 3680 53616 3689
rect 40500 3476 40552 3528
rect 43076 3476 43128 3528
rect 48228 3519 48280 3528
rect 48228 3485 48237 3519
rect 48237 3485 48271 3519
rect 48271 3485 48280 3519
rect 48228 3476 48280 3485
rect 48964 3476 49016 3528
rect 50160 3476 50212 3528
rect 50620 3519 50672 3528
rect 50620 3485 50654 3519
rect 50654 3485 50672 3519
rect 14740 3408 14792 3460
rect 18144 3408 18196 3460
rect 23204 3408 23256 3460
rect 27344 3408 27396 3460
rect 33508 3408 33560 3460
rect 34060 3408 34112 3460
rect 35900 3408 35952 3460
rect 50620 3476 50672 3485
rect 52736 3476 52788 3528
rect 52276 3408 52328 3460
rect 18052 3340 18104 3392
rect 26240 3383 26292 3392
rect 26240 3349 26249 3383
rect 26249 3349 26283 3383
rect 26283 3349 26292 3383
rect 28080 3383 28132 3392
rect 26240 3340 26292 3349
rect 28080 3349 28089 3383
rect 28089 3349 28123 3383
rect 28123 3349 28132 3383
rect 28080 3340 28132 3349
rect 33968 3383 34020 3392
rect 33968 3349 33977 3383
rect 33977 3349 34011 3383
rect 34011 3349 34020 3383
rect 33968 3340 34020 3349
rect 36084 3383 36136 3392
rect 36084 3349 36093 3383
rect 36093 3349 36127 3383
rect 36127 3349 36136 3383
rect 36084 3340 36136 3349
rect 36452 3340 36504 3392
rect 51724 3383 51776 3392
rect 51724 3349 51733 3383
rect 51733 3349 51767 3383
rect 51767 3349 51776 3383
rect 51724 3340 51776 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 14740 3179 14792 3188
rect 14740 3145 14749 3179
rect 14749 3145 14783 3179
rect 14783 3145 14792 3179
rect 14740 3136 14792 3145
rect 18144 3136 18196 3188
rect 25688 3179 25740 3188
rect 12900 3068 12952 3120
rect 13820 3068 13872 3120
rect 17316 3068 17368 3120
rect 10784 3000 10836 3052
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 13360 3043 13412 3052
rect 11520 3000 11572 3009
rect 13360 3009 13369 3043
rect 13369 3009 13403 3043
rect 13403 3009 13412 3043
rect 13360 3000 13412 3009
rect 16304 3000 16356 3052
rect 17224 3000 17276 3052
rect 19340 3068 19392 3120
rect 22744 3111 22796 3120
rect 22744 3077 22778 3111
rect 22778 3077 22796 3111
rect 22744 3068 22796 3077
rect 18604 3000 18656 3052
rect 25688 3145 25697 3179
rect 25697 3145 25731 3179
rect 25731 3145 25740 3179
rect 25688 3136 25740 3145
rect 29644 3136 29696 3188
rect 34060 3179 34112 3188
rect 34060 3145 34069 3179
rect 34069 3145 34103 3179
rect 34103 3145 34112 3179
rect 34060 3136 34112 3145
rect 35900 3179 35952 3188
rect 35900 3145 35909 3179
rect 35909 3145 35943 3179
rect 35943 3145 35952 3179
rect 35900 3136 35952 3145
rect 40408 3136 40460 3188
rect 43536 3136 43588 3188
rect 52276 3136 52328 3188
rect 26240 3068 26292 3120
rect 28080 3068 28132 3120
rect 33968 3068 34020 3120
rect 36084 3068 36136 3120
rect 38660 3068 38712 3120
rect 42708 3111 42760 3120
rect 42708 3077 42742 3111
rect 42742 3077 42760 3111
rect 42708 3068 42760 3077
rect 51724 3068 51776 3120
rect 54116 3068 54168 3120
rect 32588 3000 32640 3052
rect 34612 3000 34664 3052
rect 37280 3043 37332 3052
rect 37280 3009 37289 3043
rect 37289 3009 37323 3043
rect 37323 3009 37332 3043
rect 37280 3000 37332 3009
rect 37556 3043 37608 3052
rect 37556 3009 37590 3043
rect 37590 3009 37608 3043
rect 37556 3000 37608 3009
rect 39856 3000 39908 3052
rect 42432 3043 42484 3052
rect 42432 3009 42441 3043
rect 42441 3009 42475 3043
rect 42475 3009 42484 3043
rect 42432 3000 42484 3009
rect 48228 3000 48280 3052
rect 52736 3043 52788 3052
rect 52736 3009 52745 3043
rect 52745 3009 52779 3043
rect 52779 3009 52788 3043
rect 52736 3000 52788 3009
rect 24032 2932 24084 2984
rect 26976 2975 27028 2984
rect 26976 2941 26985 2975
rect 26985 2941 27019 2975
rect 27019 2941 27028 2975
rect 26976 2932 27028 2941
rect 12900 2839 12952 2848
rect 12900 2805 12909 2839
rect 12909 2805 12943 2839
rect 12943 2805 12952 2839
rect 12900 2796 12952 2805
rect 19984 2796 20036 2848
rect 24308 2796 24360 2848
rect 38844 2864 38896 2916
rect 54024 2864 54076 2916
rect 28356 2839 28408 2848
rect 28356 2805 28365 2839
rect 28365 2805 28399 2839
rect 28399 2805 28408 2839
rect 28356 2796 28408 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 18604 2635 18656 2644
rect 13084 2567 13136 2576
rect 13084 2533 13093 2567
rect 13093 2533 13127 2567
rect 13127 2533 13136 2567
rect 13084 2524 13136 2533
rect 18604 2601 18613 2635
rect 18613 2601 18647 2635
rect 18647 2601 18656 2635
rect 18604 2592 18656 2601
rect 23204 2635 23256 2644
rect 11520 2456 11572 2508
rect 17224 2499 17276 2508
rect 17224 2465 17233 2499
rect 17233 2465 17267 2499
rect 17267 2465 17276 2499
rect 17224 2456 17276 2465
rect 12900 2388 12952 2440
rect 18052 2388 18104 2440
rect 20 2320 72 2372
rect 19984 2388 20036 2440
rect 20628 2388 20680 2440
rect 23204 2601 23213 2635
rect 23213 2601 23247 2635
rect 23247 2601 23256 2635
rect 23204 2592 23256 2601
rect 25780 2635 25832 2644
rect 25780 2601 25789 2635
rect 25789 2601 25823 2635
rect 25823 2601 25832 2635
rect 25780 2592 25832 2601
rect 27344 2592 27396 2644
rect 33508 2592 33560 2644
rect 37556 2592 37608 2644
rect 38752 2592 38804 2644
rect 24308 2456 24360 2508
rect 26976 2499 27028 2508
rect 26976 2465 26985 2499
rect 26985 2465 27019 2499
rect 27019 2465 27028 2499
rect 26976 2456 27028 2465
rect 34612 2456 34664 2508
rect 37280 2499 37332 2508
rect 37280 2465 37289 2499
rect 37289 2465 37323 2499
rect 37323 2465 37332 2499
rect 37280 2456 37332 2465
rect 25412 2388 25464 2440
rect 28356 2388 28408 2440
rect 34244 2388 34296 2440
rect 36452 2388 36504 2440
rect 38568 2388 38620 2440
rect 28540 2320 28592 2372
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
<< metal2 >>
rect 26146 61860 26202 62660
rect 60370 61860 60426 62660
rect 4214 60412 4522 60432
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60336 4522 60356
rect 26160 60330 26188 61860
rect 34934 60412 35242 60432
rect 34934 60410 34940 60412
rect 34996 60410 35020 60412
rect 35076 60410 35100 60412
rect 35156 60410 35180 60412
rect 35236 60410 35242 60412
rect 34996 60358 34998 60410
rect 35178 60358 35180 60410
rect 34934 60356 34940 60358
rect 34996 60356 35020 60358
rect 35076 60356 35100 60358
rect 35156 60356 35180 60358
rect 35236 60356 35242 60358
rect 34934 60336 35242 60356
rect 26160 60302 26280 60330
rect 26252 60246 26280 60302
rect 60384 60246 60412 61860
rect 26240 60240 26292 60246
rect 26240 60182 26292 60188
rect 60372 60240 60424 60246
rect 60372 60182 60424 60188
rect 11520 60104 11572 60110
rect 11520 60046 11572 60052
rect 29920 60104 29972 60110
rect 29920 60046 29972 60052
rect 32128 60104 32180 60110
rect 32128 60046 32180 60052
rect 34060 60104 34112 60110
rect 34060 60046 34112 60052
rect 37556 60104 37608 60110
rect 37556 60046 37608 60052
rect 40408 60104 40460 60110
rect 40408 60046 40460 60052
rect 43628 60104 43680 60110
rect 43628 60046 43680 60052
rect 45560 60104 45612 60110
rect 45560 60046 45612 60052
rect 48964 60104 49016 60110
rect 48964 60046 49016 60052
rect 50804 60104 50856 60110
rect 50804 60046 50856 60052
rect 54116 60104 54168 60110
rect 54116 60046 54168 60052
rect 7748 60036 7800 60042
rect 7748 59978 7800 59984
rect 6920 59968 6972 59974
rect 6920 59910 6972 59916
rect 6932 59702 6960 59910
rect 7760 59770 7788 59978
rect 8484 59968 8536 59974
rect 8484 59910 8536 59916
rect 7748 59764 7800 59770
rect 7748 59706 7800 59712
rect 6920 59696 6972 59702
rect 6920 59638 6972 59644
rect 4214 59324 4522 59344
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 4214 59248 4522 59268
rect 6184 59016 6236 59022
rect 6184 58958 6236 58964
rect 6828 59016 6880 59022
rect 6932 58970 6960 59638
rect 8116 59628 8168 59634
rect 8116 59570 8168 59576
rect 8128 59226 8156 59570
rect 8116 59220 8168 59226
rect 8116 59162 8168 59168
rect 6880 58964 6960 58970
rect 6828 58958 6960 58964
rect 8208 59016 8260 59022
rect 8208 58958 8260 58964
rect 6000 58948 6052 58954
rect 6000 58890 6052 58896
rect 5172 58540 5224 58546
rect 5172 58482 5224 58488
rect 4214 58236 4522 58256
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58160 4522 58180
rect 5184 58138 5212 58482
rect 5540 58336 5592 58342
rect 5540 58278 5592 58284
rect 5172 58132 5224 58138
rect 5172 58074 5224 58080
rect 3884 57928 3936 57934
rect 3884 57870 3936 57876
rect 3896 57254 3924 57870
rect 5552 57866 5580 58278
rect 4988 57860 5040 57866
rect 4988 57802 5040 57808
rect 5540 57860 5592 57866
rect 5540 57802 5592 57808
rect 5000 57594 5028 57802
rect 6012 57798 6040 58890
rect 6196 58614 6224 58958
rect 6840 58942 6960 58958
rect 6276 58880 6328 58886
rect 6276 58822 6328 58828
rect 6288 58614 6316 58822
rect 6184 58608 6236 58614
rect 6184 58550 6236 58556
rect 6276 58608 6328 58614
rect 6276 58550 6328 58556
rect 6196 58426 6224 58550
rect 6932 58546 6960 58942
rect 7748 58948 7800 58954
rect 7748 58890 7800 58896
rect 7760 58682 7788 58890
rect 7748 58676 7800 58682
rect 7748 58618 7800 58624
rect 8220 58546 8248 58958
rect 8496 58614 8524 59910
rect 9496 59628 9548 59634
rect 9496 59570 9548 59576
rect 9508 58682 9536 59570
rect 11532 59566 11560 60046
rect 12900 60036 12952 60042
rect 12900 59978 12952 59984
rect 28448 60036 28500 60042
rect 28448 59978 28500 59984
rect 12912 59770 12940 59978
rect 13084 59968 13136 59974
rect 13084 59910 13136 59916
rect 12900 59764 12952 59770
rect 12900 59706 12952 59712
rect 12256 59628 12308 59634
rect 12256 59570 12308 59576
rect 11520 59560 11572 59566
rect 11520 59502 11572 59508
rect 9588 59424 9640 59430
rect 9588 59366 9640 59372
rect 9600 59022 9628 59366
rect 11532 59022 11560 59502
rect 9588 59016 9640 59022
rect 9588 58958 9640 58964
rect 11520 59016 11572 59022
rect 11520 58958 11572 58964
rect 10324 58880 10376 58886
rect 10324 58822 10376 58828
rect 9496 58676 9548 58682
rect 9496 58618 9548 58624
rect 8484 58608 8536 58614
rect 8484 58550 8536 58556
rect 6920 58540 6972 58546
rect 6920 58482 6972 58488
rect 8208 58540 8260 58546
rect 8208 58482 8260 58488
rect 6276 58472 6328 58478
rect 6196 58420 6276 58426
rect 6196 58414 6328 58420
rect 6196 58398 6316 58414
rect 6000 57792 6052 57798
rect 6000 57734 6052 57740
rect 4988 57588 5040 57594
rect 4988 57530 5040 57536
rect 5172 57452 5224 57458
rect 5172 57394 5224 57400
rect 3884 57248 3936 57254
rect 3884 57190 3936 57196
rect 3896 56846 3924 57190
rect 4214 57148 4522 57168
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57072 4522 57092
rect 5184 57050 5212 57394
rect 5172 57044 5224 57050
rect 5172 56986 5224 56992
rect 3884 56840 3936 56846
rect 3884 56782 3936 56788
rect 3896 56166 3924 56782
rect 4988 56772 5040 56778
rect 4988 56714 5040 56720
rect 5000 56506 5028 56714
rect 4988 56500 5040 56506
rect 4988 56442 5040 56448
rect 5172 56364 5224 56370
rect 5172 56306 5224 56312
rect 3884 56160 3936 56166
rect 3884 56102 3936 56108
rect 3896 55282 3924 56102
rect 4214 56060 4522 56080
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55984 4522 56004
rect 5184 55418 5212 56306
rect 5540 55684 5592 55690
rect 5540 55626 5592 55632
rect 5172 55412 5224 55418
rect 5172 55354 5224 55360
rect 3884 55276 3936 55282
rect 3884 55218 3936 55224
rect 3896 54670 3924 55218
rect 4214 54972 4522 54992
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54896 4522 54916
rect 3884 54664 3936 54670
rect 3884 54606 3936 54612
rect 2872 54120 2924 54126
rect 2872 54062 2924 54068
rect 2884 53650 2912 54062
rect 3896 53938 3924 54606
rect 5356 54188 5408 54194
rect 5356 54130 5408 54136
rect 3804 53910 3924 53938
rect 4620 53984 4672 53990
rect 4620 53926 4672 53932
rect 3804 53650 3832 53910
rect 4214 53884 4522 53904
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53808 4522 53828
rect 2872 53644 2924 53650
rect 2872 53586 2924 53592
rect 3792 53644 3844 53650
rect 3792 53586 3844 53592
rect 2884 53174 2912 53586
rect 4632 53582 4660 53926
rect 4620 53576 4672 53582
rect 4620 53518 4672 53524
rect 5368 53242 5396 54130
rect 5356 53236 5408 53242
rect 5356 53178 5408 53184
rect 2872 53168 2924 53174
rect 2872 53110 2924 53116
rect 3240 53100 3292 53106
rect 3240 53042 3292 53048
rect 3252 52698 3280 53042
rect 4214 52796 4522 52816
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52720 4522 52740
rect 3240 52692 3292 52698
rect 3240 52634 3292 52640
rect 1584 52488 1636 52494
rect 1584 52430 1636 52436
rect 3424 52488 3476 52494
rect 3424 52430 3476 52436
rect 1596 51950 1624 52430
rect 3436 52154 3464 52430
rect 4620 52420 4672 52426
rect 4620 52362 4672 52368
rect 3424 52148 3476 52154
rect 3424 52090 3476 52096
rect 3240 52012 3292 52018
rect 3240 51954 3292 51960
rect 1584 51944 1636 51950
rect 1584 51886 1636 51892
rect 1596 51406 1624 51886
rect 3252 51610 3280 51954
rect 4214 51708 4522 51728
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51632 4522 51652
rect 3240 51604 3292 51610
rect 3240 51546 3292 51552
rect 1584 51400 1636 51406
rect 1584 51342 1636 51348
rect 4436 51400 4488 51406
rect 4632 51388 4660 52362
rect 4488 51360 4660 51388
rect 5172 51400 5224 51406
rect 4436 51342 4488 51348
rect 5172 51342 5224 51348
rect 1596 50862 1624 51342
rect 3424 51332 3476 51338
rect 3424 51274 3476 51280
rect 3436 51066 3464 51274
rect 3424 51060 3476 51066
rect 3424 51002 3476 51008
rect 4448 50930 4476 51342
rect 3240 50924 3292 50930
rect 3240 50866 3292 50872
rect 4436 50924 4488 50930
rect 4436 50866 4488 50872
rect 1584 50856 1636 50862
rect 1584 50798 1636 50804
rect 1596 50318 1624 50798
rect 3252 50522 3280 50866
rect 3698 50688 3754 50697
rect 3698 50623 3754 50632
rect 3240 50516 3292 50522
rect 3240 50458 3292 50464
rect 1584 50312 1636 50318
rect 1584 50254 1636 50260
rect 1596 49774 1624 50254
rect 2872 50244 2924 50250
rect 2872 50186 2924 50192
rect 1584 49768 1636 49774
rect 1584 49710 1636 49716
rect 1596 49230 1624 49710
rect 2884 49434 2912 50186
rect 3516 49836 3568 49842
rect 3516 49778 3568 49784
rect 2964 49632 3016 49638
rect 2964 49574 3016 49580
rect 2872 49428 2924 49434
rect 2872 49370 2924 49376
rect 2976 49230 3004 49574
rect 1584 49224 1636 49230
rect 1584 49166 1636 49172
rect 2964 49224 3016 49230
rect 2964 49166 3016 49172
rect 1860 49088 1912 49094
rect 1860 49030 1912 49036
rect 1872 48550 1900 49030
rect 3528 48890 3556 49778
rect 3516 48884 3568 48890
rect 3516 48826 3568 48832
rect 1860 48544 1912 48550
rect 1860 48486 1912 48492
rect 1872 46510 1900 48486
rect 3240 46572 3292 46578
rect 3240 46514 3292 46520
rect 1860 46504 1912 46510
rect 1860 46446 1912 46452
rect 1872 46034 1900 46446
rect 3252 46170 3280 46514
rect 3240 46164 3292 46170
rect 3240 46106 3292 46112
rect 1860 46028 1912 46034
rect 1860 45970 1912 45976
rect 3148 45484 3200 45490
rect 3148 45426 3200 45432
rect 1676 45416 1728 45422
rect 1676 45358 1728 45364
rect 1688 44878 1716 45358
rect 3160 45082 3188 45426
rect 3148 45076 3200 45082
rect 3148 45018 3200 45024
rect 1676 44872 1728 44878
rect 1676 44814 1728 44820
rect 1688 44402 1716 44814
rect 3056 44804 3108 44810
rect 3056 44746 3108 44752
rect 3068 44538 3096 44746
rect 3056 44532 3108 44538
rect 3056 44474 3108 44480
rect 1676 44396 1728 44402
rect 1676 44338 1728 44344
rect 3056 44396 3108 44402
rect 3056 44338 3108 44344
rect 1688 43858 1716 44338
rect 1676 43852 1728 43858
rect 1676 43794 1728 43800
rect 1688 43314 1716 43794
rect 3068 43450 3096 44338
rect 3240 43648 3292 43654
rect 3240 43590 3292 43596
rect 3056 43444 3108 43450
rect 3056 43386 3108 43392
rect 3252 43382 3280 43590
rect 3240 43376 3292 43382
rect 3240 43318 3292 43324
rect 1676 43308 1728 43314
rect 1676 43250 1728 43256
rect 3240 41132 3292 41138
rect 3240 41074 3292 41080
rect 3252 40730 3280 41074
rect 3240 40724 3292 40730
rect 3240 40666 3292 40672
rect 2872 40520 2924 40526
rect 2872 40462 2924 40468
rect 2884 40118 2912 40462
rect 3240 40452 3292 40458
rect 3240 40394 3292 40400
rect 2872 40112 2924 40118
rect 2872 40054 2924 40060
rect 3252 39642 3280 40394
rect 3608 39840 3660 39846
rect 3608 39782 3660 39788
rect 3240 39636 3292 39642
rect 3240 39578 3292 39584
rect 3620 39438 3648 39782
rect 3608 39432 3660 39438
rect 3608 39374 3660 39380
rect 3332 32904 3384 32910
rect 3332 32846 3384 32852
rect 3344 32434 3372 32846
rect 3332 32428 3384 32434
rect 3332 32370 3384 32376
rect 2872 31816 2924 31822
rect 2872 31758 2924 31764
rect 2884 31346 2912 31758
rect 3712 31414 3740 50623
rect 4214 50620 4522 50640
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50544 4522 50564
rect 5184 50522 5212 51342
rect 5172 50516 5224 50522
rect 5172 50458 5224 50464
rect 5552 50318 5580 55626
rect 6288 55622 6316 58398
rect 6932 57934 6960 58482
rect 10336 57934 10364 58822
rect 11532 58478 11560 58958
rect 12164 58880 12216 58886
rect 12164 58822 12216 58828
rect 12176 58614 12204 58822
rect 12164 58608 12216 58614
rect 12164 58550 12216 58556
rect 11520 58472 11572 58478
rect 11520 58414 11572 58420
rect 6920 57928 6972 57934
rect 6920 57870 6972 57876
rect 10324 57928 10376 57934
rect 10324 57870 10376 57876
rect 10784 57928 10836 57934
rect 10784 57870 10836 57876
rect 6932 57390 6960 57870
rect 10796 57798 10824 57870
rect 8944 57792 8996 57798
rect 8944 57734 8996 57740
rect 10784 57792 10836 57798
rect 10784 57734 10836 57740
rect 8300 57452 8352 57458
rect 8300 57394 8352 57400
rect 8760 57452 8812 57458
rect 8760 57394 8812 57400
rect 6920 57384 6972 57390
rect 6920 57326 6972 57332
rect 6932 56846 6960 57326
rect 8312 57050 8340 57394
rect 8392 57248 8444 57254
rect 8392 57190 8444 57196
rect 8300 57044 8352 57050
rect 8300 56986 8352 56992
rect 6920 56840 6972 56846
rect 6920 56782 6972 56788
rect 8300 56840 8352 56846
rect 8300 56782 8352 56788
rect 6932 56302 6960 56782
rect 8312 56506 8340 56782
rect 8300 56500 8352 56506
rect 8300 56442 8352 56448
rect 8208 56364 8260 56370
rect 8208 56306 8260 56312
rect 6920 56296 6972 56302
rect 6920 56238 6972 56244
rect 6276 55616 6328 55622
rect 6276 55558 6328 55564
rect 6288 54670 6316 55558
rect 6932 55282 6960 56238
rect 8220 55418 8248 56306
rect 8208 55412 8260 55418
rect 8208 55354 8260 55360
rect 8404 55350 8432 57190
rect 8772 55690 8800 57394
rect 8956 56914 8984 57734
rect 10796 57390 10824 57734
rect 10784 57384 10836 57390
rect 10784 57326 10836 57332
rect 8944 56908 8996 56914
rect 8944 56850 8996 56856
rect 8956 56506 8984 56850
rect 11532 56846 11560 58414
rect 12164 57792 12216 57798
rect 12164 57734 12216 57740
rect 12176 57526 12204 57734
rect 12164 57520 12216 57526
rect 12164 57462 12216 57468
rect 12268 57050 12296 59570
rect 12808 58948 12860 58954
rect 12808 58890 12860 58896
rect 12820 57594 12848 58890
rect 13096 58614 13124 59910
rect 19574 59868 19882 59888
rect 19574 59866 19580 59868
rect 19636 59866 19660 59868
rect 19716 59866 19740 59868
rect 19796 59866 19820 59868
rect 19876 59866 19882 59868
rect 19636 59814 19638 59866
rect 19818 59814 19820 59866
rect 19574 59812 19580 59814
rect 19636 59812 19660 59814
rect 19716 59812 19740 59814
rect 19796 59812 19820 59814
rect 19876 59812 19882 59814
rect 19574 59792 19882 59812
rect 27528 59696 27580 59702
rect 27528 59638 27580 59644
rect 14648 59628 14700 59634
rect 14648 59570 14700 59576
rect 19984 59628 20036 59634
rect 19984 59570 20036 59576
rect 21180 59628 21232 59634
rect 21180 59570 21232 59576
rect 23848 59628 23900 59634
rect 23848 59570 23900 59576
rect 25964 59628 26016 59634
rect 25964 59570 26016 59576
rect 14096 59016 14148 59022
rect 14096 58958 14148 58964
rect 13084 58608 13136 58614
rect 13084 58550 13136 58556
rect 14108 58546 14136 58958
rect 14660 58682 14688 59570
rect 14740 59424 14792 59430
rect 14740 59366 14792 59372
rect 14752 59022 14780 59366
rect 19996 59022 20024 59570
rect 20168 59424 20220 59430
rect 20168 59366 20220 59372
rect 14740 59016 14792 59022
rect 14740 58958 14792 58964
rect 15936 59016 15988 59022
rect 15936 58958 15988 58964
rect 19984 59016 20036 59022
rect 19984 58958 20036 58964
rect 15844 58948 15896 58954
rect 15844 58890 15896 58896
rect 15476 58880 15528 58886
rect 15476 58822 15528 58828
rect 14648 58676 14700 58682
rect 14648 58618 14700 58624
rect 14096 58540 14148 58546
rect 14096 58482 14148 58488
rect 12900 58336 12952 58342
rect 12900 58278 12952 58284
rect 12808 57588 12860 57594
rect 12808 57530 12860 57536
rect 12256 57044 12308 57050
rect 12256 56986 12308 56992
rect 12912 56846 12940 58278
rect 13820 57860 13872 57866
rect 13820 57802 13872 57808
rect 13832 57458 13860 57802
rect 14096 57792 14148 57798
rect 14096 57734 14148 57740
rect 14108 57458 14136 57734
rect 15488 57526 15516 58822
rect 15476 57520 15528 57526
rect 15476 57462 15528 57468
rect 13820 57452 13872 57458
rect 13820 57394 13872 57400
rect 14096 57452 14148 57458
rect 14096 57394 14148 57400
rect 11520 56840 11572 56846
rect 11520 56782 11572 56788
rect 12900 56840 12952 56846
rect 12900 56782 12952 56788
rect 10324 56704 10376 56710
rect 10324 56646 10376 56652
rect 8944 56500 8996 56506
rect 8944 56442 8996 56448
rect 8956 55826 8984 56442
rect 10336 56438 10364 56646
rect 11532 56438 11560 56782
rect 10324 56432 10376 56438
rect 10324 56374 10376 56380
rect 11520 56432 11572 56438
rect 11520 56374 11572 56380
rect 10140 56160 10192 56166
rect 10140 56102 10192 56108
rect 8944 55820 8996 55826
rect 8944 55762 8996 55768
rect 10152 55758 10180 56102
rect 10140 55752 10192 55758
rect 10140 55694 10192 55700
rect 11704 55752 11756 55758
rect 11704 55694 11756 55700
rect 8760 55684 8812 55690
rect 8760 55626 8812 55632
rect 9312 55684 9364 55690
rect 9312 55626 9364 55632
rect 8392 55344 8444 55350
rect 8392 55286 8444 55292
rect 6920 55276 6972 55282
rect 6920 55218 6972 55224
rect 7932 55276 7984 55282
rect 7932 55218 7984 55224
rect 6932 55026 6960 55218
rect 7012 55072 7064 55078
rect 6932 55020 7012 55026
rect 6932 55014 7064 55020
rect 6932 54998 7052 55014
rect 6932 54738 6960 54998
rect 6920 54732 6972 54738
rect 6920 54674 6972 54680
rect 5632 54664 5684 54670
rect 5632 54606 5684 54612
rect 6276 54664 6328 54670
rect 6276 54606 6328 54612
rect 5644 53650 5672 54606
rect 5816 54596 5868 54602
rect 5816 54538 5868 54544
rect 5632 53644 5684 53650
rect 5632 53586 5684 53592
rect 5828 52698 5856 54538
rect 6288 54194 6316 54606
rect 7748 54596 7800 54602
rect 7748 54538 7800 54544
rect 6460 54528 6512 54534
rect 6460 54470 6512 54476
rect 7564 54528 7616 54534
rect 7564 54470 7616 54476
rect 6472 54262 6500 54470
rect 6460 54256 6512 54262
rect 6460 54198 6512 54204
rect 6276 54188 6328 54194
rect 6276 54130 6328 54136
rect 6288 53106 6316 54130
rect 7012 53440 7064 53446
rect 7012 53382 7064 53388
rect 6276 53100 6328 53106
rect 6276 53042 6328 53048
rect 5816 52692 5868 52698
rect 5816 52634 5868 52640
rect 7024 52494 7052 53382
rect 7576 53174 7604 54470
rect 7760 54330 7788 54538
rect 7748 54324 7800 54330
rect 7748 54266 7800 54272
rect 7944 53242 7972 55218
rect 9324 55214 9352 55626
rect 10324 55616 10376 55622
rect 10324 55558 10376 55564
rect 10336 55350 10364 55558
rect 10324 55344 10376 55350
rect 10324 55286 10376 55292
rect 9312 55208 9364 55214
rect 9312 55150 9364 55156
rect 9324 54194 9352 55150
rect 10692 55072 10744 55078
rect 10692 55014 10744 55020
rect 10704 54670 10732 55014
rect 9496 54664 9548 54670
rect 9496 54606 9548 54612
rect 10692 54664 10744 54670
rect 10692 54606 10744 54612
rect 9312 54188 9364 54194
rect 9312 54130 9364 54136
rect 9508 53582 9536 54606
rect 10876 54528 10928 54534
rect 10876 54470 10928 54476
rect 10888 54262 10916 54470
rect 10876 54256 10928 54262
rect 10876 54198 10928 54204
rect 11244 54188 11296 54194
rect 11244 54130 11296 54136
rect 10968 53984 11020 53990
rect 10968 53926 11020 53932
rect 10980 53582 11008 53926
rect 11256 53786 11284 54130
rect 11716 53990 11744 55694
rect 13728 55684 13780 55690
rect 13728 55626 13780 55632
rect 13740 55418 13768 55626
rect 13728 55412 13780 55418
rect 13728 55354 13780 55360
rect 11704 53984 11756 53990
rect 11704 53926 11756 53932
rect 12900 53984 12952 53990
rect 12900 53926 12952 53932
rect 11244 53780 11296 53786
rect 11244 53722 11296 53728
rect 11716 53582 11744 53926
rect 12912 53582 12940 53926
rect 9496 53576 9548 53582
rect 9496 53518 9548 53524
rect 10968 53576 11020 53582
rect 10968 53518 11020 53524
rect 11704 53576 11756 53582
rect 11704 53518 11756 53524
rect 12900 53576 12952 53582
rect 12900 53518 12952 53524
rect 7932 53236 7984 53242
rect 7932 53178 7984 53184
rect 7564 53168 7616 53174
rect 7564 53110 7616 53116
rect 9508 52698 9536 53518
rect 9496 52692 9548 52698
rect 9496 52634 9548 52640
rect 10140 52624 10192 52630
rect 10140 52566 10192 52572
rect 7012 52488 7064 52494
rect 7012 52430 7064 52436
rect 7012 52080 7064 52086
rect 7012 52022 7064 52028
rect 7024 51406 7052 52022
rect 8392 52012 8444 52018
rect 8392 51954 8444 51960
rect 7932 51808 7984 51814
rect 7932 51750 7984 51756
rect 7012 51400 7064 51406
rect 7012 51342 7064 51348
rect 6184 51332 6236 51338
rect 6184 51274 6236 51280
rect 5816 50720 5868 50726
rect 5816 50662 5868 50668
rect 5540 50312 5592 50318
rect 5540 50254 5592 50260
rect 5448 49700 5500 49706
rect 5448 49642 5500 49648
rect 4214 49532 4522 49552
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49456 4522 49476
rect 5460 49298 5488 49642
rect 4988 49292 5040 49298
rect 4988 49234 5040 49240
rect 5448 49292 5500 49298
rect 5448 49234 5500 49240
rect 5000 48754 5028 49234
rect 5552 48754 5580 50254
rect 5828 49910 5856 50662
rect 6196 50522 6224 51274
rect 6552 51264 6604 51270
rect 6552 51206 6604 51212
rect 6564 50998 6592 51206
rect 6552 50992 6604 50998
rect 6552 50934 6604 50940
rect 6184 50516 6236 50522
rect 6184 50458 6236 50464
rect 7024 50250 7052 51342
rect 7944 50318 7972 51750
rect 8404 51610 8432 51954
rect 8392 51604 8444 51610
rect 8392 51546 8444 51552
rect 9128 51332 9180 51338
rect 9128 51274 9180 51280
rect 9140 51066 9168 51274
rect 9128 51060 9180 51066
rect 9128 51002 9180 51008
rect 10152 50930 10180 52566
rect 10968 52488 11020 52494
rect 10968 52430 11020 52436
rect 11612 52488 11664 52494
rect 11716 52476 11744 53518
rect 13084 53440 13136 53446
rect 13084 53382 13136 53388
rect 13096 52494 13124 53382
rect 13832 53174 13860 57394
rect 14108 56914 14136 57394
rect 15476 57248 15528 57254
rect 15476 57190 15528 57196
rect 14096 56908 14148 56914
rect 14096 56850 14148 56856
rect 14108 56438 14136 56850
rect 15488 56846 15516 57190
rect 15856 57050 15884 58890
rect 15948 58002 15976 58958
rect 17316 58880 17368 58886
rect 17316 58822 17368 58828
rect 15936 57996 15988 58002
rect 15936 57938 15988 57944
rect 15844 57044 15896 57050
rect 15844 56986 15896 56992
rect 15476 56840 15528 56846
rect 15476 56782 15528 56788
rect 15948 56506 15976 57938
rect 15936 56500 15988 56506
rect 15936 56442 15988 56448
rect 17328 56438 17356 58822
rect 19574 58780 19882 58800
rect 19574 58778 19580 58780
rect 19636 58778 19660 58780
rect 19716 58778 19740 58780
rect 19796 58778 19820 58780
rect 19876 58778 19882 58780
rect 19636 58726 19638 58778
rect 19818 58726 19820 58778
rect 19574 58724 19580 58726
rect 19636 58724 19660 58726
rect 19716 58724 19740 58726
rect 19796 58724 19820 58726
rect 19876 58724 19882 58726
rect 19574 58704 19882 58724
rect 19996 58546 20024 58958
rect 19156 58540 19208 58546
rect 19156 58482 19208 58488
rect 19984 58540 20036 58546
rect 19984 58482 20036 58488
rect 18052 58472 18104 58478
rect 18052 58414 18104 58420
rect 18064 57934 18092 58414
rect 18052 57928 18104 57934
rect 18052 57870 18104 57876
rect 18064 57458 18092 57870
rect 18604 57860 18656 57866
rect 18604 57802 18656 57808
rect 18052 57452 18104 57458
rect 18052 57394 18104 57400
rect 18616 57050 18644 57802
rect 18696 57792 18748 57798
rect 18696 57734 18748 57740
rect 18604 57044 18656 57050
rect 18604 56986 18656 56992
rect 17868 56840 17920 56846
rect 17868 56782 17920 56788
rect 14096 56432 14148 56438
rect 14096 56374 14148 56380
rect 17316 56432 17368 56438
rect 17316 56374 17368 56380
rect 14108 55826 14136 56374
rect 15568 56364 15620 56370
rect 15568 56306 15620 56312
rect 14188 56160 14240 56166
rect 14188 56102 14240 56108
rect 14096 55820 14148 55826
rect 14096 55762 14148 55768
rect 14108 55214 14136 55762
rect 14200 55350 14228 56102
rect 14372 55616 14424 55622
rect 14372 55558 14424 55564
rect 14188 55344 14240 55350
rect 14188 55286 14240 55292
rect 14096 55208 14148 55214
rect 14096 55150 14148 55156
rect 14108 54738 14136 55150
rect 14096 54732 14148 54738
rect 14096 54674 14148 54680
rect 14384 54670 14412 55558
rect 15580 55418 15608 56306
rect 17880 56302 17908 56782
rect 17868 56296 17920 56302
rect 17868 56238 17920 56244
rect 16120 56160 16172 56166
rect 16120 56102 16172 56108
rect 16132 55758 16160 56102
rect 16120 55752 16172 55758
rect 16120 55694 16172 55700
rect 17880 55690 17908 56238
rect 18708 55758 18736 57734
rect 18696 55752 18748 55758
rect 18696 55694 18748 55700
rect 17868 55684 17920 55690
rect 17868 55626 17920 55632
rect 16028 55616 16080 55622
rect 16028 55558 16080 55564
rect 15568 55412 15620 55418
rect 15568 55354 15620 55360
rect 16040 55350 16068 55558
rect 16028 55344 16080 55350
rect 16028 55286 16080 55292
rect 17880 55282 17908 55626
rect 18696 55616 18748 55622
rect 18696 55558 18748 55564
rect 18708 55350 18736 55558
rect 19168 55418 19196 58482
rect 19340 58336 19392 58342
rect 19340 58278 19392 58284
rect 19248 56772 19300 56778
rect 19248 56714 19300 56720
rect 19260 56234 19288 56714
rect 19248 56228 19300 56234
rect 19248 56170 19300 56176
rect 19156 55412 19208 55418
rect 19156 55354 19208 55360
rect 19352 55350 19380 58278
rect 19996 58070 20024 58482
rect 19984 58064 20036 58070
rect 19984 58006 20036 58012
rect 19574 57692 19882 57712
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57616 19882 57636
rect 19996 57474 20024 58006
rect 19904 57458 20024 57474
rect 19892 57452 20024 57458
rect 19944 57446 20024 57452
rect 19892 57394 19944 57400
rect 19432 57248 19484 57254
rect 19432 57190 19484 57196
rect 19444 56438 19472 57190
rect 19904 56914 19932 57394
rect 19892 56908 19944 56914
rect 19944 56868 20024 56896
rect 19892 56850 19944 56856
rect 19574 56604 19882 56624
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56528 19882 56548
rect 19432 56432 19484 56438
rect 19432 56374 19484 56380
rect 19996 56370 20024 56868
rect 20180 56846 20208 59366
rect 21192 58682 21220 59570
rect 22468 59560 22520 59566
rect 22468 59502 22520 59508
rect 21272 58948 21324 58954
rect 21272 58890 21324 58896
rect 21180 58676 21232 58682
rect 21180 58618 21232 58624
rect 20444 57860 20496 57866
rect 20444 57802 20496 57808
rect 20168 56840 20220 56846
rect 20168 56782 20220 56788
rect 19984 56364 20036 56370
rect 19984 56306 20036 56312
rect 19996 55758 20024 56306
rect 19984 55752 20036 55758
rect 19984 55694 20036 55700
rect 19574 55516 19882 55536
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55440 19882 55460
rect 19996 55350 20024 55694
rect 18696 55344 18748 55350
rect 18696 55286 18748 55292
rect 19340 55344 19392 55350
rect 19340 55286 19392 55292
rect 19984 55344 20036 55350
rect 19984 55286 20036 55292
rect 17868 55276 17920 55282
rect 17868 55218 17920 55224
rect 14372 54664 14424 54670
rect 14372 54606 14424 54612
rect 16580 54664 16632 54670
rect 16580 54606 16632 54612
rect 16212 54596 16264 54602
rect 16212 54538 16264 54544
rect 15476 54528 15528 54534
rect 15476 54470 15528 54476
rect 15488 54262 15516 54470
rect 15476 54256 15528 54262
rect 15476 54198 15528 54204
rect 16028 53984 16080 53990
rect 16028 53926 16080 53932
rect 16040 53582 16068 53926
rect 16224 53786 16252 54538
rect 16592 54262 16620 54606
rect 16672 54528 16724 54534
rect 16672 54470 16724 54476
rect 16580 54256 16632 54262
rect 16580 54198 16632 54204
rect 16212 53780 16264 53786
rect 16212 53722 16264 53728
rect 16684 53582 16712 54470
rect 17880 54262 17908 55218
rect 19574 54428 19882 54448
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54352 19882 54372
rect 20456 54262 20484 57802
rect 21284 57594 21312 58890
rect 21916 58880 21968 58886
rect 21916 58822 21968 58828
rect 21928 58614 21956 58822
rect 21916 58608 21968 58614
rect 21916 58550 21968 58556
rect 22480 58546 22508 59502
rect 23480 59424 23532 59430
rect 23480 59366 23532 59372
rect 22468 58540 22520 58546
rect 22468 58482 22520 58488
rect 21272 57588 21324 57594
rect 21272 57530 21324 57536
rect 20628 57520 20680 57526
rect 20628 57462 20680 57468
rect 20640 55962 20668 57462
rect 22480 57390 22508 58482
rect 22468 57384 22520 57390
rect 22468 57326 22520 57332
rect 22480 56914 22508 57326
rect 22468 56908 22520 56914
rect 22468 56850 22520 56856
rect 20996 56704 21048 56710
rect 20996 56646 21048 56652
rect 21272 56704 21324 56710
rect 21272 56646 21324 56652
rect 20628 55956 20680 55962
rect 20628 55898 20680 55904
rect 21008 55418 21036 56646
rect 21284 56438 21312 56646
rect 21272 56432 21324 56438
rect 21272 56374 21324 56380
rect 22480 56370 22508 56850
rect 23492 56438 23520 59366
rect 23860 59226 23888 59570
rect 23940 59424 23992 59430
rect 23940 59366 23992 59372
rect 23848 59220 23900 59226
rect 23848 59162 23900 59168
rect 23848 58948 23900 58954
rect 23848 58890 23900 58896
rect 23756 57452 23808 57458
rect 23756 57394 23808 57400
rect 23768 56506 23796 57394
rect 23860 57050 23888 58890
rect 23952 58614 23980 59366
rect 25976 58682 26004 59570
rect 27252 59424 27304 59430
rect 27252 59366 27304 59372
rect 27264 59022 27292 59366
rect 27540 59226 27568 59638
rect 27528 59220 27580 59226
rect 27528 59162 27580 59168
rect 27540 59022 27568 59162
rect 27252 59016 27304 59022
rect 27252 58958 27304 58964
rect 27528 59016 27580 59022
rect 27528 58958 27580 58964
rect 27160 58880 27212 58886
rect 27160 58822 27212 58828
rect 25964 58676 26016 58682
rect 25964 58618 26016 58624
rect 23940 58608 23992 58614
rect 23940 58550 23992 58556
rect 26424 58540 26476 58546
rect 26424 58482 26476 58488
rect 24124 58336 24176 58342
rect 24124 58278 24176 58284
rect 24136 57526 24164 58278
rect 25044 57928 25096 57934
rect 25044 57870 25096 57876
rect 24124 57520 24176 57526
rect 24124 57462 24176 57468
rect 25056 57390 25084 57870
rect 26436 57594 26464 58482
rect 26424 57588 26476 57594
rect 26424 57530 26476 57536
rect 27172 57526 27200 58822
rect 27540 58478 27568 58958
rect 27528 58472 27580 58478
rect 27528 58414 27580 58420
rect 27540 57934 27568 58414
rect 27528 57928 27580 57934
rect 27528 57870 27580 57876
rect 27252 57792 27304 57798
rect 27252 57734 27304 57740
rect 27160 57520 27212 57526
rect 27160 57462 27212 57468
rect 25044 57384 25096 57390
rect 25044 57326 25096 57332
rect 24584 57248 24636 57254
rect 24584 57190 24636 57196
rect 23848 57044 23900 57050
rect 23848 56986 23900 56992
rect 24596 56846 24624 57190
rect 25056 57050 25084 57326
rect 25044 57044 25096 57050
rect 25044 56986 25096 56992
rect 24584 56840 24636 56846
rect 24584 56782 24636 56788
rect 26976 56840 27028 56846
rect 26976 56782 27028 56788
rect 23756 56500 23808 56506
rect 23756 56442 23808 56448
rect 23480 56432 23532 56438
rect 23480 56374 23532 56380
rect 22468 56364 22520 56370
rect 22468 56306 22520 56312
rect 25044 56364 25096 56370
rect 25044 56306 25096 56312
rect 21272 56160 21324 56166
rect 21272 56102 21324 56108
rect 21732 56160 21784 56166
rect 21732 56102 21784 56108
rect 21284 55758 21312 56102
rect 21744 55758 21772 56102
rect 22480 55758 22508 56306
rect 21272 55752 21324 55758
rect 21272 55694 21324 55700
rect 21732 55752 21784 55758
rect 21732 55694 21784 55700
rect 21824 55752 21876 55758
rect 21824 55694 21876 55700
rect 22468 55752 22520 55758
rect 22468 55694 22520 55700
rect 23664 55752 23716 55758
rect 23664 55694 23716 55700
rect 24400 55752 24452 55758
rect 24400 55694 24452 55700
rect 20996 55412 21048 55418
rect 20996 55354 21048 55360
rect 21744 54738 21772 55694
rect 21836 55214 21864 55694
rect 23204 55684 23256 55690
rect 23204 55626 23256 55632
rect 23216 55418 23244 55626
rect 23204 55412 23256 55418
rect 23204 55354 23256 55360
rect 23676 55282 23704 55694
rect 23848 55616 23900 55622
rect 23848 55558 23900 55564
rect 23112 55276 23164 55282
rect 23112 55218 23164 55224
rect 23664 55276 23716 55282
rect 23664 55218 23716 55224
rect 21824 55208 21876 55214
rect 21824 55150 21876 55156
rect 21732 54732 21784 54738
rect 21732 54674 21784 54680
rect 20720 54664 20772 54670
rect 20772 54612 20852 54618
rect 20720 54606 20852 54612
rect 20732 54590 20852 54606
rect 17868 54256 17920 54262
rect 17868 54198 17920 54204
rect 20076 54256 20128 54262
rect 20076 54198 20128 54204
rect 20444 54256 20496 54262
rect 20444 54198 20496 54204
rect 17776 54188 17828 54194
rect 17776 54130 17828 54136
rect 17788 53786 17816 54130
rect 17776 53780 17828 53786
rect 17776 53722 17828 53728
rect 17880 53582 17908 54198
rect 18052 53984 18104 53990
rect 18052 53926 18104 53932
rect 16028 53576 16080 53582
rect 16028 53518 16080 53524
rect 16672 53576 16724 53582
rect 16672 53518 16724 53524
rect 17868 53576 17920 53582
rect 17868 53518 17920 53524
rect 14648 53508 14700 53514
rect 14648 53450 14700 53456
rect 14660 53174 14688 53450
rect 18064 53174 18092 53926
rect 18512 53576 18564 53582
rect 18512 53518 18564 53524
rect 13360 53168 13412 53174
rect 13360 53110 13412 53116
rect 13820 53168 13872 53174
rect 13820 53110 13872 53116
rect 14648 53168 14700 53174
rect 14648 53110 14700 53116
rect 18052 53168 18104 53174
rect 18052 53110 18104 53116
rect 11664 52448 11744 52476
rect 11612 52430 11664 52436
rect 10980 52154 11008 52430
rect 10968 52148 11020 52154
rect 10968 52090 11020 52096
rect 11716 52034 11744 52448
rect 13084 52488 13136 52494
rect 13084 52430 13136 52436
rect 12900 52352 12952 52358
rect 12900 52294 12952 52300
rect 12912 52086 12940 52294
rect 13372 52154 13400 53110
rect 14660 52494 14688 53110
rect 18524 53106 18552 53518
rect 19984 53508 20036 53514
rect 19984 53450 20036 53456
rect 19574 53340 19882 53360
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53264 19882 53284
rect 19996 53242 20024 53450
rect 19984 53236 20036 53242
rect 19984 53178 20036 53184
rect 18512 53100 18564 53106
rect 18512 53042 18564 53048
rect 18604 53100 18656 53106
rect 18604 53042 18656 53048
rect 17408 52896 17460 52902
rect 17408 52838 17460 52844
rect 17420 52494 17448 52838
rect 18616 52698 18644 53042
rect 18604 52692 18656 52698
rect 18604 52634 18656 52640
rect 14096 52488 14148 52494
rect 14096 52430 14148 52436
rect 14648 52488 14700 52494
rect 14648 52430 14700 52436
rect 16672 52488 16724 52494
rect 16672 52430 16724 52436
rect 17408 52488 17460 52494
rect 17408 52430 17460 52436
rect 13820 52420 13872 52426
rect 13820 52362 13872 52368
rect 13360 52148 13412 52154
rect 13360 52090 13412 52096
rect 11624 52018 11744 52034
rect 12900 52080 12952 52086
rect 12900 52022 12952 52028
rect 10968 52012 11020 52018
rect 10968 51954 11020 51960
rect 11612 52012 11744 52018
rect 11664 52006 11744 52012
rect 11612 51954 11664 51960
rect 10980 51066 11008 51954
rect 11716 51406 11744 52006
rect 13636 52012 13688 52018
rect 13636 51954 13688 51960
rect 13648 51610 13676 51954
rect 13832 51882 13860 52362
rect 14108 51950 14136 52430
rect 15200 52352 15252 52358
rect 15200 52294 15252 52300
rect 14004 51944 14056 51950
rect 14004 51886 14056 51892
rect 14096 51944 14148 51950
rect 14096 51886 14148 51892
rect 13820 51876 13872 51882
rect 13820 51818 13872 51824
rect 14016 51610 14044 51886
rect 13636 51604 13688 51610
rect 13636 51546 13688 51552
rect 14004 51604 14056 51610
rect 14004 51546 14056 51552
rect 14108 51474 14136 51886
rect 14096 51468 14148 51474
rect 14096 51410 14148 51416
rect 11704 51400 11756 51406
rect 11704 51342 11756 51348
rect 11612 51264 11664 51270
rect 11612 51206 11664 51212
rect 10968 51060 11020 51066
rect 10968 51002 11020 51008
rect 11624 50998 11652 51206
rect 11612 50992 11664 50998
rect 11612 50934 11664 50940
rect 10140 50924 10192 50930
rect 10140 50866 10192 50872
rect 11244 50924 11296 50930
rect 11244 50866 11296 50872
rect 8116 50720 8168 50726
rect 8116 50662 8168 50668
rect 7932 50312 7984 50318
rect 7932 50254 7984 50260
rect 8128 50250 8156 50662
rect 11256 50522 11284 50866
rect 11716 50862 11744 51342
rect 12164 51332 12216 51338
rect 12164 51274 12216 51280
rect 12176 51066 12204 51274
rect 12164 51060 12216 51066
rect 12164 51002 12216 51008
rect 14108 50862 14136 51410
rect 15212 51338 15240 52294
rect 16684 52018 16712 52430
rect 19574 52252 19882 52272
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52176 19882 52196
rect 16672 52012 16724 52018
rect 16672 51954 16724 51960
rect 18052 52012 18104 52018
rect 18052 51954 18104 51960
rect 15476 51808 15528 51814
rect 15476 51750 15528 51756
rect 15488 51406 15516 51750
rect 16684 51406 16712 51954
rect 17776 51808 17828 51814
rect 17776 51750 17828 51756
rect 15476 51400 15528 51406
rect 15476 51342 15528 51348
rect 16672 51400 16724 51406
rect 16672 51342 16724 51348
rect 15200 51332 15252 51338
rect 15200 51274 15252 51280
rect 15568 51332 15620 51338
rect 15568 51274 15620 51280
rect 15476 51264 15528 51270
rect 15476 51206 15528 51212
rect 15488 50998 15516 51206
rect 15476 50992 15528 50998
rect 15476 50934 15528 50940
rect 11704 50856 11756 50862
rect 11704 50798 11756 50804
rect 14096 50856 14148 50862
rect 14096 50798 14148 50804
rect 14108 50522 14136 50798
rect 15476 50720 15528 50726
rect 15476 50662 15528 50668
rect 11244 50516 11296 50522
rect 11244 50458 11296 50464
rect 14096 50516 14148 50522
rect 14096 50458 14148 50464
rect 15488 50318 15516 50662
rect 15580 50522 15608 51274
rect 16684 50862 16712 51342
rect 17316 51264 17368 51270
rect 17316 51206 17368 51212
rect 16672 50856 16724 50862
rect 16672 50798 16724 50804
rect 17040 50720 17092 50726
rect 17040 50662 17092 50668
rect 15568 50516 15620 50522
rect 15568 50458 15620 50464
rect 8944 50312 8996 50318
rect 8944 50254 8996 50260
rect 13820 50312 13872 50318
rect 13820 50254 13872 50260
rect 15476 50312 15528 50318
rect 15476 50254 15528 50260
rect 7012 50244 7064 50250
rect 7012 50186 7064 50192
rect 8116 50244 8168 50250
rect 8116 50186 8168 50192
rect 6368 50176 6420 50182
rect 6368 50118 6420 50124
rect 5816 49904 5868 49910
rect 5816 49846 5868 49852
rect 6380 49774 6408 50118
rect 6460 49836 6512 49842
rect 6460 49778 6512 49784
rect 6368 49768 6420 49774
rect 6368 49710 6420 49716
rect 5816 49632 5868 49638
rect 5816 49574 5868 49580
rect 5828 48822 5856 49574
rect 6472 49434 6500 49778
rect 7748 49632 7800 49638
rect 7748 49574 7800 49580
rect 6460 49428 6512 49434
rect 6460 49370 6512 49376
rect 7760 49230 7788 49574
rect 7748 49224 7800 49230
rect 7748 49166 7800 49172
rect 5816 48816 5868 48822
rect 5816 48758 5868 48764
rect 8128 48754 8156 50186
rect 8956 49774 8984 50254
rect 10784 50244 10836 50250
rect 10784 50186 10836 50192
rect 10232 49836 10284 49842
rect 10232 49778 10284 49784
rect 8944 49768 8996 49774
rect 8944 49710 8996 49716
rect 8956 49230 8984 49710
rect 8944 49224 8996 49230
rect 8944 49166 8996 49172
rect 4988 48748 5040 48754
rect 4988 48690 5040 48696
rect 5540 48748 5592 48754
rect 5540 48690 5592 48696
rect 8116 48748 8168 48754
rect 8116 48690 8168 48696
rect 4214 48444 4522 48464
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48368 4522 48388
rect 5000 48210 5028 48690
rect 4988 48204 5040 48210
rect 4988 48146 5040 48152
rect 5000 47734 5028 48146
rect 8956 48142 8984 49166
rect 10244 48890 10272 49778
rect 10416 49632 10468 49638
rect 10416 49574 10468 49580
rect 10324 49088 10376 49094
rect 10324 49030 10376 49036
rect 10232 48884 10284 48890
rect 10232 48826 10284 48832
rect 10336 48822 10364 49030
rect 10324 48816 10376 48822
rect 10324 48758 10376 48764
rect 10428 48142 10456 49574
rect 10796 48278 10824 50186
rect 13544 50176 13596 50182
rect 13544 50118 13596 50124
rect 13556 49230 13584 50118
rect 13728 49836 13780 49842
rect 13832 49824 13860 50254
rect 16120 50244 16172 50250
rect 16120 50186 16172 50192
rect 16132 49978 16160 50186
rect 16120 49972 16172 49978
rect 16120 49914 16172 49920
rect 16028 49904 16080 49910
rect 16028 49846 16080 49852
rect 13780 49796 13860 49824
rect 13728 49778 13780 49784
rect 13832 49366 13860 49796
rect 13912 49836 13964 49842
rect 13912 49778 13964 49784
rect 13924 49434 13952 49778
rect 14740 49768 14792 49774
rect 14740 49710 14792 49716
rect 14372 49632 14424 49638
rect 14372 49574 14424 49580
rect 13912 49428 13964 49434
rect 13912 49370 13964 49376
rect 13820 49360 13872 49366
rect 13820 49302 13872 49308
rect 14384 49230 14412 49574
rect 14752 49450 14780 49710
rect 14752 49434 14872 49450
rect 14740 49428 14872 49434
rect 14792 49422 14872 49428
rect 14740 49370 14792 49376
rect 14752 49339 14780 49370
rect 12164 49224 12216 49230
rect 12164 49166 12216 49172
rect 13544 49224 13596 49230
rect 13544 49166 13596 49172
rect 14372 49224 14424 49230
rect 14372 49166 14424 49172
rect 12176 48822 12204 49166
rect 12164 48816 12216 48822
rect 12164 48758 12216 48764
rect 12900 48748 12952 48754
rect 12900 48690 12952 48696
rect 13636 48748 13688 48754
rect 13636 48690 13688 48696
rect 11888 48544 11940 48550
rect 11888 48486 11940 48492
rect 10784 48272 10836 48278
rect 10784 48214 10836 48220
rect 8944 48136 8996 48142
rect 8944 48078 8996 48084
rect 10416 48136 10468 48142
rect 10416 48078 10468 48084
rect 11520 48136 11572 48142
rect 11520 48078 11572 48084
rect 5908 48068 5960 48074
rect 5908 48010 5960 48016
rect 4988 47728 5040 47734
rect 4988 47670 5040 47676
rect 5000 47598 5028 47670
rect 5172 47660 5224 47666
rect 5172 47602 5224 47608
rect 4988 47592 5040 47598
rect 4988 47534 5040 47540
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 5184 47258 5212 47602
rect 5448 47592 5500 47598
rect 5448 47534 5500 47540
rect 5172 47252 5224 47258
rect 5172 47194 5224 47200
rect 5460 47122 5488 47534
rect 5724 47456 5776 47462
rect 5724 47398 5776 47404
rect 5448 47116 5500 47122
rect 5448 47058 5500 47064
rect 4344 47048 4396 47054
rect 4344 46990 4396 46996
rect 4356 46578 4384 46990
rect 4620 46640 4672 46646
rect 4620 46582 4672 46588
rect 4344 46572 4396 46578
rect 4344 46514 4396 46520
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4632 46050 4660 46582
rect 5460 46510 5488 47058
rect 5736 47054 5764 47398
rect 5816 47252 5868 47258
rect 5816 47194 5868 47200
rect 5724 47048 5776 47054
rect 5724 46990 5776 46996
rect 5540 46980 5592 46986
rect 5540 46922 5592 46928
rect 5552 46714 5580 46922
rect 5540 46708 5592 46714
rect 5540 46650 5592 46656
rect 5448 46504 5500 46510
rect 5448 46446 5500 46452
rect 5460 46170 5488 46446
rect 5448 46164 5500 46170
rect 5448 46106 5500 46112
rect 4540 46034 4660 46050
rect 4528 46028 4660 46034
rect 4580 46022 4660 46028
rect 4528 45970 4580 45976
rect 5828 45966 5856 47194
rect 5920 46170 5948 48010
rect 6368 48000 6420 48006
rect 6368 47942 6420 47948
rect 6380 46646 6408 47942
rect 7748 47660 7800 47666
rect 7748 47602 7800 47608
rect 7288 47456 7340 47462
rect 7288 47398 7340 47404
rect 6368 46640 6420 46646
rect 6368 46582 6420 46588
rect 5908 46164 5960 46170
rect 5908 46106 5960 46112
rect 7300 45966 7328 47398
rect 7760 46714 7788 47602
rect 11428 47048 11480 47054
rect 11532 47036 11560 48078
rect 11900 47734 11928 48486
rect 12912 48278 12940 48690
rect 12900 48272 12952 48278
rect 12900 48214 12952 48220
rect 12900 48068 12952 48074
rect 12900 48010 12952 48016
rect 11888 47728 11940 47734
rect 11888 47670 11940 47676
rect 11480 47008 11560 47036
rect 11428 46990 11480 46996
rect 7748 46708 7800 46714
rect 7748 46650 7800 46656
rect 7840 46572 7892 46578
rect 7840 46514 7892 46520
rect 7852 46170 7880 46514
rect 11532 46510 11560 47008
rect 12164 46980 12216 46986
rect 12164 46922 12216 46928
rect 11980 46912 12032 46918
rect 11980 46854 12032 46860
rect 11992 46646 12020 46854
rect 11980 46640 12032 46646
rect 11980 46582 12032 46588
rect 11520 46504 11572 46510
rect 11520 46446 11572 46452
rect 8944 46368 8996 46374
rect 8944 46310 8996 46316
rect 9588 46368 9640 46374
rect 9588 46310 9640 46316
rect 7840 46164 7892 46170
rect 7840 46106 7892 46112
rect 8956 45966 8984 46310
rect 5816 45960 5868 45966
rect 5816 45902 5868 45908
rect 7288 45960 7340 45966
rect 7288 45902 7340 45908
rect 8944 45960 8996 45966
rect 8944 45902 8996 45908
rect 4620 45892 4672 45898
rect 4620 45834 4672 45840
rect 8576 45892 8628 45898
rect 8576 45834 8628 45840
rect 4632 45626 4660 45834
rect 8588 45626 8616 45834
rect 4620 45620 4672 45626
rect 4620 45562 4672 45568
rect 8576 45620 8628 45626
rect 8576 45562 8628 45568
rect 9600 45490 9628 46310
rect 11532 45966 11560 46446
rect 12176 46170 12204 46922
rect 12912 46714 12940 48010
rect 13648 47598 13676 48690
rect 14188 48544 14240 48550
rect 14188 48486 14240 48492
rect 14200 47666 14228 48486
rect 14844 48346 14872 49422
rect 15476 48748 15528 48754
rect 15476 48690 15528 48696
rect 14924 48544 14976 48550
rect 14924 48486 14976 48492
rect 14832 48340 14884 48346
rect 14832 48282 14884 48288
rect 14936 48142 14964 48486
rect 14924 48136 14976 48142
rect 14924 48078 14976 48084
rect 14832 48068 14884 48074
rect 14832 48010 14884 48016
rect 14188 47660 14240 47666
rect 14188 47602 14240 47608
rect 13636 47592 13688 47598
rect 13636 47534 13688 47540
rect 12900 46708 12952 46714
rect 12900 46650 12952 46656
rect 13648 46578 13676 47534
rect 14844 47462 14872 48010
rect 15488 47802 15516 48690
rect 16040 48278 16068 49846
rect 17052 49298 17080 50662
rect 17328 50318 17356 51206
rect 17408 50924 17460 50930
rect 17408 50866 17460 50872
rect 17420 50522 17448 50866
rect 17408 50516 17460 50522
rect 17408 50458 17460 50464
rect 17316 50312 17368 50318
rect 17316 50254 17368 50260
rect 17040 49292 17092 49298
rect 17040 49234 17092 49240
rect 17052 48754 17080 49234
rect 17788 49230 17816 51750
rect 18064 51066 18092 51954
rect 19248 51944 19300 51950
rect 19248 51886 19300 51892
rect 18052 51060 18104 51066
rect 18052 51002 18104 51008
rect 19260 50726 19288 51886
rect 20088 51542 20116 54198
rect 20824 54126 20852 54590
rect 21088 54596 21140 54602
rect 21088 54538 21140 54544
rect 20812 54120 20864 54126
rect 20812 54062 20864 54068
rect 20824 53582 20852 54062
rect 21100 53786 21128 54538
rect 21272 54528 21324 54534
rect 21272 54470 21324 54476
rect 21284 54262 21312 54470
rect 21272 54256 21324 54262
rect 21272 54198 21324 54204
rect 21836 54126 21864 55150
rect 23124 54874 23152 55218
rect 23860 55214 23888 55558
rect 24412 55350 24440 55694
rect 25056 55418 25084 56306
rect 25596 56160 25648 56166
rect 25596 56102 25648 56108
rect 25412 55684 25464 55690
rect 25412 55626 25464 55632
rect 25044 55412 25096 55418
rect 25044 55354 25096 55360
rect 24400 55344 24452 55350
rect 24400 55286 24452 55292
rect 23860 55186 23980 55214
rect 23112 54868 23164 54874
rect 23112 54810 23164 54816
rect 23664 54664 23716 54670
rect 23664 54606 23716 54612
rect 23204 54596 23256 54602
rect 23204 54538 23256 54544
rect 23216 54330 23244 54538
rect 23204 54324 23256 54330
rect 23204 54266 23256 54272
rect 23676 54194 23704 54606
rect 23952 54262 23980 55186
rect 24412 54670 24440 55286
rect 25044 55276 25096 55282
rect 25044 55218 25096 55224
rect 24400 54664 24452 54670
rect 24400 54606 24452 54612
rect 25056 54330 25084 55218
rect 25424 54874 25452 55626
rect 25412 54868 25464 54874
rect 25412 54810 25464 54816
rect 25608 54670 25636 56102
rect 26988 55758 27016 56782
rect 27264 55758 27292 57734
rect 27540 57390 27568 57870
rect 27528 57384 27580 57390
rect 27528 57326 27580 57332
rect 27540 56846 27568 57326
rect 27528 56840 27580 56846
rect 27528 56782 27580 56788
rect 27620 56772 27672 56778
rect 27620 56714 27672 56720
rect 27632 56438 27660 56714
rect 27620 56432 27672 56438
rect 27620 56374 27672 56380
rect 26976 55752 27028 55758
rect 26976 55694 27028 55700
rect 27252 55752 27304 55758
rect 27252 55694 27304 55700
rect 26988 55078 27016 55694
rect 26976 55072 27028 55078
rect 26976 55014 27028 55020
rect 26988 54670 27016 55014
rect 25596 54664 25648 54670
rect 25596 54606 25648 54612
rect 26976 54664 27028 54670
rect 26976 54606 27028 54612
rect 25044 54324 25096 54330
rect 25044 54266 25096 54272
rect 23940 54256 23992 54262
rect 23940 54198 23992 54204
rect 26988 54194 27016 54606
rect 23664 54188 23716 54194
rect 23664 54130 23716 54136
rect 26976 54188 27028 54194
rect 26976 54130 27028 54136
rect 27252 54188 27304 54194
rect 27252 54130 27304 54136
rect 21824 54120 21876 54126
rect 21824 54062 21876 54068
rect 21088 53780 21140 53786
rect 21088 53722 21140 53728
rect 21836 53582 21864 54062
rect 26988 53582 27016 54130
rect 27264 53786 27292 54130
rect 27252 53780 27304 53786
rect 27252 53722 27304 53728
rect 20812 53576 20864 53582
rect 20812 53518 20864 53524
rect 21824 53576 21876 53582
rect 21824 53518 21876 53524
rect 25044 53576 25096 53582
rect 25044 53518 25096 53524
rect 26976 53576 27028 53582
rect 26976 53518 27028 53524
rect 20720 53508 20772 53514
rect 20720 53450 20772 53456
rect 20628 53440 20680 53446
rect 20628 53382 20680 53388
rect 20640 52494 20668 53382
rect 20628 52488 20680 52494
rect 20628 52430 20680 52436
rect 20732 52154 20760 53450
rect 20824 52426 20852 53518
rect 25056 53106 25084 53518
rect 26424 53508 26476 53514
rect 26424 53450 26476 53456
rect 26436 53242 26464 53450
rect 26424 53236 26476 53242
rect 26424 53178 26476 53184
rect 24860 53100 24912 53106
rect 24860 53042 24912 53048
rect 25044 53100 25096 53106
rect 25044 53042 25096 53048
rect 26240 53100 26292 53106
rect 26240 53042 26292 53048
rect 23020 52624 23072 52630
rect 23020 52566 23072 52572
rect 21732 52488 21784 52494
rect 21732 52430 21784 52436
rect 20812 52420 20864 52426
rect 20812 52362 20864 52368
rect 20720 52148 20772 52154
rect 20720 52090 20772 52096
rect 19340 51536 19392 51542
rect 19340 51478 19392 51484
rect 20076 51536 20128 51542
rect 20076 51478 20128 51484
rect 20720 51536 20772 51542
rect 20720 51478 20772 51484
rect 19248 50720 19300 50726
rect 19248 50662 19300 50668
rect 19260 50386 19288 50662
rect 19248 50380 19300 50386
rect 19248 50322 19300 50328
rect 19260 49910 19288 50322
rect 19248 49904 19300 49910
rect 19248 49846 19300 49852
rect 19352 49842 19380 51478
rect 20088 51270 20116 51478
rect 20076 51264 20128 51270
rect 20076 51206 20128 51212
rect 19574 51164 19882 51184
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51088 19882 51108
rect 20076 50720 20128 50726
rect 20076 50662 20128 50668
rect 19574 50076 19882 50096
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50000 19882 50020
rect 20088 49910 20116 50662
rect 20076 49904 20128 49910
rect 20076 49846 20128 49852
rect 19340 49836 19392 49842
rect 19340 49778 19392 49784
rect 19708 49836 19760 49842
rect 19708 49778 19760 49784
rect 19720 49298 19748 49778
rect 19432 49292 19484 49298
rect 19432 49234 19484 49240
rect 19708 49292 19760 49298
rect 19708 49234 19760 49240
rect 17776 49224 17828 49230
rect 17776 49166 17828 49172
rect 18604 49088 18656 49094
rect 18604 49030 18656 49036
rect 18616 48822 18644 49030
rect 18604 48816 18656 48822
rect 18604 48758 18656 48764
rect 19444 48754 19472 49234
rect 19574 48988 19882 49008
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48912 19882 48932
rect 17040 48748 17092 48754
rect 17040 48690 17092 48696
rect 19432 48748 19484 48754
rect 19432 48690 19484 48696
rect 17052 48346 17080 48690
rect 18328 48544 18380 48550
rect 18328 48486 18380 48492
rect 17040 48340 17092 48346
rect 17040 48282 17092 48288
rect 16028 48272 16080 48278
rect 16028 48214 16080 48220
rect 15476 47796 15528 47802
rect 15476 47738 15528 47744
rect 17052 47666 17080 48282
rect 18340 48142 18368 48486
rect 19444 48210 19472 48690
rect 19432 48204 19484 48210
rect 19432 48146 19484 48152
rect 18328 48136 18380 48142
rect 18328 48078 18380 48084
rect 18420 48000 18472 48006
rect 18420 47942 18472 47948
rect 18432 47734 18460 47942
rect 18420 47728 18472 47734
rect 18420 47670 18472 47676
rect 19444 47666 19472 48146
rect 19574 47900 19882 47920
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47824 19882 47844
rect 17040 47660 17092 47666
rect 17040 47602 17092 47608
rect 19432 47660 19484 47666
rect 19432 47602 19484 47608
rect 14832 47456 14884 47462
rect 14832 47398 14884 47404
rect 14844 47054 14872 47398
rect 17052 47138 17080 47602
rect 18328 47456 18380 47462
rect 18328 47398 18380 47404
rect 16960 47110 17080 47138
rect 16960 47054 16988 47110
rect 18340 47054 18368 47398
rect 19444 47122 19472 47602
rect 19432 47116 19484 47122
rect 19432 47058 19484 47064
rect 14832 47048 14884 47054
rect 14832 46990 14884 46996
rect 16948 47048 17000 47054
rect 16948 46990 17000 46996
rect 18328 47048 18380 47054
rect 18328 46990 18380 46996
rect 13636 46572 13688 46578
rect 13636 46514 13688 46520
rect 12164 46164 12216 46170
rect 12164 46106 12216 46112
rect 11520 45960 11572 45966
rect 11520 45902 11572 45908
rect 10324 45824 10376 45830
rect 10324 45766 10376 45772
rect 10336 45558 10364 45766
rect 10324 45552 10376 45558
rect 10324 45494 10376 45500
rect 11532 45490 11560 45902
rect 12900 45892 12952 45898
rect 12900 45834 12952 45840
rect 12912 45626 12940 45834
rect 12900 45620 12952 45626
rect 12900 45562 12952 45568
rect 13648 45558 13676 46514
rect 14844 45898 14872 46990
rect 16212 46912 16264 46918
rect 16212 46854 16264 46860
rect 16224 46646 16252 46854
rect 16212 46640 16264 46646
rect 16212 46582 16264 46588
rect 16120 46368 16172 46374
rect 16120 46310 16172 46316
rect 16132 45966 16160 46310
rect 16960 46170 16988 46990
rect 17960 46980 18012 46986
rect 17960 46922 18012 46928
rect 16948 46164 17000 46170
rect 16948 46106 17000 46112
rect 16120 45960 16172 45966
rect 16120 45902 16172 45908
rect 14832 45892 14884 45898
rect 14832 45834 14884 45840
rect 15752 45824 15804 45830
rect 15752 45766 15804 45772
rect 15764 45558 15792 45766
rect 13636 45552 13688 45558
rect 13636 45494 13688 45500
rect 15752 45552 15804 45558
rect 15752 45494 15804 45500
rect 9588 45484 9640 45490
rect 9588 45426 9640 45432
rect 11520 45484 11572 45490
rect 11520 45426 11572 45432
rect 12900 45484 12952 45490
rect 12900 45426 12952 45432
rect 7196 45416 7248 45422
rect 7196 45358 7248 45364
rect 9036 45416 9088 45422
rect 9036 45358 9088 45364
rect 7208 45286 7236 45358
rect 6368 45280 6420 45286
rect 6368 45222 6420 45228
rect 7196 45280 7248 45286
rect 7196 45222 7248 45228
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 6380 44878 6408 45222
rect 6368 44872 6420 44878
rect 6368 44814 6420 44820
rect 5356 44396 5408 44402
rect 5356 44338 5408 44344
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 5368 43450 5396 44338
rect 6380 44334 6408 44814
rect 7208 44470 7236 45222
rect 9048 44878 9076 45358
rect 10416 45280 10468 45286
rect 10416 45222 10468 45228
rect 9036 44872 9088 44878
rect 9036 44814 9088 44820
rect 9496 44872 9548 44878
rect 9496 44814 9548 44820
rect 7656 44804 7708 44810
rect 7656 44746 7708 44752
rect 7668 44538 7696 44746
rect 7748 44736 7800 44742
rect 7748 44678 7800 44684
rect 7656 44532 7708 44538
rect 7656 44474 7708 44480
rect 7196 44464 7248 44470
rect 7196 44406 7248 44412
rect 7472 44396 7524 44402
rect 7472 44338 7524 44344
rect 6368 44328 6420 44334
rect 6368 44270 6420 44276
rect 5724 44192 5776 44198
rect 5724 44134 5776 44140
rect 5632 43716 5684 43722
rect 5632 43658 5684 43664
rect 5356 43444 5408 43450
rect 5356 43386 5408 43392
rect 5172 43308 5224 43314
rect 5172 43250 5224 43256
rect 3792 43240 3844 43246
rect 3792 43182 3844 43188
rect 3804 42022 3832 43182
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 5184 42906 5212 43250
rect 5172 42900 5224 42906
rect 5172 42842 5224 42848
rect 5172 42628 5224 42634
rect 5172 42570 5224 42576
rect 3792 42016 3844 42022
rect 3792 41958 3844 41964
rect 4068 42016 4120 42022
rect 4068 41958 4120 41964
rect 3804 41614 3832 41958
rect 4080 41614 4108 41958
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 5184 41818 5212 42570
rect 5448 42220 5500 42226
rect 5448 42162 5500 42168
rect 5172 41812 5224 41818
rect 5172 41754 5224 41760
rect 3792 41608 3844 41614
rect 3792 41550 3844 41556
rect 4068 41608 4120 41614
rect 4068 41550 4120 41556
rect 3804 41070 3832 41550
rect 5460 41274 5488 42162
rect 5448 41268 5500 41274
rect 5448 41210 5500 41216
rect 3792 41064 3844 41070
rect 3792 41006 3844 41012
rect 3804 40118 3832 41006
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 5644 40118 5672 43658
rect 5736 43382 5764 44134
rect 6380 43994 6408 44270
rect 6368 43988 6420 43994
rect 6368 43930 6420 43936
rect 6828 43988 6880 43994
rect 6828 43930 6880 43936
rect 6840 43382 6868 43930
rect 7484 43450 7512 44338
rect 7760 43790 7788 44678
rect 9508 44334 9536 44814
rect 9588 44804 9640 44810
rect 9588 44746 9640 44752
rect 9600 44538 9628 44746
rect 9588 44532 9640 44538
rect 9588 44474 9640 44480
rect 10428 44470 10456 45222
rect 10784 44872 10836 44878
rect 10784 44814 10836 44820
rect 10416 44464 10468 44470
rect 10416 44406 10468 44412
rect 10796 44402 10824 44814
rect 12164 44736 12216 44742
rect 12164 44678 12216 44684
rect 12176 44470 12204 44678
rect 12912 44538 12940 45426
rect 12900 44532 12952 44538
rect 12900 44474 12952 44480
rect 12164 44464 12216 44470
rect 12164 44406 12216 44412
rect 13648 44402 13676 45494
rect 16672 45416 16724 45422
rect 16672 45358 16724 45364
rect 15476 45280 15528 45286
rect 15476 45222 15528 45228
rect 15488 44878 15516 45222
rect 16684 44946 16712 45358
rect 17972 45354 18000 46922
rect 18236 46912 18288 46918
rect 18236 46854 18288 46860
rect 18248 46646 18276 46854
rect 18236 46640 18288 46646
rect 18236 46582 18288 46588
rect 19444 46578 19472 47058
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19432 46572 19484 46578
rect 19432 46514 19484 46520
rect 18144 46368 18196 46374
rect 18144 46310 18196 46316
rect 18156 45966 18184 46310
rect 19444 46034 19472 46514
rect 19432 46028 19484 46034
rect 19432 45970 19484 45976
rect 18144 45960 18196 45966
rect 18144 45902 18196 45908
rect 18052 45824 18104 45830
rect 18052 45766 18104 45772
rect 18064 45558 18092 45766
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 18052 45552 18104 45558
rect 20732 45554 20760 51478
rect 20824 51406 20852 52362
rect 21364 52352 21416 52358
rect 21364 52294 21416 52300
rect 21376 52086 21404 52294
rect 21364 52080 21416 52086
rect 21364 52022 21416 52028
rect 20812 51400 20864 51406
rect 20812 51342 20864 51348
rect 21272 51332 21324 51338
rect 21272 51274 21324 51280
rect 21180 51264 21232 51270
rect 21180 51206 21232 51212
rect 21088 50244 21140 50250
rect 21088 50186 21140 50192
rect 21100 49978 21128 50186
rect 21088 49972 21140 49978
rect 21088 49914 21140 49920
rect 21088 49836 21140 49842
rect 21088 49778 21140 49784
rect 21100 49434 21128 49778
rect 21088 49428 21140 49434
rect 21088 49370 21140 49376
rect 20996 49156 21048 49162
rect 20996 49098 21048 49104
rect 21008 48890 21036 49098
rect 20996 48884 21048 48890
rect 20996 48826 21048 48832
rect 20812 48748 20864 48754
rect 20812 48690 20864 48696
rect 20824 48278 20852 48690
rect 20812 48272 20864 48278
rect 20812 48214 20864 48220
rect 21192 48142 21220 51206
rect 21284 51066 21312 51274
rect 21272 51060 21324 51066
rect 21272 51002 21324 51008
rect 21744 50386 21772 52430
rect 21824 51944 21876 51950
rect 21824 51886 21876 51892
rect 21836 51406 21864 51886
rect 21824 51400 21876 51406
rect 21824 51342 21876 51348
rect 22100 51264 22152 51270
rect 22100 51206 22152 51212
rect 22112 50998 22140 51206
rect 22100 50992 22152 50998
rect 22100 50934 22152 50940
rect 22468 50720 22520 50726
rect 22468 50662 22520 50668
rect 21732 50380 21784 50386
rect 21732 50322 21784 50328
rect 21744 49774 21772 50322
rect 21732 49768 21784 49774
rect 21732 49710 21784 49716
rect 21744 49298 21772 49710
rect 21732 49292 21784 49298
rect 21732 49234 21784 49240
rect 22480 48754 22508 50662
rect 22468 48748 22520 48754
rect 22468 48690 22520 48696
rect 22480 48346 22508 48690
rect 22468 48340 22520 48346
rect 22468 48282 22520 48288
rect 21180 48136 21232 48142
rect 21180 48078 21232 48084
rect 20904 48068 20956 48074
rect 20904 48010 20956 48016
rect 20916 47802 20944 48010
rect 20904 47796 20956 47802
rect 22480 47784 22508 48282
rect 22480 47756 22600 47784
rect 20904 47738 20956 47744
rect 20904 47660 20956 47666
rect 20904 47602 20956 47608
rect 22468 47660 22520 47666
rect 22468 47602 22520 47608
rect 20916 47258 20944 47602
rect 20904 47252 20956 47258
rect 20904 47194 20956 47200
rect 22480 47122 22508 47602
rect 22468 47116 22520 47122
rect 22468 47058 22520 47064
rect 20996 46980 21048 46986
rect 20996 46922 21048 46928
rect 21008 46714 21036 46922
rect 20996 46708 21048 46714
rect 20996 46650 21048 46656
rect 22572 46578 22600 47756
rect 21088 46572 21140 46578
rect 21088 46514 21140 46520
rect 22560 46572 22612 46578
rect 22560 46514 22612 46520
rect 21100 46170 21128 46514
rect 21088 46164 21140 46170
rect 21088 46106 21140 46112
rect 22572 45966 22600 46514
rect 22560 45960 22612 45966
rect 22560 45902 22612 45908
rect 21272 45892 21324 45898
rect 21272 45834 21324 45840
rect 21284 45626 21312 45834
rect 21272 45620 21324 45626
rect 21272 45562 21324 45568
rect 20732 45526 20852 45554
rect 18052 45494 18104 45500
rect 19984 45484 20036 45490
rect 19984 45426 20036 45432
rect 17960 45348 18012 45354
rect 17960 45290 18012 45296
rect 19996 44946 20024 45426
rect 20260 45280 20312 45286
rect 20260 45222 20312 45228
rect 16672 44940 16724 44946
rect 16672 44882 16724 44888
rect 19984 44940 20036 44946
rect 19984 44882 20036 44888
rect 14096 44872 14148 44878
rect 14096 44814 14148 44820
rect 15476 44872 15528 44878
rect 15476 44814 15528 44820
rect 10784 44396 10836 44402
rect 10784 44338 10836 44344
rect 13636 44396 13688 44402
rect 13636 44338 13688 44344
rect 9496 44328 9548 44334
rect 11428 44328 11480 44334
rect 9548 44276 9628 44282
rect 9496 44270 9628 44276
rect 11428 44270 11480 44276
rect 9508 44254 9628 44270
rect 9508 44205 9536 44254
rect 9600 43790 9628 44254
rect 11440 43790 11468 44270
rect 14108 43858 14136 44814
rect 15476 44736 15528 44742
rect 15476 44678 15528 44684
rect 15488 44470 15516 44678
rect 15476 44464 15528 44470
rect 15476 44406 15528 44412
rect 16684 44402 16712 44882
rect 20272 44878 20300 45222
rect 20260 44872 20312 44878
rect 20260 44814 20312 44820
rect 18236 44736 18288 44742
rect 18236 44678 18288 44684
rect 18248 44470 18276 44678
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 18236 44464 18288 44470
rect 18236 44406 18288 44412
rect 16672 44396 16724 44402
rect 16672 44338 16724 44344
rect 14372 44192 14424 44198
rect 14372 44134 14424 44140
rect 14096 43852 14148 43858
rect 14096 43794 14148 43800
rect 7748 43784 7800 43790
rect 7748 43726 7800 43732
rect 9588 43784 9640 43790
rect 9588 43726 9640 43732
rect 11428 43784 11480 43790
rect 11428 43726 11480 43732
rect 7472 43444 7524 43450
rect 7472 43386 7524 43392
rect 5724 43376 5776 43382
rect 5724 43318 5776 43324
rect 6828 43376 6880 43382
rect 6828 43318 6880 43324
rect 6840 42770 6868 43318
rect 9600 43246 9628 43726
rect 9680 43716 9732 43722
rect 9680 43658 9732 43664
rect 10876 43716 10928 43722
rect 10876 43658 10928 43664
rect 9588 43240 9640 43246
rect 9588 43182 9640 43188
rect 9496 43104 9548 43110
rect 9496 43046 9548 43052
rect 6828 42764 6880 42770
rect 6828 42706 6880 42712
rect 6840 42226 6868 42706
rect 8300 42628 8352 42634
rect 8300 42570 8352 42576
rect 7656 42560 7708 42566
rect 7656 42502 7708 42508
rect 6828 42220 6880 42226
rect 6828 42162 6880 42168
rect 6840 41682 6868 42162
rect 6828 41676 6880 41682
rect 6828 41618 6880 41624
rect 7668 41206 7696 42502
rect 8312 41818 8340 42570
rect 8944 42152 8996 42158
rect 8944 42094 8996 42100
rect 8576 42016 8628 42022
rect 8576 41958 8628 41964
rect 8300 41812 8352 41818
rect 8300 41754 8352 41760
rect 8588 41614 8616 41958
rect 8576 41608 8628 41614
rect 8576 41550 8628 41556
rect 7656 41200 7708 41206
rect 7656 41142 7708 41148
rect 8956 41070 8984 42094
rect 9508 41206 9536 43046
rect 9600 42158 9628 43182
rect 9692 42702 9720 43658
rect 9680 42696 9732 42702
rect 9680 42638 9732 42644
rect 9588 42152 9640 42158
rect 9588 42094 9640 42100
rect 9496 41200 9548 41206
rect 9496 41142 9548 41148
rect 6460 41064 6512 41070
rect 6460 41006 6512 41012
rect 8944 41064 8996 41070
rect 8944 41006 8996 41012
rect 5816 40520 5868 40526
rect 5816 40462 5868 40468
rect 3792 40112 3844 40118
rect 3792 40054 3844 40060
rect 5632 40112 5684 40118
rect 5632 40054 5684 40060
rect 3804 39438 3832 40054
rect 3976 40044 4028 40050
rect 3976 39986 4028 39992
rect 3988 39642 4016 39986
rect 5828 39982 5856 40462
rect 6472 40050 6500 41006
rect 7840 40928 7892 40934
rect 7840 40870 7892 40876
rect 7852 40526 7880 40870
rect 8956 40526 8984 41006
rect 10600 40928 10652 40934
rect 10600 40870 10652 40876
rect 10612 40526 10640 40870
rect 10888 40730 10916 43658
rect 10968 43308 11020 43314
rect 10968 43250 11020 43256
rect 10980 42362 11008 43250
rect 11440 43246 11468 43726
rect 11520 43648 11572 43654
rect 11520 43590 11572 43596
rect 13544 43648 13596 43654
rect 13544 43590 13596 43596
rect 11428 43240 11480 43246
rect 11428 43182 11480 43188
rect 11440 42906 11468 43182
rect 11428 42900 11480 42906
rect 11428 42842 11480 42848
rect 11336 42696 11388 42702
rect 11336 42638 11388 42644
rect 10968 42356 11020 42362
rect 10968 42298 11020 42304
rect 11348 41750 11376 42638
rect 11336 41744 11388 41750
rect 11336 41686 11388 41692
rect 10876 40724 10928 40730
rect 10876 40666 10928 40672
rect 7840 40520 7892 40526
rect 7840 40462 7892 40468
rect 8944 40520 8996 40526
rect 8944 40462 8996 40468
rect 10600 40520 10652 40526
rect 10600 40462 10652 40468
rect 7564 40384 7616 40390
rect 7564 40326 7616 40332
rect 7576 40050 7604 40326
rect 6460 40044 6512 40050
rect 6460 39986 6512 39992
rect 7564 40044 7616 40050
rect 7564 39986 7616 39992
rect 7840 40044 7892 40050
rect 7840 39986 7892 39992
rect 5816 39976 5868 39982
rect 5816 39918 5868 39924
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 3976 39636 4028 39642
rect 3976 39578 4028 39584
rect 5828 39438 5856 39918
rect 7748 39840 7800 39846
rect 7748 39782 7800 39788
rect 7760 39438 7788 39782
rect 7852 39642 7880 39986
rect 8208 39976 8260 39982
rect 8260 39924 8340 39930
rect 8208 39918 8340 39924
rect 8220 39902 8340 39918
rect 7840 39636 7892 39642
rect 7840 39578 7892 39584
rect 8312 39506 8340 39902
rect 8392 39840 8444 39846
rect 8392 39782 8444 39788
rect 8300 39500 8352 39506
rect 8300 39442 8352 39448
rect 3792 39432 3844 39438
rect 3792 39374 3844 39380
rect 5816 39432 5868 39438
rect 5816 39374 5868 39380
rect 7748 39432 7800 39438
rect 7748 39374 7800 39380
rect 3804 38894 3832 39374
rect 4068 39364 4120 39370
rect 4068 39306 4120 39312
rect 6828 39364 6880 39370
rect 6828 39306 6880 39312
rect 3792 38888 3844 38894
rect 3792 38830 3844 38836
rect 4080 38010 4108 39306
rect 6840 38962 6868 39306
rect 8404 39030 8432 39782
rect 8956 39506 8984 40462
rect 11348 39642 11376 41686
rect 11440 41682 11468 42842
rect 11428 41676 11480 41682
rect 11428 41618 11480 41624
rect 11532 40526 11560 43590
rect 13360 43308 13412 43314
rect 13360 43250 13412 43256
rect 12624 43104 12676 43110
rect 12624 43046 12676 43052
rect 11612 42220 11664 42226
rect 11612 42162 11664 42168
rect 11624 41818 11652 42162
rect 11612 41812 11664 41818
rect 11612 41754 11664 41760
rect 12636 41614 12664 43046
rect 13372 42362 13400 43250
rect 13360 42356 13412 42362
rect 13360 42298 13412 42304
rect 13556 42294 13584 43590
rect 14108 43314 14136 43794
rect 14384 43790 14412 44134
rect 16684 43858 16712 44338
rect 18328 44192 18380 44198
rect 18328 44134 18380 44140
rect 16672 43852 16724 43858
rect 16672 43794 16724 43800
rect 17132 43852 17184 43858
rect 17132 43794 17184 43800
rect 14372 43784 14424 43790
rect 14372 43726 14424 43732
rect 14832 43716 14884 43722
rect 14832 43658 14884 43664
rect 14844 43450 14872 43658
rect 15476 43648 15528 43654
rect 15476 43590 15528 43596
rect 14832 43444 14884 43450
rect 14832 43386 14884 43392
rect 15488 43382 15516 43590
rect 15476 43376 15528 43382
rect 15476 43318 15528 43324
rect 17144 43314 17172 43794
rect 18340 43790 18368 44134
rect 18328 43784 18380 43790
rect 18328 43726 18380 43732
rect 20536 43716 20588 43722
rect 20536 43658 20588 43664
rect 18512 43648 18564 43654
rect 18512 43590 18564 43596
rect 18524 43382 18552 43590
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 20548 43450 20576 43658
rect 20536 43444 20588 43450
rect 20536 43386 20588 43392
rect 18512 43376 18564 43382
rect 18512 43318 18564 43324
rect 14096 43308 14148 43314
rect 14096 43250 14148 43256
rect 17132 43308 17184 43314
rect 17132 43250 17184 43256
rect 19248 43308 19300 43314
rect 19248 43250 19300 43256
rect 19340 43308 19392 43314
rect 19340 43250 19392 43256
rect 12808 42288 12860 42294
rect 12808 42230 12860 42236
rect 13544 42288 13596 42294
rect 13544 42230 13596 42236
rect 12624 41608 12676 41614
rect 12624 41550 12676 41556
rect 12164 41472 12216 41478
rect 12164 41414 12216 41420
rect 12176 41138 12204 41414
rect 12164 41132 12216 41138
rect 12164 41074 12216 41080
rect 11520 40520 11572 40526
rect 11520 40462 11572 40468
rect 12176 40458 12204 41074
rect 12820 40730 12848 42230
rect 14108 42226 14136 43250
rect 17144 42770 17172 43250
rect 18604 43104 18656 43110
rect 18604 43046 18656 43052
rect 18788 43104 18840 43110
rect 18788 43046 18840 43052
rect 17132 42764 17184 42770
rect 17132 42706 17184 42712
rect 18616 42702 18644 43046
rect 15292 42696 15344 42702
rect 15292 42638 15344 42644
rect 18604 42696 18656 42702
rect 18604 42638 18656 42644
rect 14096 42220 14148 42226
rect 14096 42162 14148 42168
rect 14108 41478 14136 42162
rect 14096 41472 14148 41478
rect 14096 41414 14148 41420
rect 14108 41206 14136 41414
rect 14096 41200 14148 41206
rect 14096 41142 14148 41148
rect 14108 41070 14136 41142
rect 14832 41132 14884 41138
rect 14832 41074 14884 41080
rect 14096 41064 14148 41070
rect 14096 41006 14148 41012
rect 14740 41064 14792 41070
rect 14740 41006 14792 41012
rect 14280 40928 14332 40934
rect 14280 40870 14332 40876
rect 12808 40724 12860 40730
rect 12808 40666 12860 40672
rect 12164 40452 12216 40458
rect 12164 40394 12216 40400
rect 12176 40050 12204 40394
rect 14292 40050 14320 40870
rect 14752 40050 14780 41006
rect 12164 40044 12216 40050
rect 12164 39986 12216 39992
rect 14280 40044 14332 40050
rect 14280 39986 14332 39992
rect 14740 40044 14792 40050
rect 14740 39986 14792 39992
rect 11336 39636 11388 39642
rect 11336 39578 11388 39584
rect 12176 39506 12204 39986
rect 13544 39840 13596 39846
rect 13544 39782 13596 39788
rect 8944 39500 8996 39506
rect 8944 39442 8996 39448
rect 12164 39500 12216 39506
rect 12164 39442 12216 39448
rect 8484 39364 8536 39370
rect 8484 39306 8536 39312
rect 8496 39098 8524 39306
rect 8484 39092 8536 39098
rect 8484 39034 8536 39040
rect 8392 39024 8444 39030
rect 8392 38966 8444 38972
rect 8956 38962 8984 39442
rect 10324 39296 10376 39302
rect 10324 39238 10376 39244
rect 10336 39030 10364 39238
rect 10324 39024 10376 39030
rect 10324 38966 10376 38972
rect 12176 38962 12204 39442
rect 13556 39438 13584 39782
rect 13544 39432 13596 39438
rect 13544 39374 13596 39380
rect 14752 39370 14780 39986
rect 13360 39364 13412 39370
rect 13360 39306 13412 39312
rect 14740 39364 14792 39370
rect 14740 39306 14792 39312
rect 5724 38956 5776 38962
rect 5724 38898 5776 38904
rect 6828 38956 6880 38962
rect 6828 38898 6880 38904
rect 8944 38956 8996 38962
rect 8944 38898 8996 38904
rect 12164 38956 12216 38962
rect 12164 38898 12216 38904
rect 4988 38752 5040 38758
rect 4988 38694 5040 38700
rect 5172 38752 5224 38758
rect 5172 38694 5224 38700
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 5000 38350 5028 38694
rect 4988 38344 5040 38350
rect 4988 38286 5040 38292
rect 4068 38004 4120 38010
rect 4068 37946 4120 37952
rect 4620 37664 4672 37670
rect 4620 37606 4672 37612
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4632 36802 4660 37606
rect 5000 37262 5028 38286
rect 5184 37874 5212 38694
rect 5736 38010 5764 38898
rect 5816 38276 5868 38282
rect 5816 38218 5868 38224
rect 5724 38004 5776 38010
rect 5724 37946 5776 37952
rect 5172 37868 5224 37874
rect 5172 37810 5224 37816
rect 4988 37256 5040 37262
rect 4988 37198 5040 37204
rect 5828 36922 5856 38218
rect 6368 38208 6420 38214
rect 6368 38150 6420 38156
rect 6380 37942 6408 38150
rect 6368 37936 6420 37942
rect 6368 37878 6420 37884
rect 6644 37800 6696 37806
rect 6644 37742 6696 37748
rect 6552 37120 6604 37126
rect 6552 37062 6604 37068
rect 5816 36916 5868 36922
rect 5816 36858 5868 36864
rect 6564 36854 6592 37062
rect 4540 36786 4660 36802
rect 6552 36848 6604 36854
rect 6552 36790 6604 36796
rect 6656 36786 6684 37742
rect 6840 37262 6868 38898
rect 10324 38752 10376 38758
rect 10324 38694 10376 38700
rect 10336 38350 10364 38694
rect 12176 38350 12204 38898
rect 8944 38344 8996 38350
rect 8944 38286 8996 38292
rect 10324 38344 10376 38350
rect 10324 38286 10376 38292
rect 12164 38344 12216 38350
rect 12164 38286 12216 38292
rect 8956 37330 8984 38286
rect 10324 38208 10376 38214
rect 10324 38150 10376 38156
rect 10336 37942 10364 38150
rect 10324 37936 10376 37942
rect 10324 37878 10376 37884
rect 11520 37800 11572 37806
rect 11520 37742 11572 37748
rect 9772 37664 9824 37670
rect 9772 37606 9824 37612
rect 8944 37324 8996 37330
rect 8944 37266 8996 37272
rect 6828 37256 6880 37262
rect 6828 37198 6880 37204
rect 8956 37210 8984 37266
rect 9784 37262 9812 37606
rect 11532 37262 11560 37742
rect 13176 37664 13228 37670
rect 13176 37606 13228 37612
rect 13188 37262 13216 37606
rect 9772 37256 9824 37262
rect 6736 37188 6788 37194
rect 8956 37182 9168 37210
rect 9772 37198 9824 37204
rect 11520 37256 11572 37262
rect 11520 37198 11572 37204
rect 13176 37256 13228 37262
rect 13176 37198 13228 37204
rect 6736 37130 6788 37136
rect 4528 36780 4660 36786
rect 4580 36774 4660 36780
rect 4988 36780 5040 36786
rect 4528 36722 4580 36728
rect 4988 36722 5040 36728
rect 6644 36780 6696 36786
rect 6644 36722 6696 36728
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 3976 35692 4028 35698
rect 3976 35634 4028 35640
rect 3988 34678 4016 35634
rect 5000 35494 5028 36722
rect 6656 36174 6684 36722
rect 6368 36168 6420 36174
rect 6368 36110 6420 36116
rect 6644 36168 6696 36174
rect 6644 36110 6696 36116
rect 6380 35630 6408 36110
rect 6748 35834 6776 37130
rect 9140 37126 9168 37182
rect 9680 37188 9732 37194
rect 9680 37130 9732 37136
rect 9036 37120 9088 37126
rect 9036 37062 9088 37068
rect 9128 37120 9180 37126
rect 9128 37062 9180 37068
rect 8484 36848 8536 36854
rect 8484 36790 8536 36796
rect 8392 36712 8444 36718
rect 8392 36654 8444 36660
rect 7932 36576 7984 36582
rect 7932 36518 7984 36524
rect 7944 36174 7972 36518
rect 8404 36242 8432 36654
rect 8496 36378 8524 36790
rect 8484 36372 8536 36378
rect 8484 36314 8536 36320
rect 8392 36236 8444 36242
rect 8392 36178 8444 36184
rect 8944 36236 8996 36242
rect 8944 36178 8996 36184
rect 7932 36168 7984 36174
rect 7932 36110 7984 36116
rect 7932 36032 7984 36038
rect 7932 35974 7984 35980
rect 6736 35828 6788 35834
rect 6736 35770 6788 35776
rect 7944 35766 7972 35974
rect 7932 35760 7984 35766
rect 7932 35702 7984 35708
rect 6368 35624 6420 35630
rect 6368 35566 6420 35572
rect 4988 35488 5040 35494
rect 4988 35430 5040 35436
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 3976 34672 4028 34678
rect 3976 34614 4028 34620
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 3792 33992 3844 33998
rect 3792 33934 3844 33940
rect 3804 33454 3832 33934
rect 3792 33448 3844 33454
rect 3792 33390 3844 33396
rect 3804 32910 3832 33390
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 3792 32904 3844 32910
rect 3792 32846 3844 32852
rect 4712 32836 4764 32842
rect 4712 32778 4764 32784
rect 4724 32570 4752 32778
rect 4712 32564 4764 32570
rect 4712 32506 4764 32512
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 5000 32026 5028 35430
rect 6380 34474 6408 35566
rect 6828 35148 6880 35154
rect 6828 35090 6880 35096
rect 6840 34474 6868 35090
rect 8300 34944 8352 34950
rect 8300 34886 8352 34892
rect 6368 34468 6420 34474
rect 6368 34410 6420 34416
rect 6828 34468 6880 34474
rect 6828 34410 6880 34416
rect 6380 33998 6408 34410
rect 6368 33992 6420 33998
rect 6368 33934 6420 33940
rect 6000 33924 6052 33930
rect 6000 33866 6052 33872
rect 5172 33516 5224 33522
rect 5172 33458 5224 33464
rect 5184 33114 5212 33458
rect 5908 33312 5960 33318
rect 5908 33254 5960 33260
rect 5172 33108 5224 33114
rect 5172 33050 5224 33056
rect 5920 32842 5948 33254
rect 6012 33114 6040 33866
rect 6276 33856 6328 33862
rect 6276 33798 6328 33804
rect 6288 33590 6316 33798
rect 6276 33584 6328 33590
rect 6276 33526 6328 33532
rect 6380 33522 6408 33934
rect 7748 33924 7800 33930
rect 7748 33866 7800 33872
rect 7760 33658 7788 33866
rect 8116 33856 8168 33862
rect 8116 33798 8168 33804
rect 7748 33652 7800 33658
rect 7748 33594 7800 33600
rect 6368 33516 6420 33522
rect 6368 33458 6420 33464
rect 6920 33516 6972 33522
rect 6920 33458 6972 33464
rect 6000 33108 6052 33114
rect 6000 33050 6052 33056
rect 6932 32842 6960 33458
rect 5908 32836 5960 32842
rect 5908 32778 5960 32784
rect 6920 32836 6972 32842
rect 6920 32778 6972 32784
rect 6932 32434 6960 32778
rect 8128 32502 8156 33798
rect 8312 32502 8340 34886
rect 8956 34610 8984 36178
rect 9048 36174 9076 37062
rect 9692 36922 9720 37130
rect 10324 37120 10376 37126
rect 10324 37062 10376 37068
rect 9680 36916 9732 36922
rect 9680 36858 9732 36864
rect 10336 36854 10364 37062
rect 10324 36848 10376 36854
rect 10324 36790 10376 36796
rect 11532 36786 11560 37198
rect 12900 37120 12952 37126
rect 12900 37062 12952 37068
rect 12912 36854 12940 37062
rect 13372 36854 13400 39306
rect 14844 39302 14872 41074
rect 15304 40594 15332 42638
rect 16028 42628 16080 42634
rect 16028 42570 16080 42576
rect 16040 41002 16068 42570
rect 16856 42560 16908 42566
rect 16856 42502 16908 42508
rect 18696 42560 18748 42566
rect 18696 42502 18748 42508
rect 16120 42016 16172 42022
rect 16120 41958 16172 41964
rect 16132 41206 16160 41958
rect 16120 41200 16172 41206
rect 16120 41142 16172 41148
rect 16028 40996 16080 41002
rect 16028 40938 16080 40944
rect 15292 40588 15344 40594
rect 15292 40530 15344 40536
rect 16868 40526 16896 42502
rect 18708 42294 18736 42502
rect 18696 42288 18748 42294
rect 18696 42230 18748 42236
rect 18604 42220 18656 42226
rect 18604 42162 18656 42168
rect 17316 42152 17368 42158
rect 17316 42094 17368 42100
rect 17328 41614 17356 42094
rect 17316 41608 17368 41614
rect 17316 41550 17368 41556
rect 17328 41070 17356 41550
rect 17316 41064 17368 41070
rect 17316 41006 17368 41012
rect 17328 40526 17356 41006
rect 18616 40730 18644 42162
rect 18800 41614 18828 43046
rect 19260 42838 19288 43250
rect 19248 42832 19300 42838
rect 19248 42774 19300 42780
rect 19352 42362 19380 43250
rect 19984 42764 20036 42770
rect 19984 42706 20036 42712
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 19340 42356 19392 42362
rect 19340 42298 19392 42304
rect 19996 42226 20024 42706
rect 19984 42220 20036 42226
rect 19984 42162 20036 42168
rect 19996 41682 20024 42162
rect 19984 41676 20036 41682
rect 19984 41618 20036 41624
rect 18788 41608 18840 41614
rect 18788 41550 18840 41556
rect 18696 41472 18748 41478
rect 18696 41414 18748 41420
rect 18708 41206 18736 41414
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 18696 41200 18748 41206
rect 18696 41142 18748 41148
rect 19996 41138 20024 41618
rect 19984 41132 20036 41138
rect 19984 41074 20036 41080
rect 19064 40928 19116 40934
rect 19064 40870 19116 40876
rect 18604 40724 18656 40730
rect 18604 40666 18656 40672
rect 19076 40526 19104 40870
rect 16856 40520 16908 40526
rect 16856 40462 16908 40468
rect 17316 40520 17368 40526
rect 17316 40462 17368 40468
rect 19064 40520 19116 40526
rect 19064 40462 19116 40468
rect 15292 40384 15344 40390
rect 15292 40326 15344 40332
rect 15304 40050 15332 40326
rect 17328 40118 17356 40462
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19340 40180 19392 40186
rect 19340 40122 19392 40128
rect 17316 40112 17368 40118
rect 17316 40054 17368 40060
rect 15292 40044 15344 40050
rect 15292 39986 15344 39992
rect 16120 39840 16172 39846
rect 16120 39782 16172 39788
rect 16132 39438 16160 39782
rect 17328 39438 17356 40054
rect 18052 40044 18104 40050
rect 18052 39986 18104 39992
rect 18064 39642 18092 39986
rect 18052 39636 18104 39642
rect 18052 39578 18104 39584
rect 19352 39438 19380 40122
rect 19996 40050 20024 41074
rect 20548 40458 20576 43386
rect 20536 40452 20588 40458
rect 20536 40394 20588 40400
rect 19984 40044 20036 40050
rect 19984 39986 20036 39992
rect 16120 39432 16172 39438
rect 16120 39374 16172 39380
rect 17316 39432 17368 39438
rect 17316 39374 17368 39380
rect 18512 39432 18564 39438
rect 18512 39374 18564 39380
rect 19340 39432 19392 39438
rect 19340 39374 19392 39380
rect 18328 39364 18380 39370
rect 18328 39306 18380 39312
rect 13544 39296 13596 39302
rect 13544 39238 13596 39244
rect 14832 39296 14884 39302
rect 14832 39238 14884 39244
rect 13556 39030 13584 39238
rect 18340 39098 18368 39306
rect 18328 39092 18380 39098
rect 18328 39034 18380 39040
rect 13544 39024 13596 39030
rect 13544 38966 13596 38972
rect 18052 38956 18104 38962
rect 18052 38898 18104 38904
rect 16672 38888 16724 38894
rect 16672 38830 16724 38836
rect 13544 38752 13596 38758
rect 13544 38694 13596 38700
rect 13556 38350 13584 38694
rect 13544 38344 13596 38350
rect 13544 38286 13596 38292
rect 14740 38344 14792 38350
rect 14740 38286 14792 38292
rect 13452 38208 13504 38214
rect 13452 38150 13504 38156
rect 13464 37942 13492 38150
rect 13452 37936 13504 37942
rect 13452 37878 13504 37884
rect 14752 37330 14780 38286
rect 15844 38276 15896 38282
rect 15844 38218 15896 38224
rect 15856 38010 15884 38218
rect 15844 38004 15896 38010
rect 15844 37946 15896 37952
rect 15292 37868 15344 37874
rect 15292 37810 15344 37816
rect 15304 37346 15332 37810
rect 16684 37806 16712 38830
rect 17960 38276 18012 38282
rect 17960 38218 18012 38224
rect 16948 38208 17000 38214
rect 16948 38150 17000 38156
rect 17868 38208 17920 38214
rect 17868 38150 17920 38156
rect 16672 37800 16724 37806
rect 16672 37742 16724 37748
rect 14740 37324 14792 37330
rect 15304 37318 15424 37346
rect 14740 37266 14792 37272
rect 14752 36922 14780 37266
rect 15292 37188 15344 37194
rect 15292 37130 15344 37136
rect 14740 36916 14792 36922
rect 14740 36858 14792 36864
rect 12900 36848 12952 36854
rect 12900 36790 12952 36796
rect 13360 36848 13412 36854
rect 13360 36790 13412 36796
rect 11520 36780 11572 36786
rect 11520 36722 11572 36728
rect 11532 36242 11560 36722
rect 12900 36576 12952 36582
rect 12900 36518 12952 36524
rect 11520 36236 11572 36242
rect 11520 36178 11572 36184
rect 9036 36168 9088 36174
rect 9036 36110 9088 36116
rect 11532 35698 11560 36178
rect 12912 36174 12940 36518
rect 12900 36168 12952 36174
rect 12900 36110 12952 36116
rect 12900 36032 12952 36038
rect 12900 35974 12952 35980
rect 12912 35766 12940 35974
rect 12900 35760 12952 35766
rect 12900 35702 12952 35708
rect 11520 35692 11572 35698
rect 11520 35634 11572 35640
rect 11532 35154 11560 35634
rect 12900 35488 12952 35494
rect 12900 35430 12952 35436
rect 11520 35148 11572 35154
rect 11520 35090 11572 35096
rect 12912 35086 12940 35430
rect 12900 35080 12952 35086
rect 12900 35022 12952 35028
rect 9588 35012 9640 35018
rect 9588 34954 9640 34960
rect 8944 34604 8996 34610
rect 8944 34546 8996 34552
rect 8956 34066 8984 34546
rect 8944 34060 8996 34066
rect 8944 34002 8996 34008
rect 8576 33584 8628 33590
rect 8576 33526 8628 33532
rect 8588 32570 8616 33526
rect 8956 33522 8984 34002
rect 9600 33658 9628 34954
rect 11060 34740 11112 34746
rect 11060 34682 11112 34688
rect 10324 34604 10376 34610
rect 10324 34546 10376 34552
rect 10336 34202 10364 34546
rect 10784 34536 10836 34542
rect 10784 34478 10836 34484
rect 10324 34196 10376 34202
rect 10324 34138 10376 34144
rect 10796 33998 10824 34478
rect 10784 33992 10836 33998
rect 10784 33934 10836 33940
rect 10324 33924 10376 33930
rect 10324 33866 10376 33872
rect 9588 33652 9640 33658
rect 9588 33594 9640 33600
rect 8944 33516 8996 33522
rect 8944 33458 8996 33464
rect 8956 32978 8984 33458
rect 10336 33114 10364 33866
rect 10324 33108 10376 33114
rect 10324 33050 10376 33056
rect 8944 32972 8996 32978
rect 8944 32914 8996 32920
rect 11072 32910 11100 34682
rect 11888 34672 11940 34678
rect 11888 34614 11940 34620
rect 11900 33590 11928 34614
rect 13084 34536 13136 34542
rect 13084 34478 13136 34484
rect 12072 33924 12124 33930
rect 12072 33866 12124 33872
rect 11888 33584 11940 33590
rect 11888 33526 11940 33532
rect 12084 33114 12112 33866
rect 12532 33856 12584 33862
rect 12532 33798 12584 33804
rect 12072 33108 12124 33114
rect 12072 33050 12124 33056
rect 10232 32904 10284 32910
rect 10232 32846 10284 32852
rect 11060 32904 11112 32910
rect 11060 32846 11112 32852
rect 9588 32836 9640 32842
rect 9588 32778 9640 32784
rect 9600 32570 9628 32778
rect 8576 32564 8628 32570
rect 8576 32506 8628 32512
rect 9588 32564 9640 32570
rect 9588 32506 9640 32512
rect 8116 32496 8168 32502
rect 8116 32438 8168 32444
rect 8300 32496 8352 32502
rect 8300 32438 8352 32444
rect 5172 32428 5224 32434
rect 5172 32370 5224 32376
rect 6920 32428 6972 32434
rect 6920 32370 6972 32376
rect 5184 32026 5212 32370
rect 4988 32020 5040 32026
rect 4988 31962 5040 31968
rect 5172 32020 5224 32026
rect 5172 31962 5224 31968
rect 10244 31890 10272 32846
rect 12544 32502 12572 33798
rect 13096 33318 13124 34478
rect 13372 33590 13400 36790
rect 14752 36174 14780 36858
rect 14004 36168 14056 36174
rect 14004 36110 14056 36116
rect 14740 36168 14792 36174
rect 14740 36110 14792 36116
rect 13820 36100 13872 36106
rect 13820 36042 13872 36048
rect 13452 35692 13504 35698
rect 13452 35634 13504 35640
rect 13464 34746 13492 35634
rect 13636 35488 13688 35494
rect 13636 35430 13688 35436
rect 13452 34740 13504 34746
rect 13452 34682 13504 34688
rect 13648 34678 13676 35430
rect 13832 35290 13860 36042
rect 14016 35766 14044 36110
rect 15200 36032 15252 36038
rect 15200 35974 15252 35980
rect 14004 35760 14056 35766
rect 14004 35702 14056 35708
rect 13820 35284 13872 35290
rect 13820 35226 13872 35232
rect 14016 35086 14044 35702
rect 14004 35080 14056 35086
rect 14004 35022 14056 35028
rect 13636 34672 13688 34678
rect 13636 34614 13688 34620
rect 14016 33998 14044 35022
rect 14740 35012 14792 35018
rect 14740 34954 14792 34960
rect 14752 34746 14780 34954
rect 14740 34740 14792 34746
rect 14740 34682 14792 34688
rect 15212 34610 15240 35974
rect 15200 34604 15252 34610
rect 15200 34546 15252 34552
rect 15304 34202 15332 37130
rect 15292 34196 15344 34202
rect 15292 34138 15344 34144
rect 14004 33992 14056 33998
rect 14004 33934 14056 33940
rect 13360 33584 13412 33590
rect 13360 33526 13412 33532
rect 14016 33454 14044 33934
rect 14740 33516 14792 33522
rect 14740 33458 14792 33464
rect 14004 33448 14056 33454
rect 14004 33390 14056 33396
rect 13084 33312 13136 33318
rect 13084 33254 13136 33260
rect 12532 32496 12584 32502
rect 12532 32438 12584 32444
rect 13096 32434 13124 33254
rect 14016 32978 14044 33390
rect 14004 32972 14056 32978
rect 14004 32914 14056 32920
rect 13084 32428 13136 32434
rect 13084 32370 13136 32376
rect 13820 32428 13872 32434
rect 13820 32370 13872 32376
rect 12072 32360 12124 32366
rect 12072 32302 12124 32308
rect 10508 32224 10560 32230
rect 10508 32166 10560 32172
rect 10232 31884 10284 31890
rect 10232 31826 10284 31832
rect 10520 31822 10548 32166
rect 12084 31822 12112 32302
rect 13096 31890 13124 32370
rect 13084 31884 13136 31890
rect 13084 31826 13136 31832
rect 10508 31816 10560 31822
rect 10508 31758 10560 31764
rect 11520 31816 11572 31822
rect 11520 31758 11572 31764
rect 12072 31816 12124 31822
rect 12072 31758 12124 31764
rect 4252 31748 4304 31754
rect 4252 31690 4304 31696
rect 4264 31482 4292 31690
rect 4252 31476 4304 31482
rect 4252 31418 4304 31424
rect 3700 31408 3752 31414
rect 3700 31350 3752 31356
rect 11532 31346 11560 31758
rect 2872 31340 2924 31346
rect 2872 31282 2924 31288
rect 3976 31340 4028 31346
rect 3976 31282 4028 31288
rect 11520 31340 11572 31346
rect 11520 31282 11572 31288
rect 3988 30394 4016 31282
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 11532 30802 11560 31282
rect 13096 31278 13124 31826
rect 13452 31680 13504 31686
rect 13452 31622 13504 31628
rect 13464 31346 13492 31622
rect 13452 31340 13504 31346
rect 13452 31282 13504 31288
rect 13084 31272 13136 31278
rect 13084 31214 13136 31220
rect 12900 31136 12952 31142
rect 12900 31078 12952 31084
rect 11520 30796 11572 30802
rect 11520 30738 11572 30744
rect 12912 30734 12940 31078
rect 13832 30938 13860 32370
rect 13912 32224 13964 32230
rect 13912 32166 13964 32172
rect 13924 31346 13952 32166
rect 13912 31340 13964 31346
rect 13912 31282 13964 31288
rect 13820 30932 13872 30938
rect 13820 30874 13872 30880
rect 4528 30728 4580 30734
rect 4528 30670 4580 30676
rect 7012 30728 7064 30734
rect 7012 30670 7064 30676
rect 9312 30728 9364 30734
rect 9312 30670 9364 30676
rect 12900 30728 12952 30734
rect 12900 30670 12952 30676
rect 3976 30388 4028 30394
rect 3976 30330 4028 30336
rect 4540 30258 4568 30670
rect 5816 30660 5868 30666
rect 5816 30602 5868 30608
rect 5264 30592 5316 30598
rect 5264 30534 5316 30540
rect 3976 30252 4028 30258
rect 3976 30194 4028 30200
rect 4528 30252 4580 30258
rect 4528 30194 4580 30200
rect 3988 29306 4016 30194
rect 4540 30138 4568 30194
rect 4540 30110 4660 30138
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4632 29578 4660 30110
rect 4436 29572 4488 29578
rect 4436 29514 4488 29520
rect 4620 29572 4672 29578
rect 4620 29514 4672 29520
rect 4988 29572 5040 29578
rect 4988 29514 5040 29520
rect 3976 29300 4028 29306
rect 3976 29242 4028 29248
rect 4448 29170 4476 29514
rect 4436 29164 4488 29170
rect 4436 29106 4488 29112
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 5000 28626 5028 29514
rect 5276 29238 5304 30534
rect 5828 30394 5856 30602
rect 6184 30592 6236 30598
rect 6184 30534 6236 30540
rect 5816 30388 5868 30394
rect 5816 30330 5868 30336
rect 5816 30252 5868 30258
rect 5816 30194 5868 30200
rect 5828 29306 5856 30194
rect 6196 29646 6224 30534
rect 7024 30274 7052 30670
rect 8208 30660 8260 30666
rect 8208 30602 8260 30608
rect 6932 30246 7052 30274
rect 6932 30190 6960 30246
rect 6920 30184 6972 30190
rect 6920 30126 6972 30132
rect 6184 29640 6236 29646
rect 6184 29582 6236 29588
rect 6932 29578 6960 30126
rect 6920 29572 6972 29578
rect 6920 29514 6972 29520
rect 6552 29504 6604 29510
rect 6552 29446 6604 29452
rect 5816 29300 5868 29306
rect 5816 29242 5868 29248
rect 5264 29232 5316 29238
rect 5264 29174 5316 29180
rect 6368 29164 6420 29170
rect 6368 29106 6420 29112
rect 6380 28762 6408 29106
rect 6368 28756 6420 28762
rect 6368 28698 6420 28704
rect 4988 28620 5040 28626
rect 4988 28562 5040 28568
rect 6564 28558 6592 29446
rect 6932 29034 6960 29514
rect 7104 29504 7156 29510
rect 7104 29446 7156 29452
rect 6920 29028 6972 29034
rect 6920 28970 6972 28976
rect 6552 28552 6604 28558
rect 6552 28494 6604 28500
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 6932 27470 6960 28970
rect 7116 27470 7144 29446
rect 8220 27606 8248 30602
rect 8392 30252 8444 30258
rect 8392 30194 8444 30200
rect 8404 28762 8432 30194
rect 9324 30190 9352 30670
rect 10968 30660 11020 30666
rect 10968 30602 11020 30608
rect 9680 30592 9732 30598
rect 9680 30534 9732 30540
rect 9312 30184 9364 30190
rect 9312 30126 9364 30132
rect 9588 30184 9640 30190
rect 9588 30126 9640 30132
rect 9128 30048 9180 30054
rect 9128 29990 9180 29996
rect 9140 29646 9168 29990
rect 9600 29646 9628 30126
rect 9128 29640 9180 29646
rect 9128 29582 9180 29588
rect 9588 29640 9640 29646
rect 9588 29582 9640 29588
rect 9600 29102 9628 29582
rect 9588 29096 9640 29102
rect 9588 29038 9640 29044
rect 8392 28756 8444 28762
rect 8392 28698 8444 28704
rect 8300 28552 8352 28558
rect 8300 28494 8352 28500
rect 8312 28082 8340 28494
rect 9128 28484 9180 28490
rect 9128 28426 9180 28432
rect 9140 28218 9168 28426
rect 9128 28212 9180 28218
rect 9128 28154 9180 28160
rect 8300 28076 8352 28082
rect 8300 28018 8352 28024
rect 9600 28014 9628 29038
rect 9692 28150 9720 30534
rect 10980 30394 11008 30602
rect 10968 30388 11020 30394
rect 10968 30330 11020 30336
rect 14016 30258 14044 32914
rect 14752 31482 14780 33458
rect 14740 31476 14792 31482
rect 14740 31418 14792 31424
rect 14096 30728 14148 30734
rect 14096 30670 14148 30676
rect 10876 30252 10928 30258
rect 10876 30194 10928 30200
rect 11520 30252 11572 30258
rect 11520 30194 11572 30200
rect 13268 30252 13320 30258
rect 13268 30194 13320 30200
rect 14004 30252 14056 30258
rect 14004 30194 14056 30200
rect 10888 29306 10916 30194
rect 11532 29714 11560 30194
rect 12440 30048 12492 30054
rect 12440 29990 12492 29996
rect 11520 29708 11572 29714
rect 11520 29650 11572 29656
rect 10968 29572 11020 29578
rect 10968 29514 11020 29520
rect 10876 29300 10928 29306
rect 10876 29242 10928 29248
rect 10692 29164 10744 29170
rect 10692 29106 10744 29112
rect 10704 28558 10732 29106
rect 10692 28552 10744 28558
rect 10692 28494 10744 28500
rect 10980 28218 11008 29514
rect 11428 29504 11480 29510
rect 11428 29446 11480 29452
rect 11440 29238 11468 29446
rect 11428 29232 11480 29238
rect 11428 29174 11480 29180
rect 11532 28762 11560 29650
rect 11520 28756 11572 28762
rect 11520 28698 11572 28704
rect 10968 28212 11020 28218
rect 10968 28154 11020 28160
rect 12452 28150 12480 29990
rect 13280 29850 13308 30194
rect 13268 29844 13320 29850
rect 13268 29786 13320 29792
rect 13544 29572 13596 29578
rect 13544 29514 13596 29520
rect 12532 28552 12584 28558
rect 12532 28494 12584 28500
rect 9680 28144 9732 28150
rect 9680 28086 9732 28092
rect 12440 28144 12492 28150
rect 12440 28086 12492 28092
rect 12256 28076 12308 28082
rect 12256 28018 12308 28024
rect 9588 28008 9640 28014
rect 9588 27950 9640 27956
rect 8208 27600 8260 27606
rect 8208 27542 8260 27548
rect 6920 27464 6972 27470
rect 6920 27406 6972 27412
rect 7104 27464 7156 27470
rect 7104 27406 7156 27412
rect 6932 26994 6960 27406
rect 6920 26988 6972 26994
rect 6920 26930 6972 26936
rect 8484 26988 8536 26994
rect 8484 26930 8536 26936
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 6932 26586 6960 26930
rect 6920 26580 6972 26586
rect 6920 26522 6972 26528
rect 6932 25906 6960 26522
rect 8024 26240 8076 26246
rect 8024 26182 8076 26188
rect 8036 25974 8064 26182
rect 8496 26042 8524 26930
rect 9036 26784 9088 26790
rect 9036 26726 9088 26732
rect 9128 26784 9180 26790
rect 9128 26726 9180 26732
rect 8484 26036 8536 26042
rect 8484 25978 8536 25984
rect 9048 25974 9076 26726
rect 9140 26382 9168 26726
rect 9128 26376 9180 26382
rect 9128 26318 9180 26324
rect 8024 25968 8076 25974
rect 8024 25910 8076 25916
rect 9036 25968 9088 25974
rect 9036 25910 9088 25916
rect 9600 25906 9628 27950
rect 12268 27470 12296 28018
rect 12256 27464 12308 27470
rect 12256 27406 12308 27412
rect 12268 27062 12296 27406
rect 12544 27062 12572 28494
rect 13556 27606 13584 29514
rect 14108 29170 14136 30670
rect 15396 30122 15424 37318
rect 16684 37262 16712 37742
rect 16960 37262 16988 38150
rect 17880 37942 17908 38150
rect 17868 37936 17920 37942
rect 17868 37878 17920 37884
rect 17972 37466 18000 38218
rect 18064 38010 18092 38898
rect 18524 38894 18552 39374
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 18512 38888 18564 38894
rect 18512 38830 18564 38836
rect 18524 38282 18552 38830
rect 20548 38758 20576 40394
rect 20824 39642 20852 45526
rect 21364 45484 21416 45490
rect 21364 45426 21416 45432
rect 21376 45082 21404 45426
rect 21824 45416 21876 45422
rect 21824 45358 21876 45364
rect 21364 45076 21416 45082
rect 21364 45018 21416 45024
rect 21548 44872 21600 44878
rect 21548 44814 21600 44820
rect 21560 43790 21588 44814
rect 21836 44402 21864 45358
rect 23032 44878 23060 52566
rect 24872 52562 24900 53042
rect 26252 52698 26280 53042
rect 26792 52896 26844 52902
rect 26792 52838 26844 52844
rect 26240 52692 26292 52698
rect 26240 52634 26292 52640
rect 24860 52556 24912 52562
rect 24860 52498 24912 52504
rect 23756 52488 23808 52494
rect 23756 52430 23808 52436
rect 23204 52012 23256 52018
rect 23204 51954 23256 51960
rect 23216 51066 23244 51954
rect 23664 51944 23716 51950
rect 23664 51886 23716 51892
rect 23480 51264 23532 51270
rect 23480 51206 23532 51212
rect 23204 51060 23256 51066
rect 23204 51002 23256 51008
rect 23112 50924 23164 50930
rect 23112 50866 23164 50872
rect 23124 50522 23152 50866
rect 23112 50516 23164 50522
rect 23112 50458 23164 50464
rect 23492 49910 23520 51206
rect 23676 50930 23704 51886
rect 23664 50924 23716 50930
rect 23664 50866 23716 50872
rect 23676 50726 23704 50866
rect 23664 50720 23716 50726
rect 23664 50662 23716 50668
rect 23480 49904 23532 49910
rect 23480 49846 23532 49852
rect 23112 49088 23164 49094
rect 23112 49030 23164 49036
rect 23124 45966 23152 49030
rect 23768 46170 23796 52430
rect 24872 52426 24900 52498
rect 26804 52494 26832 52838
rect 25688 52488 25740 52494
rect 25688 52430 25740 52436
rect 26792 52488 26844 52494
rect 26792 52430 26844 52436
rect 24860 52420 24912 52426
rect 24860 52362 24912 52368
rect 24492 52012 24544 52018
rect 24492 51954 24544 51960
rect 23940 51808 23992 51814
rect 23940 51750 23992 51756
rect 23952 50998 23980 51750
rect 23940 50992 23992 50998
rect 23940 50934 23992 50940
rect 24504 49978 24532 51954
rect 24872 51626 24900 52362
rect 24952 51808 25004 51814
rect 24952 51750 25004 51756
rect 24780 51610 24900 51626
rect 24768 51604 24900 51610
rect 24820 51598 24900 51604
rect 24768 51546 24820 51552
rect 24964 50318 24992 51750
rect 25044 51332 25096 51338
rect 25044 51274 25096 51280
rect 25056 51066 25084 51274
rect 25044 51060 25096 51066
rect 25044 51002 25096 51008
rect 25700 50522 25728 52430
rect 26976 52352 27028 52358
rect 26976 52294 27028 52300
rect 26988 51950 27016 52294
rect 26976 51944 27028 51950
rect 26976 51886 27028 51892
rect 25780 51400 25832 51406
rect 25780 51342 25832 51348
rect 25688 50516 25740 50522
rect 25688 50458 25740 50464
rect 24952 50312 25004 50318
rect 24952 50254 25004 50260
rect 24860 50244 24912 50250
rect 24860 50186 24912 50192
rect 24492 49972 24544 49978
rect 24492 49914 24544 49920
rect 24872 49842 24900 50186
rect 24860 49836 24912 49842
rect 24860 49778 24912 49784
rect 24872 49298 24900 49778
rect 24860 49292 24912 49298
rect 24860 49234 24912 49240
rect 24032 49156 24084 49162
rect 24032 49098 24084 49104
rect 23848 48544 23900 48550
rect 23848 48486 23900 48492
rect 23860 47054 23888 48486
rect 23848 47048 23900 47054
rect 23848 46990 23900 46996
rect 23848 46912 23900 46918
rect 23848 46854 23900 46860
rect 23860 46646 23888 46854
rect 24044 46714 24072 49098
rect 24872 48754 24900 49234
rect 24400 48748 24452 48754
rect 24400 48690 24452 48696
rect 24860 48748 24912 48754
rect 24860 48690 24912 48696
rect 24412 47802 24440 48690
rect 24872 48346 24900 48690
rect 24860 48340 24912 48346
rect 24860 48282 24912 48288
rect 24400 47796 24452 47802
rect 24400 47738 24452 47744
rect 24872 47666 24900 48282
rect 25792 48142 25820 51342
rect 26988 50862 27016 51886
rect 27632 51406 27660 56374
rect 28356 56364 28408 56370
rect 28356 56306 28408 56312
rect 28264 56296 28316 56302
rect 28264 56238 28316 56244
rect 28276 55350 28304 56238
rect 28368 55622 28396 56306
rect 28356 55616 28408 55622
rect 28356 55558 28408 55564
rect 28264 55344 28316 55350
rect 28264 55286 28316 55292
rect 28172 55276 28224 55282
rect 28172 55218 28224 55224
rect 28184 54874 28212 55218
rect 28172 54868 28224 54874
rect 28172 54810 28224 54816
rect 28356 54596 28408 54602
rect 28356 54538 28408 54544
rect 28368 54330 28396 54538
rect 28356 54324 28408 54330
rect 28356 54266 28408 54272
rect 28080 52352 28132 52358
rect 28080 52294 28132 52300
rect 28092 52086 28120 52294
rect 28080 52080 28132 52086
rect 28080 52022 28132 52028
rect 28356 51808 28408 51814
rect 28356 51750 28408 51756
rect 27620 51400 27672 51406
rect 27620 51342 27672 51348
rect 28368 50998 28396 51750
rect 28356 50992 28408 50998
rect 28356 50934 28408 50940
rect 26976 50856 27028 50862
rect 26976 50798 27028 50804
rect 26988 50318 27016 50798
rect 28356 50720 28408 50726
rect 28356 50662 28408 50668
rect 28368 50318 28396 50662
rect 26976 50312 27028 50318
rect 26976 50254 27028 50260
rect 28356 50312 28408 50318
rect 28356 50254 28408 50260
rect 26240 49972 26292 49978
rect 26240 49914 26292 49920
rect 25780 48136 25832 48142
rect 25780 48078 25832 48084
rect 26252 47734 26280 49914
rect 26988 49842 27016 50254
rect 28356 50176 28408 50182
rect 28356 50118 28408 50124
rect 28368 49910 28396 50118
rect 28356 49904 28408 49910
rect 28356 49846 28408 49852
rect 26424 49836 26476 49842
rect 26424 49778 26476 49784
rect 26976 49836 27028 49842
rect 26976 49778 27028 49784
rect 26436 49434 26464 49778
rect 26424 49428 26476 49434
rect 26424 49370 26476 49376
rect 26332 49156 26384 49162
rect 26332 49098 26384 49104
rect 26344 48890 26372 49098
rect 26332 48884 26384 48890
rect 26332 48826 26384 48832
rect 26424 48748 26476 48754
rect 26424 48690 26476 48696
rect 26436 47802 26464 48690
rect 26424 47796 26476 47802
rect 26424 47738 26476 47744
rect 26240 47728 26292 47734
rect 26240 47670 26292 47676
rect 24860 47660 24912 47666
rect 24860 47602 24912 47608
rect 26792 47660 26844 47666
rect 26792 47602 26844 47608
rect 24872 47122 24900 47602
rect 26804 47258 26832 47602
rect 27620 47592 27672 47598
rect 27620 47534 27672 47540
rect 26792 47252 26844 47258
rect 26792 47194 26844 47200
rect 27632 47122 27660 47534
rect 24860 47116 24912 47122
rect 24860 47058 24912 47064
rect 27620 47116 27672 47122
rect 27620 47058 27672 47064
rect 24032 46708 24084 46714
rect 24032 46650 24084 46656
rect 23848 46640 23900 46646
rect 23848 46582 23900 46588
rect 24872 46578 24900 47058
rect 26424 46980 26476 46986
rect 26424 46922 26476 46928
rect 26436 46714 26464 46922
rect 26424 46708 26476 46714
rect 26424 46650 26476 46656
rect 24860 46572 24912 46578
rect 24860 46514 24912 46520
rect 26240 46572 26292 46578
rect 26240 46514 26292 46520
rect 23756 46164 23808 46170
rect 23756 46106 23808 46112
rect 24872 46034 24900 46514
rect 26252 46170 26280 46514
rect 26240 46164 26292 46170
rect 26240 46106 26292 46112
rect 27632 46034 27660 47058
rect 24860 46028 24912 46034
rect 24860 45970 24912 45976
rect 27620 46028 27672 46034
rect 27620 45970 27672 45976
rect 23112 45960 23164 45966
rect 23112 45902 23164 45908
rect 24952 45892 25004 45898
rect 24952 45834 25004 45840
rect 23204 45484 23256 45490
rect 23204 45426 23256 45432
rect 23216 45082 23244 45426
rect 23204 45076 23256 45082
rect 23204 45018 23256 45024
rect 23020 44872 23072 44878
rect 23020 44814 23072 44820
rect 23112 44804 23164 44810
rect 23112 44746 23164 44752
rect 23124 44538 23152 44746
rect 23112 44532 23164 44538
rect 23112 44474 23164 44480
rect 21824 44396 21876 44402
rect 21824 44338 21876 44344
rect 23848 44396 23900 44402
rect 23848 44338 23900 44344
rect 21548 43784 21600 43790
rect 21548 43726 21600 43732
rect 21560 43654 21588 43726
rect 21548 43648 21600 43654
rect 21548 43590 21600 43596
rect 21560 42702 21588 43590
rect 21836 43314 21864 44338
rect 23860 43994 23888 44338
rect 23848 43988 23900 43994
rect 23848 43930 23900 43936
rect 23204 43716 23256 43722
rect 23204 43658 23256 43664
rect 23216 43450 23244 43658
rect 23204 43444 23256 43450
rect 23204 43386 23256 43392
rect 22652 43376 22704 43382
rect 22652 43318 22704 43324
rect 21824 43308 21876 43314
rect 21824 43250 21876 43256
rect 21548 42696 21600 42702
rect 21548 42638 21600 42644
rect 22008 42696 22060 42702
rect 22008 42638 22060 42644
rect 21272 42628 21324 42634
rect 21272 42570 21324 42576
rect 21284 42362 21312 42570
rect 21272 42356 21324 42362
rect 21272 42298 21324 42304
rect 21548 42220 21600 42226
rect 21548 42162 21600 42168
rect 21560 41818 21588 42162
rect 21548 41812 21600 41818
rect 21548 41754 21600 41760
rect 22020 41682 22048 42638
rect 22664 42634 22692 43318
rect 23664 43308 23716 43314
rect 23664 43250 23716 43256
rect 23676 42906 23704 43250
rect 23664 42900 23716 42906
rect 23664 42842 23716 42848
rect 22652 42628 22704 42634
rect 22652 42570 22704 42576
rect 22664 42226 22692 42570
rect 24964 42362 24992 45834
rect 25044 45552 25096 45558
rect 25044 45494 25096 45500
rect 25056 44402 25084 45494
rect 25780 45484 25832 45490
rect 25780 45426 25832 45432
rect 25688 45280 25740 45286
rect 25688 45222 25740 45228
rect 25044 44396 25096 44402
rect 25044 44338 25096 44344
rect 25056 43858 25084 44338
rect 25044 43852 25096 43858
rect 25044 43794 25096 43800
rect 25596 43852 25648 43858
rect 25596 43794 25648 43800
rect 25608 43450 25636 43794
rect 25596 43444 25648 43450
rect 25596 43386 25648 43392
rect 24952 42356 25004 42362
rect 24952 42298 25004 42304
rect 25700 42294 25728 45222
rect 25792 42566 25820 45426
rect 27712 45416 27764 45422
rect 27712 45358 27764 45364
rect 27724 44878 27752 45358
rect 27712 44872 27764 44878
rect 27712 44814 27764 44820
rect 27528 44804 27580 44810
rect 27528 44746 27580 44752
rect 27160 44736 27212 44742
rect 27160 44678 27212 44684
rect 27068 44396 27120 44402
rect 27068 44338 27120 44344
rect 26424 44192 26476 44198
rect 26424 44134 26476 44140
rect 26436 42702 26464 44134
rect 27080 43994 27108 44338
rect 27068 43988 27120 43994
rect 27068 43930 27120 43936
rect 27172 43790 27200 44678
rect 27540 43994 27568 44746
rect 27724 44334 27752 44814
rect 27712 44328 27764 44334
rect 27712 44270 27764 44276
rect 27528 43988 27580 43994
rect 27528 43930 27580 43936
rect 27160 43784 27212 43790
rect 27160 43726 27212 43732
rect 27724 43722 27752 44270
rect 27712 43716 27764 43722
rect 27712 43658 27764 43664
rect 27724 43382 27752 43658
rect 27344 43376 27396 43382
rect 27344 43318 27396 43324
rect 27712 43376 27764 43382
rect 27712 43318 27764 43324
rect 26424 42696 26476 42702
rect 26424 42638 26476 42644
rect 27356 42634 27384 43318
rect 27436 43104 27488 43110
rect 27436 43046 27488 43052
rect 27344 42628 27396 42634
rect 27344 42570 27396 42576
rect 25780 42560 25832 42566
rect 25780 42502 25832 42508
rect 25688 42288 25740 42294
rect 25688 42230 25740 42236
rect 22652 42220 22704 42226
rect 22652 42162 22704 42168
rect 26148 42220 26200 42226
rect 26148 42162 26200 42168
rect 22008 41676 22060 41682
rect 22008 41618 22060 41624
rect 21272 41540 21324 41546
rect 21272 41482 21324 41488
rect 21284 41274 21312 41482
rect 21272 41268 21324 41274
rect 21272 41210 21324 41216
rect 22664 41138 22692 42162
rect 25872 42016 25924 42022
rect 25872 41958 25924 41964
rect 24952 41608 25004 41614
rect 24952 41550 25004 41556
rect 23756 41540 23808 41546
rect 23756 41482 23808 41488
rect 23204 41472 23256 41478
rect 23204 41414 23256 41420
rect 21272 41132 21324 41138
rect 21272 41074 21324 41080
rect 22652 41132 22704 41138
rect 22652 41074 22704 41080
rect 21088 40384 21140 40390
rect 21088 40326 21140 40332
rect 20812 39636 20864 39642
rect 20812 39578 20864 39584
rect 20628 39296 20680 39302
rect 20628 39238 20680 39244
rect 20640 39030 20668 39238
rect 20628 39024 20680 39030
rect 20628 38966 20680 38972
rect 20824 38962 20852 39578
rect 20812 38956 20864 38962
rect 20812 38898 20864 38904
rect 19524 38752 19576 38758
rect 19524 38694 19576 38700
rect 20536 38752 20588 38758
rect 20536 38694 20588 38700
rect 19536 38350 19564 38694
rect 19524 38344 19576 38350
rect 19524 38286 19576 38292
rect 18512 38276 18564 38282
rect 18512 38218 18564 38224
rect 18052 38004 18104 38010
rect 18052 37946 18104 37952
rect 18524 37874 18552 38218
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 18512 37868 18564 37874
rect 18512 37810 18564 37816
rect 19892 37664 19944 37670
rect 19892 37606 19944 37612
rect 17960 37460 18012 37466
rect 17960 37402 18012 37408
rect 19904 37262 19932 37606
rect 16672 37256 16724 37262
rect 16672 37198 16724 37204
rect 16948 37256 17000 37262
rect 16948 37198 17000 37204
rect 19892 37256 19944 37262
rect 19892 37198 19944 37204
rect 15660 37120 15712 37126
rect 15660 37062 15712 37068
rect 15476 34944 15528 34950
rect 15476 34886 15528 34892
rect 15488 33998 15516 34886
rect 15476 33992 15528 33998
rect 15476 33934 15528 33940
rect 15476 33312 15528 33318
rect 15476 33254 15528 33260
rect 15488 31822 15516 33254
rect 15476 31816 15528 31822
rect 15476 31758 15528 31764
rect 15568 31748 15620 31754
rect 15568 31690 15620 31696
rect 15476 31680 15528 31686
rect 15476 31622 15528 31628
rect 15488 30734 15516 31622
rect 15580 30938 15608 31690
rect 15568 30932 15620 30938
rect 15568 30874 15620 30880
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 15672 30326 15700 37062
rect 16684 36786 16712 37198
rect 20260 37188 20312 37194
rect 20260 37130 20312 37136
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 20272 36922 20300 37130
rect 19432 36916 19484 36922
rect 19432 36858 19484 36864
rect 20260 36916 20312 36922
rect 20260 36858 20312 36864
rect 16672 36780 16724 36786
rect 16672 36722 16724 36728
rect 18052 36780 18104 36786
rect 18052 36722 18104 36728
rect 16684 36242 16712 36722
rect 18064 36378 18092 36722
rect 18052 36372 18104 36378
rect 18052 36314 18104 36320
rect 16672 36236 16724 36242
rect 16672 36178 16724 36184
rect 16684 35494 16712 36178
rect 17868 36168 17920 36174
rect 17868 36110 17920 36116
rect 17776 36100 17828 36106
rect 17776 36042 17828 36048
rect 16672 35488 16724 35494
rect 16672 35430 16724 35436
rect 16684 35290 16712 35430
rect 17788 35290 17816 36042
rect 17880 35494 17908 36110
rect 17868 35488 17920 35494
rect 17868 35430 17920 35436
rect 19248 35488 19300 35494
rect 19248 35430 19300 35436
rect 19444 35442 19472 36858
rect 20548 36666 20576 38694
rect 21100 38350 21128 40326
rect 21284 40186 21312 41074
rect 22664 40610 22692 41074
rect 22572 40582 22692 40610
rect 22572 40526 22600 40582
rect 22560 40520 22612 40526
rect 22560 40462 22612 40468
rect 21272 40180 21324 40186
rect 21272 40122 21324 40128
rect 22572 39982 22600 40462
rect 23216 40050 23244 41414
rect 23768 40730 23796 41482
rect 24964 41070 24992 41550
rect 25884 41206 25912 41958
rect 25872 41200 25924 41206
rect 25872 41142 25924 41148
rect 24952 41064 25004 41070
rect 24952 41006 25004 41012
rect 24584 40928 24636 40934
rect 24584 40870 24636 40876
rect 23756 40724 23808 40730
rect 23756 40666 23808 40672
rect 24596 40526 24624 40870
rect 24964 40594 24992 41006
rect 24952 40588 25004 40594
rect 24952 40530 25004 40536
rect 24584 40520 24636 40526
rect 24584 40462 24636 40468
rect 24964 40118 24992 40530
rect 26160 40186 26188 42162
rect 26608 41472 26660 41478
rect 26608 41414 26660 41420
rect 26424 40928 26476 40934
rect 26424 40870 26476 40876
rect 26148 40180 26200 40186
rect 26148 40122 26200 40128
rect 24952 40112 25004 40118
rect 24952 40054 25004 40060
rect 26436 40050 26464 40870
rect 26620 40526 26648 41414
rect 27160 41132 27212 41138
rect 27160 41074 27212 41080
rect 27172 40730 27200 41074
rect 27160 40724 27212 40730
rect 27160 40666 27212 40672
rect 26608 40520 26660 40526
rect 26608 40462 26660 40468
rect 23020 40044 23072 40050
rect 23020 39986 23072 39992
rect 23204 40044 23256 40050
rect 23204 39986 23256 39992
rect 26424 40044 26476 40050
rect 26424 39986 26476 39992
rect 22560 39976 22612 39982
rect 22560 39918 22612 39924
rect 22572 39438 22600 39918
rect 22560 39432 22612 39438
rect 22560 39374 22612 39380
rect 23032 39098 23060 39986
rect 24308 39840 24360 39846
rect 24308 39782 24360 39788
rect 24320 39438 24348 39782
rect 24308 39432 24360 39438
rect 24308 39374 24360 39380
rect 24400 39432 24452 39438
rect 24400 39374 24452 39380
rect 23848 39296 23900 39302
rect 23848 39238 23900 39244
rect 23020 39092 23072 39098
rect 23020 39034 23072 39040
rect 23860 39030 23888 39238
rect 23848 39024 23900 39030
rect 23848 38966 23900 38972
rect 24412 38962 24440 39374
rect 24400 38956 24452 38962
rect 24400 38898 24452 38904
rect 24412 38350 24440 38898
rect 21088 38344 21140 38350
rect 21088 38286 21140 38292
rect 21824 38344 21876 38350
rect 21824 38286 21876 38292
rect 24400 38344 24452 38350
rect 24400 38286 24452 38292
rect 26240 38344 26292 38350
rect 26240 38286 26292 38292
rect 20628 38208 20680 38214
rect 20628 38150 20680 38156
rect 20640 37942 20668 38150
rect 20628 37936 20680 37942
rect 20628 37878 20680 37884
rect 21836 37874 21864 38286
rect 22376 38276 22428 38282
rect 22376 38218 22428 38224
rect 22192 38208 22244 38214
rect 22192 38150 22244 38156
rect 21824 37868 21876 37874
rect 21824 37810 21876 37816
rect 22100 37664 22152 37670
rect 22100 37606 22152 37612
rect 21088 37256 21140 37262
rect 21088 37198 21140 37204
rect 20628 37120 20680 37126
rect 20628 37062 20680 37068
rect 20640 36854 20668 37062
rect 20628 36848 20680 36854
rect 20628 36790 20680 36796
rect 21100 36786 21128 37198
rect 21088 36780 21140 36786
rect 21088 36722 21140 36728
rect 20548 36638 20668 36666
rect 20536 36100 20588 36106
rect 20536 36042 20588 36048
rect 20168 36032 20220 36038
rect 20168 35974 20220 35980
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 16672 35284 16724 35290
rect 16672 35226 16724 35232
rect 17776 35284 17828 35290
rect 17776 35226 17828 35232
rect 16684 34610 16712 35226
rect 19260 35154 19288 35430
rect 19444 35414 19564 35442
rect 19248 35148 19300 35154
rect 19248 35090 19300 35096
rect 19536 35086 19564 35414
rect 19524 35080 19576 35086
rect 19524 35022 19576 35028
rect 18236 35012 18288 35018
rect 18236 34954 18288 34960
rect 18248 34746 18276 34954
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 18236 34740 18288 34746
rect 18236 34682 18288 34688
rect 16672 34604 16724 34610
rect 16672 34546 16724 34552
rect 18512 34604 18564 34610
rect 18512 34546 18564 34552
rect 16684 34066 16712 34546
rect 18524 34202 18552 34546
rect 19248 34536 19300 34542
rect 19248 34478 19300 34484
rect 18512 34196 18564 34202
rect 18512 34138 18564 34144
rect 16672 34060 16724 34066
rect 16672 34002 16724 34008
rect 16684 32978 16712 34002
rect 19260 33998 19288 34478
rect 19248 33992 19300 33998
rect 19248 33934 19300 33940
rect 18420 33924 18472 33930
rect 18420 33866 18472 33872
rect 18432 33658 18460 33866
rect 18420 33652 18472 33658
rect 18420 33594 18472 33600
rect 19260 33590 19288 33934
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19248 33584 19300 33590
rect 19248 33526 19300 33532
rect 18880 33516 18932 33522
rect 18880 33458 18932 33464
rect 16672 32972 16724 32978
rect 16672 32914 16724 32920
rect 16580 32836 16632 32842
rect 16580 32778 16632 32784
rect 16212 32768 16264 32774
rect 16212 32710 16264 32716
rect 16224 30734 16252 32710
rect 16592 32026 16620 32778
rect 16684 32434 16712 32914
rect 17960 32836 18012 32842
rect 17960 32778 18012 32784
rect 16672 32428 16724 32434
rect 16672 32370 16724 32376
rect 17316 32428 17368 32434
rect 17316 32370 17368 32376
rect 16580 32020 16632 32026
rect 16580 31962 16632 31968
rect 16684 31822 16712 32370
rect 16672 31816 16724 31822
rect 16672 31758 16724 31764
rect 16684 31346 16712 31758
rect 16672 31340 16724 31346
rect 16672 31282 16724 31288
rect 17328 30938 17356 32370
rect 17972 32298 18000 32778
rect 18052 32768 18104 32774
rect 18052 32710 18104 32716
rect 18064 32502 18092 32710
rect 18892 32570 18920 33458
rect 19260 33454 19288 33526
rect 19248 33448 19300 33454
rect 19248 33390 19300 33396
rect 19260 32910 19288 33390
rect 20180 32910 20208 35974
rect 20548 33386 20576 36042
rect 20640 35894 20668 36638
rect 21100 36242 21128 36722
rect 21088 36236 21140 36242
rect 21088 36178 21140 36184
rect 20640 35866 20760 35894
rect 20732 35698 20760 35866
rect 22112 35766 22140 37606
rect 22204 36174 22232 38150
rect 22388 37466 22416 38218
rect 24412 37942 24440 38286
rect 24400 37936 24452 37942
rect 24400 37878 24452 37884
rect 23204 37868 23256 37874
rect 23204 37810 23256 37816
rect 22376 37460 22428 37466
rect 22376 37402 22428 37408
rect 23216 36922 23244 37810
rect 24412 37262 24440 37878
rect 24952 37868 25004 37874
rect 24952 37810 25004 37816
rect 24400 37256 24452 37262
rect 24400 37198 24452 37204
rect 24964 36922 24992 37810
rect 26252 37806 26280 38286
rect 26332 38208 26384 38214
rect 26332 38150 26384 38156
rect 26240 37800 26292 37806
rect 26240 37742 26292 37748
rect 25044 37664 25096 37670
rect 25044 37606 25096 37612
rect 25056 37262 25084 37606
rect 25044 37256 25096 37262
rect 25044 37198 25096 37204
rect 26252 37126 26280 37742
rect 26344 37262 26372 38150
rect 26332 37256 26384 37262
rect 26332 37198 26384 37204
rect 25780 37120 25832 37126
rect 25780 37062 25832 37068
rect 26240 37120 26292 37126
rect 26240 37062 26292 37068
rect 23204 36916 23256 36922
rect 23204 36858 23256 36864
rect 24952 36916 25004 36922
rect 24952 36858 25004 36864
rect 22468 36780 22520 36786
rect 22468 36722 22520 36728
rect 25044 36780 25096 36786
rect 25044 36722 25096 36728
rect 22480 36378 22508 36722
rect 23664 36712 23716 36718
rect 23664 36654 23716 36660
rect 22468 36372 22520 36378
rect 22468 36314 22520 36320
rect 22192 36168 22244 36174
rect 22192 36110 22244 36116
rect 23676 35834 23704 36654
rect 24400 36168 24452 36174
rect 24400 36110 24452 36116
rect 24412 35834 24440 36110
rect 25056 35834 25084 36722
rect 25792 36174 25820 37062
rect 26252 36174 26280 37062
rect 27356 36854 27384 42570
rect 27448 41614 27476 43046
rect 27724 42566 27752 43318
rect 27712 42560 27764 42566
rect 27712 42502 27764 42508
rect 27724 42158 27752 42502
rect 27712 42152 27764 42158
rect 27712 42094 27764 42100
rect 27724 41614 27752 42094
rect 27436 41608 27488 41614
rect 27436 41550 27488 41556
rect 27712 41608 27764 41614
rect 27712 41550 27764 41556
rect 27724 41070 27752 41550
rect 27712 41064 27764 41070
rect 27712 41006 27764 41012
rect 27724 40526 27752 41006
rect 27712 40520 27764 40526
rect 27712 40462 27764 40468
rect 27724 40050 27752 40462
rect 27712 40044 27764 40050
rect 27712 39986 27764 39992
rect 27528 39364 27580 39370
rect 27528 39306 27580 39312
rect 27540 38554 27568 39306
rect 27620 39296 27672 39302
rect 27620 39238 27672 39244
rect 27528 38548 27580 38554
rect 27528 38490 27580 38496
rect 27632 37942 27660 39238
rect 27724 39030 27752 39986
rect 28460 39098 28488 59978
rect 29368 59968 29420 59974
rect 29368 59910 29420 59916
rect 28540 59628 28592 59634
rect 28540 59570 28592 59576
rect 28552 55962 28580 59570
rect 29380 59022 29408 59910
rect 29932 59634 29960 60046
rect 31576 60036 31628 60042
rect 31576 59978 31628 59984
rect 31588 59770 31616 59978
rect 31576 59764 31628 59770
rect 31576 59706 31628 59712
rect 29920 59628 29972 59634
rect 29920 59570 29972 59576
rect 30288 59628 30340 59634
rect 30288 59570 30340 59576
rect 31760 59628 31812 59634
rect 31760 59570 31812 59576
rect 30300 59022 30328 59570
rect 29368 59016 29420 59022
rect 29368 58958 29420 58964
rect 30288 59016 30340 59022
rect 30288 58958 30340 58964
rect 29000 58880 29052 58886
rect 29000 58822 29052 58828
rect 29012 58614 29040 58822
rect 29000 58608 29052 58614
rect 29000 58550 29052 58556
rect 30300 58546 30328 58958
rect 31668 58880 31720 58886
rect 31668 58822 31720 58828
rect 31680 58614 31708 58822
rect 31772 58682 31800 59570
rect 32140 59566 32168 60046
rect 34072 59702 34100 60046
rect 36728 59968 36780 59974
rect 36728 59910 36780 59916
rect 34060 59696 34112 59702
rect 34060 59638 34112 59644
rect 35440 59628 35492 59634
rect 35440 59570 35492 59576
rect 32128 59560 32180 59566
rect 32128 59502 32180 59508
rect 34428 59560 34480 59566
rect 34480 59508 34560 59514
rect 34428 59502 34560 59508
rect 34440 59486 34560 59502
rect 32864 59424 32916 59430
rect 32864 59366 32916 59372
rect 32876 59022 32904 59366
rect 34532 59022 34560 59486
rect 34612 59424 34664 59430
rect 34612 59366 34664 59372
rect 32864 59016 32916 59022
rect 32864 58958 32916 58964
rect 34520 59016 34572 59022
rect 34520 58958 34572 58964
rect 31852 58948 31904 58954
rect 31852 58890 31904 58896
rect 31760 58676 31812 58682
rect 31760 58618 31812 58624
rect 31668 58608 31720 58614
rect 31668 58550 31720 58556
rect 30288 58540 30340 58546
rect 30288 58482 30340 58488
rect 29276 58336 29328 58342
rect 29276 58278 29328 58284
rect 29288 57934 29316 58278
rect 30300 57934 30328 58482
rect 29276 57928 29328 57934
rect 29276 57870 29328 57876
rect 30288 57928 30340 57934
rect 30288 57870 30340 57876
rect 28908 57860 28960 57866
rect 28908 57802 28960 57808
rect 28920 57050 28948 57802
rect 29000 57792 29052 57798
rect 29000 57734 29052 57740
rect 29012 57526 29040 57734
rect 29000 57520 29052 57526
rect 29000 57462 29052 57468
rect 30300 57458 30328 57870
rect 31864 57594 31892 58890
rect 32876 57934 32904 58958
rect 34624 57934 34652 59366
rect 34934 59324 35242 59344
rect 34934 59322 34940 59324
rect 34996 59322 35020 59324
rect 35076 59322 35100 59324
rect 35156 59322 35180 59324
rect 35236 59322 35242 59324
rect 34996 59270 34998 59322
rect 35178 59270 35180 59322
rect 34934 59268 34940 59270
rect 34996 59268 35020 59270
rect 35076 59268 35100 59270
rect 35156 59268 35180 59270
rect 35236 59268 35242 59270
rect 34934 59248 35242 59268
rect 35348 59016 35400 59022
rect 35348 58958 35400 58964
rect 35360 58342 35388 58958
rect 35348 58336 35400 58342
rect 35348 58278 35400 58284
rect 34934 58236 35242 58256
rect 34934 58234 34940 58236
rect 34996 58234 35020 58236
rect 35076 58234 35100 58236
rect 35156 58234 35180 58236
rect 35236 58234 35242 58236
rect 34996 58182 34998 58234
rect 35178 58182 35180 58234
rect 34934 58180 34940 58182
rect 34996 58180 35020 58182
rect 35076 58180 35100 58182
rect 35156 58180 35180 58182
rect 35236 58180 35242 58182
rect 34934 58160 35242 58180
rect 35360 57934 35388 58278
rect 32864 57928 32916 57934
rect 32864 57870 32916 57876
rect 34612 57928 34664 57934
rect 34612 57870 34664 57876
rect 34704 57928 34756 57934
rect 34704 57870 34756 57876
rect 35348 57928 35400 57934
rect 35348 57870 35400 57876
rect 32220 57860 32272 57866
rect 32220 57802 32272 57808
rect 31852 57588 31904 57594
rect 31852 57530 31904 57536
rect 30288 57452 30340 57458
rect 30288 57394 30340 57400
rect 29000 57248 29052 57254
rect 29000 57190 29052 57196
rect 31208 57248 31260 57254
rect 31208 57190 31260 57196
rect 28908 57044 28960 57050
rect 28908 56986 28960 56992
rect 29012 56846 29040 57190
rect 31220 56846 31248 57190
rect 32232 57050 32260 57802
rect 32312 57792 32364 57798
rect 32312 57734 32364 57740
rect 32324 57526 32352 57734
rect 32312 57520 32364 57526
rect 32312 57462 32364 57468
rect 32772 57384 32824 57390
rect 32772 57326 32824 57332
rect 32220 57044 32272 57050
rect 32220 56986 32272 56992
rect 32784 56914 32812 57326
rect 32772 56908 32824 56914
rect 32772 56850 32824 56856
rect 29000 56840 29052 56846
rect 29000 56782 29052 56788
rect 31208 56840 31260 56846
rect 31208 56782 31260 56788
rect 32784 56778 32812 56850
rect 32876 56846 32904 57870
rect 34152 57792 34204 57798
rect 34152 57734 34204 57740
rect 34164 57526 34192 57734
rect 34152 57520 34204 57526
rect 34152 57462 34204 57468
rect 34060 57452 34112 57458
rect 34060 57394 34112 57400
rect 34072 57050 34100 57394
rect 34716 57390 34744 57870
rect 35452 57798 35480 59570
rect 36740 59022 36768 59910
rect 37568 59634 37596 60046
rect 38752 60036 38804 60042
rect 38752 59978 38804 59984
rect 38764 59770 38792 59978
rect 38752 59764 38804 59770
rect 38752 59706 38804 59712
rect 37556 59628 37608 59634
rect 37556 59570 37608 59576
rect 39028 59628 39080 59634
rect 39028 59570 39080 59576
rect 37568 59090 37596 59570
rect 39040 59226 39068 59570
rect 40420 59566 40448 60046
rect 41880 59628 41932 59634
rect 41880 59570 41932 59576
rect 40408 59560 40460 59566
rect 40408 59502 40460 59508
rect 39028 59220 39080 59226
rect 39028 59162 39080 59168
rect 37556 59084 37608 59090
rect 37556 59026 37608 59032
rect 36728 59016 36780 59022
rect 36728 58958 36780 58964
rect 37004 58880 37056 58886
rect 37004 58822 37056 58828
rect 37016 57934 37044 58822
rect 37568 58546 37596 59026
rect 38844 58948 38896 58954
rect 38844 58890 38896 58896
rect 38856 58682 38884 58890
rect 38844 58676 38896 58682
rect 38844 58618 38896 58624
rect 39028 58608 39080 58614
rect 39028 58550 39080 58556
rect 37280 58540 37332 58546
rect 37280 58482 37332 58488
rect 37556 58540 37608 58546
rect 37556 58482 37608 58488
rect 38568 58540 38620 58546
rect 38568 58482 38620 58488
rect 37292 57934 37320 58482
rect 38580 58138 38608 58482
rect 38568 58132 38620 58138
rect 38568 58074 38620 58080
rect 37004 57928 37056 57934
rect 37004 57870 37056 57876
rect 37280 57928 37332 57934
rect 37280 57870 37332 57876
rect 35440 57792 35492 57798
rect 35440 57734 35492 57740
rect 34704 57384 34756 57390
rect 34704 57326 34756 57332
rect 34060 57044 34112 57050
rect 34060 56986 34112 56992
rect 34716 56846 34744 57326
rect 36084 57248 36136 57254
rect 36084 57190 36136 57196
rect 34934 57148 35242 57168
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57072 35242 57092
rect 36096 56846 36124 57190
rect 37292 56914 37320 57870
rect 38660 57860 38712 57866
rect 38660 57802 38712 57808
rect 38672 57050 38700 57802
rect 39040 57526 39068 58550
rect 40420 58478 40448 59502
rect 40684 59424 40736 59430
rect 40684 59366 40736 59372
rect 40408 58472 40460 58478
rect 40408 58414 40460 58420
rect 40420 58002 40448 58414
rect 40408 57996 40460 58002
rect 40408 57938 40460 57944
rect 40420 57594 40448 57938
rect 40696 57934 40724 59366
rect 41892 58682 41920 59570
rect 43640 59566 43668 60046
rect 44180 59968 44232 59974
rect 44180 59910 44232 59916
rect 43628 59560 43680 59566
rect 43628 59502 43680 59508
rect 43352 59424 43404 59430
rect 43352 59366 43404 59372
rect 42800 59016 42852 59022
rect 42800 58958 42852 58964
rect 42616 58880 42668 58886
rect 42616 58822 42668 58828
rect 41880 58676 41932 58682
rect 41880 58618 41932 58624
rect 42628 58614 42656 58822
rect 42616 58608 42668 58614
rect 42616 58550 42668 58556
rect 40684 57928 40736 57934
rect 40684 57870 40736 57876
rect 41144 57792 41196 57798
rect 41144 57734 41196 57740
rect 40408 57588 40460 57594
rect 40408 57530 40460 57536
rect 39028 57520 39080 57526
rect 39028 57462 39080 57468
rect 38660 57044 38712 57050
rect 38660 56986 38712 56992
rect 40420 56914 40448 57530
rect 37280 56908 37332 56914
rect 37280 56850 37332 56856
rect 40408 56908 40460 56914
rect 40408 56850 40460 56856
rect 32864 56840 32916 56846
rect 32864 56782 32916 56788
rect 34704 56840 34756 56846
rect 34704 56782 34756 56788
rect 36084 56840 36136 56846
rect 36084 56782 36136 56788
rect 32772 56772 32824 56778
rect 32772 56714 32824 56720
rect 29184 56160 29236 56166
rect 29184 56102 29236 56108
rect 30380 56160 30432 56166
rect 30380 56102 30432 56108
rect 28540 55956 28592 55962
rect 28540 55898 28592 55904
rect 29196 55214 29224 56102
rect 29828 55412 29880 55418
rect 29828 55354 29880 55360
rect 29276 55276 29328 55282
rect 29276 55218 29328 55224
rect 29184 55208 29236 55214
rect 29184 55150 29236 55156
rect 29288 54602 29316 55218
rect 29460 55072 29512 55078
rect 29460 55014 29512 55020
rect 29472 54670 29500 55014
rect 29460 54664 29512 54670
rect 29460 54606 29512 54612
rect 29276 54596 29328 54602
rect 29276 54538 29328 54544
rect 29472 53106 29500 54606
rect 29552 54188 29604 54194
rect 29552 54130 29604 54136
rect 29564 53582 29592 54130
rect 29840 53582 29868 55354
rect 30196 55276 30248 55282
rect 30196 55218 30248 55224
rect 30208 54330 30236 55218
rect 30196 54324 30248 54330
rect 30196 54266 30248 54272
rect 29552 53576 29604 53582
rect 29552 53518 29604 53524
rect 29828 53576 29880 53582
rect 29828 53518 29880 53524
rect 30392 53242 30420 56102
rect 32784 55758 32812 56714
rect 32876 56370 32904 56782
rect 34244 56772 34296 56778
rect 34244 56714 34296 56720
rect 34256 56506 34284 56714
rect 34244 56500 34296 56506
rect 34244 56442 34296 56448
rect 32864 56364 32916 56370
rect 32864 56306 32916 56312
rect 34716 56302 34744 56782
rect 36084 56704 36136 56710
rect 36084 56646 36136 56652
rect 36096 56438 36124 56646
rect 36084 56432 36136 56438
rect 36084 56374 36136 56380
rect 37292 56370 37320 56850
rect 39028 56772 39080 56778
rect 39028 56714 39080 56720
rect 39040 56506 39068 56714
rect 39028 56500 39080 56506
rect 39028 56442 39080 56448
rect 40420 56370 40448 56850
rect 41156 56846 41184 57734
rect 42812 57526 42840 58958
rect 43168 58948 43220 58954
rect 43168 58890 43220 58896
rect 43180 57798 43208 58890
rect 43364 57934 43392 59366
rect 43640 58546 43668 59502
rect 44192 58614 44220 59910
rect 45572 59634 45600 60046
rect 46940 60036 46992 60042
rect 46940 59978 46992 59984
rect 46952 59770 46980 59978
rect 48780 59968 48832 59974
rect 48780 59910 48832 59916
rect 46940 59764 46992 59770
rect 46940 59706 46992 59712
rect 44456 59628 44508 59634
rect 44456 59570 44508 59576
rect 45560 59628 45612 59634
rect 45560 59570 45612 59576
rect 47032 59628 47084 59634
rect 47032 59570 47084 59576
rect 44468 59226 44496 59570
rect 44456 59220 44508 59226
rect 44456 59162 44508 59168
rect 45192 58948 45244 58954
rect 45192 58890 45244 58896
rect 45204 58682 45232 58890
rect 45192 58676 45244 58682
rect 45192 58618 45244 58624
rect 44180 58608 44232 58614
rect 44180 58550 44232 58556
rect 45572 58546 45600 59570
rect 47044 58682 47072 59570
rect 48504 59424 48556 59430
rect 48504 59366 48556 59372
rect 47308 58948 47360 58954
rect 47308 58890 47360 58896
rect 47032 58676 47084 58682
rect 47032 58618 47084 58624
rect 43628 58540 43680 58546
rect 43628 58482 43680 58488
rect 45560 58540 45612 58546
rect 45560 58482 45612 58488
rect 47124 58540 47176 58546
rect 47124 58482 47176 58488
rect 43352 57928 43404 57934
rect 43352 57870 43404 57876
rect 44272 57860 44324 57866
rect 44272 57802 44324 57808
rect 43168 57792 43220 57798
rect 43168 57734 43220 57740
rect 41788 57520 41840 57526
rect 41788 57462 41840 57468
rect 42800 57520 42852 57526
rect 42800 57462 42852 57468
rect 41144 56840 41196 56846
rect 41144 56782 41196 56788
rect 37280 56364 37332 56370
rect 37280 56306 37332 56312
rect 37648 56364 37700 56370
rect 37648 56306 37700 56312
rect 39028 56364 39080 56370
rect 39028 56306 39080 56312
rect 40408 56364 40460 56370
rect 40408 56306 40460 56312
rect 34704 56296 34756 56302
rect 34704 56238 34756 56244
rect 35348 56160 35400 56166
rect 35348 56102 35400 56108
rect 34934 56060 35242 56080
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55984 35242 56004
rect 35360 55758 35388 56102
rect 37660 55826 37688 56306
rect 39040 55962 39068 56306
rect 39028 55956 39080 55962
rect 39028 55898 39080 55904
rect 37648 55820 37700 55826
rect 37648 55762 37700 55768
rect 32128 55752 32180 55758
rect 32128 55694 32180 55700
rect 32772 55752 32824 55758
rect 32772 55694 32824 55700
rect 35348 55752 35400 55758
rect 35348 55694 35400 55700
rect 32140 55214 32168 55694
rect 33140 55684 33192 55690
rect 33140 55626 33192 55632
rect 32404 55412 32456 55418
rect 32404 55354 32456 55360
rect 32128 55208 32180 55214
rect 32128 55150 32180 55156
rect 30932 54528 30984 54534
rect 30932 54470 30984 54476
rect 30944 54262 30972 54470
rect 30932 54256 30984 54262
rect 30932 54198 30984 54204
rect 32140 54194 32168 55150
rect 32128 54188 32180 54194
rect 32128 54130 32180 54136
rect 32140 53582 32168 54130
rect 32128 53576 32180 53582
rect 32128 53518 32180 53524
rect 30840 53508 30892 53514
rect 30840 53450 30892 53456
rect 30852 53242 30880 53450
rect 30932 53440 30984 53446
rect 30932 53382 30984 53388
rect 30380 53236 30432 53242
rect 30380 53178 30432 53184
rect 30840 53236 30892 53242
rect 30840 53178 30892 53184
rect 30944 53174 30972 53382
rect 32416 53174 32444 55354
rect 32496 54596 32548 54602
rect 32496 54538 32548 54544
rect 30932 53168 30984 53174
rect 30932 53110 30984 53116
rect 32404 53168 32456 53174
rect 32404 53110 32456 53116
rect 29460 53100 29512 53106
rect 29460 53042 29512 53048
rect 28908 52012 28960 52018
rect 28908 51954 28960 51960
rect 29920 52012 29972 52018
rect 29920 51954 29972 51960
rect 28920 51270 28948 51954
rect 28908 51264 28960 51270
rect 28960 51224 29040 51252
rect 28908 51206 28960 51212
rect 28908 50924 28960 50930
rect 28908 50866 28960 50872
rect 28724 49768 28776 49774
rect 28920 49756 28948 50866
rect 29012 50318 29040 51224
rect 29092 50720 29144 50726
rect 29092 50662 29144 50668
rect 29000 50312 29052 50318
rect 29000 50254 29052 50260
rect 29104 49910 29132 50662
rect 29552 50312 29604 50318
rect 29552 50254 29604 50260
rect 29092 49904 29144 49910
rect 29092 49846 29144 49852
rect 29564 49842 29592 50254
rect 29932 49978 29960 51954
rect 30196 51808 30248 51814
rect 30196 51750 30248 51756
rect 30104 51400 30156 51406
rect 30104 51342 30156 51348
rect 30116 50998 30144 51342
rect 30104 50992 30156 50998
rect 30104 50934 30156 50940
rect 30116 50250 30144 50934
rect 30208 50318 30236 51750
rect 30472 51332 30524 51338
rect 30472 51274 30524 51280
rect 30288 51264 30340 51270
rect 30288 51206 30340 51212
rect 30196 50312 30248 50318
rect 30196 50254 30248 50260
rect 30104 50244 30156 50250
rect 30104 50186 30156 50192
rect 29920 49972 29972 49978
rect 29920 49914 29972 49920
rect 29552 49836 29604 49842
rect 29552 49778 29604 49784
rect 28776 49728 28948 49756
rect 28724 49710 28776 49716
rect 29564 49298 29592 49778
rect 29552 49292 29604 49298
rect 29552 49234 29604 49240
rect 30116 48686 30144 50186
rect 30300 49162 30328 51206
rect 30484 50522 30512 51274
rect 30472 50516 30524 50522
rect 30472 50458 30524 50464
rect 31300 50244 31352 50250
rect 31300 50186 31352 50192
rect 31312 49434 31340 50186
rect 32508 49910 32536 54538
rect 32772 54188 32824 54194
rect 32772 54130 32824 54136
rect 32784 53786 32812 54130
rect 32772 53780 32824 53786
rect 32772 53722 32824 53728
rect 33152 53242 33180 55626
rect 33508 55616 33560 55622
rect 33508 55558 33560 55564
rect 33416 55276 33468 55282
rect 33416 55218 33468 55224
rect 33428 54330 33456 55218
rect 33416 54324 33468 54330
rect 33416 54266 33468 54272
rect 33520 54194 33548 55558
rect 35360 55282 35388 55694
rect 36728 55684 36780 55690
rect 36728 55626 36780 55632
rect 36740 55418 36768 55626
rect 36728 55412 36780 55418
rect 36728 55354 36780 55360
rect 35348 55276 35400 55282
rect 35348 55218 35400 55224
rect 36636 55276 36688 55282
rect 36636 55218 36688 55224
rect 34934 54972 35242 54992
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54896 35242 54916
rect 36648 54874 36676 55218
rect 36636 54868 36688 54874
rect 36636 54810 36688 54816
rect 37660 54670 37688 55762
rect 40132 55752 40184 55758
rect 40132 55694 40184 55700
rect 38936 55412 38988 55418
rect 38936 55354 38988 55360
rect 37648 54664 37700 54670
rect 37648 54606 37700 54612
rect 33968 54596 34020 54602
rect 33968 54538 34020 54544
rect 33980 54262 34008 54538
rect 33968 54256 34020 54262
rect 33968 54198 34020 54204
rect 33508 54188 33560 54194
rect 33508 54130 33560 54136
rect 33980 54126 34008 54198
rect 33968 54120 34020 54126
rect 33968 54062 34020 54068
rect 33232 53984 33284 53990
rect 33232 53926 33284 53932
rect 33140 53236 33192 53242
rect 33140 53178 33192 53184
rect 33244 52494 33272 53926
rect 33980 53106 34008 54062
rect 38660 53984 38712 53990
rect 38660 53926 38712 53932
rect 34934 53884 35242 53904
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53808 35242 53828
rect 38672 53582 38700 53926
rect 34704 53576 34756 53582
rect 34704 53518 34756 53524
rect 37924 53576 37976 53582
rect 37924 53518 37976 53524
rect 38660 53576 38712 53582
rect 38660 53518 38712 53524
rect 34060 53508 34112 53514
rect 34060 53450 34112 53456
rect 33968 53100 34020 53106
rect 33968 53042 34020 53048
rect 34072 52698 34100 53450
rect 34716 53106 34744 53518
rect 36084 53440 36136 53446
rect 36084 53382 36136 53388
rect 36096 53174 36124 53382
rect 36084 53168 36136 53174
rect 36084 53110 36136 53116
rect 37936 53106 37964 53518
rect 38948 53174 38976 55354
rect 40144 55350 40172 55694
rect 41800 55690 41828 57462
rect 42812 56930 42840 57462
rect 44284 57458 44312 57802
rect 43812 57452 43864 57458
rect 43812 57394 43864 57400
rect 44272 57452 44324 57458
rect 44272 57394 44324 57400
rect 45652 57452 45704 57458
rect 45652 57394 45704 57400
rect 42720 56914 42932 56930
rect 42708 56908 42932 56914
rect 42760 56902 42932 56908
rect 42708 56850 42760 56856
rect 42800 56772 42852 56778
rect 42800 56714 42852 56720
rect 42248 56704 42300 56710
rect 42248 56646 42300 56652
rect 42340 56704 42392 56710
rect 42340 56646 42392 56652
rect 42260 56438 42288 56646
rect 42248 56432 42300 56438
rect 42248 56374 42300 56380
rect 41880 56364 41932 56370
rect 41880 56306 41932 56312
rect 41788 55684 41840 55690
rect 41788 55626 41840 55632
rect 41420 55616 41472 55622
rect 41420 55558 41472 55564
rect 41432 55350 41460 55558
rect 40132 55344 40184 55350
rect 40132 55286 40184 55292
rect 40500 55344 40552 55350
rect 40500 55286 40552 55292
rect 41420 55344 41472 55350
rect 41420 55286 41472 55292
rect 40512 55214 40540 55286
rect 41328 55276 41380 55282
rect 41328 55218 41380 55224
rect 40500 55208 40552 55214
rect 40500 55150 40552 55156
rect 40512 54618 40540 55150
rect 41340 54874 41368 55218
rect 41800 55214 41828 55626
rect 41892 55418 41920 56306
rect 42352 55758 42380 56646
rect 42812 56506 42840 56714
rect 42800 56500 42852 56506
rect 42800 56442 42852 56448
rect 42904 56250 42932 56902
rect 43824 56506 43852 57394
rect 44284 56914 44312 57394
rect 44548 57248 44600 57254
rect 44548 57190 44600 57196
rect 45560 57248 45612 57254
rect 45560 57190 45612 57196
rect 44272 56908 44324 56914
rect 44272 56850 44324 56856
rect 43812 56500 43864 56506
rect 43812 56442 43864 56448
rect 44560 56438 44588 57190
rect 45008 56908 45060 56914
rect 45008 56850 45060 56856
rect 44548 56432 44600 56438
rect 44548 56374 44600 56380
rect 42812 56222 42932 56250
rect 42812 56166 42840 56222
rect 42800 56160 42852 56166
rect 42800 56102 42852 56108
rect 42812 55962 42840 56102
rect 42800 55956 42852 55962
rect 42800 55898 42852 55904
rect 43076 55956 43128 55962
rect 43076 55898 43128 55904
rect 42340 55752 42392 55758
rect 42340 55694 42392 55700
rect 41880 55412 41932 55418
rect 41880 55354 41932 55360
rect 41708 55186 41828 55214
rect 41328 54868 41380 54874
rect 41328 54810 41380 54816
rect 40592 54664 40644 54670
rect 40512 54612 40592 54618
rect 40512 54606 40644 54612
rect 39304 54596 39356 54602
rect 39304 54538 39356 54544
rect 40512 54590 40632 54606
rect 39316 53786 39344 54538
rect 40512 54262 40540 54590
rect 40500 54256 40552 54262
rect 40500 54198 40552 54204
rect 40040 54188 40092 54194
rect 40040 54130 40092 54136
rect 39304 53780 39356 53786
rect 39304 53722 39356 53728
rect 40052 53242 40080 54130
rect 40512 54126 40540 54198
rect 40500 54120 40552 54126
rect 40500 54062 40552 54068
rect 40512 53582 40540 54062
rect 41420 53984 41472 53990
rect 41420 53926 41472 53932
rect 40500 53576 40552 53582
rect 40500 53518 40552 53524
rect 40040 53236 40092 53242
rect 40040 53178 40092 53184
rect 38936 53168 38988 53174
rect 38936 53110 38988 53116
rect 40512 53106 40540 53518
rect 34704 53100 34756 53106
rect 34704 53042 34756 53048
rect 37924 53100 37976 53106
rect 37924 53042 37976 53048
rect 40500 53100 40552 53106
rect 40500 53042 40552 53048
rect 34060 52692 34112 52698
rect 34060 52634 34112 52640
rect 33232 52488 33284 52494
rect 33232 52430 33284 52436
rect 33232 52352 33284 52358
rect 33232 52294 33284 52300
rect 33244 52018 33272 52294
rect 34716 52018 34744 53042
rect 35348 52896 35400 52902
rect 35348 52838 35400 52844
rect 34934 52796 35242 52816
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52720 35242 52740
rect 35360 52086 35388 52838
rect 41432 52494 41460 53926
rect 39856 52488 39908 52494
rect 39856 52430 39908 52436
rect 41420 52488 41472 52494
rect 41420 52430 41472 52436
rect 35348 52080 35400 52086
rect 35348 52022 35400 52028
rect 33232 52012 33284 52018
rect 33232 51954 33284 51960
rect 34704 52012 34756 52018
rect 34704 51954 34756 51960
rect 35992 52012 36044 52018
rect 35992 51954 36044 51960
rect 33048 51808 33100 51814
rect 33048 51750 33100 51756
rect 33060 51406 33088 51750
rect 33048 51400 33100 51406
rect 33048 51342 33100 51348
rect 33244 51338 33272 51954
rect 34934 51708 35242 51728
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51632 35242 51652
rect 33232 51332 33284 51338
rect 33232 51274 33284 51280
rect 34612 51332 34664 51338
rect 34612 51274 34664 51280
rect 33244 50930 33272 51274
rect 34152 51264 34204 51270
rect 34152 51206 34204 51212
rect 34164 50998 34192 51206
rect 34624 51066 34652 51274
rect 34612 51060 34664 51066
rect 34612 51002 34664 51008
rect 34152 50992 34204 50998
rect 34152 50934 34204 50940
rect 33232 50924 33284 50930
rect 33232 50866 33284 50872
rect 32772 50176 32824 50182
rect 32772 50118 32824 50124
rect 32496 49904 32548 49910
rect 32496 49846 32548 49852
rect 31300 49428 31352 49434
rect 31300 49370 31352 49376
rect 32784 49230 32812 50118
rect 33244 49978 33272 50866
rect 34934 50620 35242 50640
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50544 35242 50564
rect 34704 50312 34756 50318
rect 34704 50254 34756 50260
rect 33232 49972 33284 49978
rect 33232 49914 33284 49920
rect 34716 49842 34744 50254
rect 34796 49904 34848 49910
rect 34796 49846 34848 49852
rect 34704 49836 34756 49842
rect 34704 49778 34756 49784
rect 34808 49230 34836 49846
rect 36004 49774 36032 51954
rect 37188 51944 37240 51950
rect 37188 51886 37240 51892
rect 36636 51808 36688 51814
rect 36636 51750 36688 51756
rect 36544 51400 36596 51406
rect 36544 51342 36596 51348
rect 36084 51264 36136 51270
rect 36084 51206 36136 51212
rect 36096 50998 36124 51206
rect 36084 50992 36136 50998
rect 36084 50934 36136 50940
rect 36556 50930 36584 51342
rect 36544 50924 36596 50930
rect 36544 50866 36596 50872
rect 36452 50720 36504 50726
rect 36452 50662 36504 50668
rect 36464 50318 36492 50662
rect 36556 50386 36584 50866
rect 36544 50380 36596 50386
rect 36544 50322 36596 50328
rect 36452 50312 36504 50318
rect 36452 50254 36504 50260
rect 36084 50176 36136 50182
rect 36084 50118 36136 50124
rect 36096 49910 36124 50118
rect 36084 49904 36136 49910
rect 36084 49846 36136 49852
rect 36556 49842 36584 50322
rect 36648 50318 36676 51750
rect 37200 51406 37228 51886
rect 39868 51474 39896 52430
rect 41708 52154 41736 55186
rect 41788 54596 41840 54602
rect 41788 54538 41840 54544
rect 41800 52698 41828 54538
rect 42616 54188 42668 54194
rect 42616 54130 42668 54136
rect 42628 53786 42656 54130
rect 42616 53780 42668 53786
rect 42616 53722 42668 53728
rect 43088 53650 43116 55898
rect 45020 55826 45048 56850
rect 45008 55820 45060 55826
rect 45008 55762 45060 55768
rect 45572 55758 45600 57190
rect 45664 56506 45692 57394
rect 46296 56772 46348 56778
rect 46296 56714 46348 56720
rect 45652 56500 45704 56506
rect 45652 56442 45704 56448
rect 46308 55962 46336 56714
rect 46388 56704 46440 56710
rect 46388 56646 46440 56652
rect 46296 55956 46348 55962
rect 46296 55898 46348 55904
rect 45560 55752 45612 55758
rect 45560 55694 45612 55700
rect 46400 55350 46428 56646
rect 46388 55344 46440 55350
rect 46388 55286 46440 55292
rect 45192 55276 45244 55282
rect 45192 55218 45244 55224
rect 45204 54754 45232 55218
rect 46480 55072 46532 55078
rect 46480 55014 46532 55020
rect 45204 54726 45324 54754
rect 45296 54670 45324 54726
rect 46492 54670 46520 55014
rect 45284 54664 45336 54670
rect 45284 54606 45336 54612
rect 46480 54664 46532 54670
rect 46480 54606 46532 54612
rect 44548 54596 44600 54602
rect 44548 54538 44600 54544
rect 44180 54528 44232 54534
rect 44180 54470 44232 54476
rect 43076 53644 43128 53650
rect 43076 53586 43128 53592
rect 41880 53508 41932 53514
rect 41880 53450 41932 53456
rect 41892 53242 41920 53450
rect 41880 53236 41932 53242
rect 41880 53178 41932 53184
rect 44192 53174 44220 54470
rect 44364 53508 44416 53514
rect 44364 53450 44416 53456
rect 44180 53168 44232 53174
rect 44180 53110 44232 53116
rect 43076 52896 43128 52902
rect 43076 52838 43128 52844
rect 41788 52692 41840 52698
rect 41788 52634 41840 52640
rect 43088 52562 43116 52838
rect 44376 52698 44404 53450
rect 44456 53440 44508 53446
rect 44456 53382 44508 53388
rect 44364 52692 44416 52698
rect 44364 52634 44416 52640
rect 43076 52556 43128 52562
rect 43076 52498 43128 52504
rect 40316 52148 40368 52154
rect 40316 52090 40368 52096
rect 41696 52148 41748 52154
rect 41696 52090 41748 52096
rect 43076 52148 43128 52154
rect 43076 52090 43128 52096
rect 39948 52012 40000 52018
rect 39948 51954 40000 51960
rect 39856 51468 39908 51474
rect 39856 51410 39908 51416
rect 37188 51400 37240 51406
rect 37188 51342 37240 51348
rect 37200 50930 37228 51342
rect 37832 51332 37884 51338
rect 37832 51274 37884 51280
rect 37188 50924 37240 50930
rect 37188 50866 37240 50872
rect 37844 50522 37872 51274
rect 37924 51264 37976 51270
rect 37924 51206 37976 51212
rect 37936 50998 37964 51206
rect 37924 50992 37976 50998
rect 37924 50934 37976 50940
rect 38752 50924 38804 50930
rect 38752 50866 38804 50872
rect 38660 50720 38712 50726
rect 38660 50662 38712 50668
rect 37832 50516 37884 50522
rect 37832 50458 37884 50464
rect 36636 50312 36688 50318
rect 36636 50254 36688 50260
rect 38672 49910 38700 50662
rect 38660 49904 38712 49910
rect 38660 49846 38712 49852
rect 36544 49836 36596 49842
rect 36544 49778 36596 49784
rect 37280 49836 37332 49842
rect 37280 49778 37332 49784
rect 35992 49768 36044 49774
rect 35992 49710 36044 49716
rect 34934 49532 35242 49552
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49456 35242 49476
rect 36556 49434 36584 49778
rect 36544 49428 36596 49434
rect 36544 49370 36596 49376
rect 31760 49224 31812 49230
rect 31760 49166 31812 49172
rect 32772 49224 32824 49230
rect 32772 49166 32824 49172
rect 34796 49224 34848 49230
rect 34796 49166 34848 49172
rect 30288 49156 30340 49162
rect 30288 49098 30340 49104
rect 31772 48686 31800 49166
rect 33140 49088 33192 49094
rect 33140 49030 33192 49036
rect 33152 48822 33180 49030
rect 33140 48816 33192 48822
rect 33140 48758 33192 48764
rect 34336 48816 34388 48822
rect 34336 48758 34388 48764
rect 32956 48748 33008 48754
rect 32956 48690 33008 48696
rect 30104 48680 30156 48686
rect 30104 48622 30156 48628
rect 31760 48680 31812 48686
rect 31760 48622 31812 48628
rect 30116 48142 30144 48622
rect 31576 48544 31628 48550
rect 31576 48486 31628 48492
rect 31588 48142 31616 48486
rect 32968 48346 32996 48690
rect 33508 48544 33560 48550
rect 33508 48486 33560 48492
rect 34244 48544 34296 48550
rect 34244 48486 34296 48492
rect 32956 48340 33008 48346
rect 32956 48282 33008 48288
rect 33520 48142 33548 48486
rect 30104 48136 30156 48142
rect 30104 48078 30156 48084
rect 31576 48136 31628 48142
rect 31576 48078 31628 48084
rect 32220 48136 32272 48142
rect 32220 48078 32272 48084
rect 33508 48136 33560 48142
rect 33508 48078 33560 48084
rect 29000 47728 29052 47734
rect 29000 47670 29052 47676
rect 29012 46170 29040 47670
rect 30012 47456 30064 47462
rect 30012 47398 30064 47404
rect 29184 47184 29236 47190
rect 29184 47126 29236 47132
rect 29092 46572 29144 46578
rect 29092 46514 29144 46520
rect 29000 46164 29052 46170
rect 29000 46106 29052 46112
rect 29104 45082 29132 46514
rect 29092 45076 29144 45082
rect 29092 45018 29144 45024
rect 29196 43790 29224 47126
rect 30024 47054 30052 47398
rect 30116 47054 30144 48078
rect 31760 48000 31812 48006
rect 31760 47942 31812 47948
rect 31772 47734 31800 47942
rect 31760 47728 31812 47734
rect 31760 47670 31812 47676
rect 32232 47666 32260 48078
rect 32220 47660 32272 47666
rect 32220 47602 32272 47608
rect 33784 47456 33836 47462
rect 33784 47398 33836 47404
rect 33796 47054 33824 47398
rect 30012 47048 30064 47054
rect 30012 46990 30064 46996
rect 30104 47048 30156 47054
rect 30104 46990 30156 46996
rect 33784 47048 33836 47054
rect 33784 46990 33836 46996
rect 30116 46866 30144 46990
rect 30024 46838 30144 46866
rect 32496 46912 32548 46918
rect 32496 46854 32548 46860
rect 30024 46374 30052 46838
rect 32508 46646 32536 46854
rect 34256 46646 34284 48486
rect 34348 48142 34376 48758
rect 35624 48748 35676 48754
rect 35624 48690 35676 48696
rect 34934 48444 35242 48464
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48368 35242 48388
rect 34336 48136 34388 48142
rect 34336 48078 34388 48084
rect 34348 47666 34376 48078
rect 35636 47802 35664 48690
rect 36556 48210 36584 49370
rect 37292 48754 37320 49778
rect 38764 49774 38792 50866
rect 39868 50726 39896 51410
rect 39960 51066 39988 51954
rect 40132 51808 40184 51814
rect 40132 51750 40184 51756
rect 39948 51060 40000 51066
rect 39948 51002 40000 51008
rect 39856 50720 39908 50726
rect 39856 50662 39908 50668
rect 39868 50386 39896 50662
rect 39856 50380 39908 50386
rect 39856 50322 39908 50328
rect 38752 49768 38804 49774
rect 38752 49710 38804 49716
rect 39868 49298 39896 50322
rect 40144 50318 40172 51750
rect 40132 50312 40184 50318
rect 40132 50254 40184 50260
rect 39856 49292 39908 49298
rect 39856 49234 39908 49240
rect 40328 49094 40356 52090
rect 40960 52012 41012 52018
rect 40960 51954 41012 51960
rect 40408 49700 40460 49706
rect 40408 49642 40460 49648
rect 40316 49088 40368 49094
rect 40316 49030 40368 49036
rect 37280 48748 37332 48754
rect 37280 48690 37332 48696
rect 38752 48748 38804 48754
rect 38752 48690 38804 48696
rect 38016 48544 38068 48550
rect 38016 48486 38068 48492
rect 36544 48204 36596 48210
rect 36544 48146 36596 48152
rect 35992 48068 36044 48074
rect 35992 48010 36044 48016
rect 35624 47796 35676 47802
rect 35624 47738 35676 47744
rect 34336 47660 34388 47666
rect 34336 47602 34388 47608
rect 34520 47660 34572 47666
rect 34520 47602 34572 47608
rect 34348 47546 34376 47602
rect 34348 47518 34468 47546
rect 34440 47054 34468 47518
rect 34428 47048 34480 47054
rect 34428 46990 34480 46996
rect 34440 46646 34468 46990
rect 32496 46640 32548 46646
rect 32496 46582 32548 46588
rect 34244 46640 34296 46646
rect 34244 46582 34296 46588
rect 34428 46640 34480 46646
rect 34428 46582 34480 46588
rect 30012 46368 30064 46374
rect 30012 46310 30064 46316
rect 30196 46368 30248 46374
rect 30196 46310 30248 46316
rect 33508 46368 33560 46374
rect 33508 46310 33560 46316
rect 30024 46034 30052 46310
rect 30012 46028 30064 46034
rect 30012 45970 30064 45976
rect 30208 45966 30236 46310
rect 33520 45966 33548 46310
rect 34440 46034 34468 46582
rect 34532 46170 34560 47602
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 36004 47258 36032 48010
rect 36556 47666 36584 48146
rect 37924 48000 37976 48006
rect 37924 47942 37976 47948
rect 36544 47660 36596 47666
rect 36544 47602 36596 47608
rect 37372 47660 37424 47666
rect 37372 47602 37424 47608
rect 35992 47252 36044 47258
rect 35992 47194 36044 47200
rect 35348 46980 35400 46986
rect 35348 46922 35400 46928
rect 35360 46714 35388 46922
rect 37280 46912 37332 46918
rect 37280 46854 37332 46860
rect 35348 46708 35400 46714
rect 35348 46650 35400 46656
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 34520 46164 34572 46170
rect 34520 46106 34572 46112
rect 34428 46028 34480 46034
rect 34428 45970 34480 45976
rect 37292 45966 37320 46854
rect 37384 46170 37412 47602
rect 37936 47054 37964 47942
rect 37924 47048 37976 47054
rect 37924 46990 37976 46996
rect 37464 46980 37516 46986
rect 37464 46922 37516 46928
rect 37476 46374 37504 46922
rect 37464 46368 37516 46374
rect 37464 46310 37516 46316
rect 37372 46164 37424 46170
rect 37372 46106 37424 46112
rect 37476 46034 37504 46310
rect 37464 46028 37516 46034
rect 37464 45970 37516 45976
rect 38028 45966 38056 48486
rect 38660 47456 38712 47462
rect 38660 47398 38712 47404
rect 38672 46646 38700 47398
rect 38660 46640 38712 46646
rect 38660 46582 38712 46588
rect 38764 46442 38792 48690
rect 40328 47734 40356 49030
rect 40420 48686 40448 49642
rect 40500 49632 40552 49638
rect 40500 49574 40552 49580
rect 40512 49230 40540 49574
rect 40500 49224 40552 49230
rect 40500 49166 40552 49172
rect 40408 48680 40460 48686
rect 40408 48622 40460 48628
rect 40420 48142 40448 48622
rect 40408 48136 40460 48142
rect 40408 48078 40460 48084
rect 40316 47728 40368 47734
rect 40316 47670 40368 47676
rect 40420 47054 40448 48078
rect 40408 47048 40460 47054
rect 40408 46990 40460 46996
rect 40132 46980 40184 46986
rect 40132 46922 40184 46928
rect 38752 46436 38804 46442
rect 38752 46378 38804 46384
rect 40144 46170 40172 46922
rect 40420 46578 40448 46990
rect 40408 46572 40460 46578
rect 40408 46514 40460 46520
rect 40684 46368 40736 46374
rect 40684 46310 40736 46316
rect 40132 46164 40184 46170
rect 40132 46106 40184 46112
rect 40696 45966 40724 46310
rect 30196 45960 30248 45966
rect 30196 45902 30248 45908
rect 33508 45960 33560 45966
rect 33508 45902 33560 45908
rect 37280 45960 37332 45966
rect 37280 45902 37332 45908
rect 38016 45960 38068 45966
rect 38016 45902 38068 45908
rect 40592 45960 40644 45966
rect 40592 45902 40644 45908
rect 40684 45960 40736 45966
rect 40684 45902 40736 45908
rect 31208 45892 31260 45898
rect 31208 45834 31260 45840
rect 30288 45824 30340 45830
rect 30288 45766 30340 45772
rect 30104 45484 30156 45490
rect 30104 45426 30156 45432
rect 29736 45280 29788 45286
rect 29736 45222 29788 45228
rect 29748 44878 29776 45222
rect 29736 44872 29788 44878
rect 29736 44814 29788 44820
rect 29736 44192 29788 44198
rect 29736 44134 29788 44140
rect 29184 43784 29236 43790
rect 29184 43726 29236 43732
rect 29748 43382 29776 44134
rect 30116 43450 30144 45426
rect 30300 44470 30328 45766
rect 30380 45280 30432 45286
rect 30380 45222 30432 45228
rect 30392 44878 30420 45222
rect 31220 45082 31248 45834
rect 40604 45558 40632 45902
rect 40592 45552 40644 45558
rect 40592 45494 40644 45500
rect 31484 45484 31536 45490
rect 31484 45426 31536 45432
rect 34796 45484 34848 45490
rect 34796 45426 34848 45432
rect 36544 45484 36596 45490
rect 36544 45426 36596 45432
rect 39212 45484 39264 45490
rect 39212 45426 39264 45432
rect 31208 45076 31260 45082
rect 31208 45018 31260 45024
rect 30380 44872 30432 44878
rect 30380 44814 30432 44820
rect 30392 44470 30420 44814
rect 31496 44538 31524 45426
rect 31668 45416 31720 45422
rect 31668 45358 31720 45364
rect 31576 45280 31628 45286
rect 31576 45222 31628 45228
rect 31484 44532 31536 44538
rect 31484 44474 31536 44480
rect 30288 44464 30340 44470
rect 30288 44406 30340 44412
rect 30380 44464 30432 44470
rect 30380 44406 30432 44412
rect 30392 43858 30420 44406
rect 30380 43852 30432 43858
rect 30380 43794 30432 43800
rect 30104 43444 30156 43450
rect 30104 43386 30156 43392
rect 29736 43376 29788 43382
rect 29736 43318 29788 43324
rect 28908 43308 28960 43314
rect 28908 43250 28960 43256
rect 28920 42362 28948 43250
rect 31588 42702 31616 45222
rect 31680 44878 31708 45358
rect 33784 45280 33836 45286
rect 33784 45222 33836 45228
rect 31668 44872 31720 44878
rect 31668 44814 31720 44820
rect 32036 44804 32088 44810
rect 32036 44746 32088 44752
rect 31944 44736 31996 44742
rect 31944 44678 31996 44684
rect 31956 43790 31984 44678
rect 31944 43784 31996 43790
rect 31944 43726 31996 43732
rect 31576 42696 31628 42702
rect 31576 42638 31628 42644
rect 32048 42566 32076 44746
rect 33796 44470 33824 45222
rect 34060 44804 34112 44810
rect 34060 44746 34112 44752
rect 33784 44464 33836 44470
rect 33784 44406 33836 44412
rect 32220 44396 32272 44402
rect 32220 44338 32272 44344
rect 32232 43994 32260 44338
rect 32772 44328 32824 44334
rect 32772 44270 32824 44276
rect 32220 43988 32272 43994
rect 32220 43930 32272 43936
rect 32784 43790 32812 44270
rect 33324 44192 33376 44198
rect 33324 44134 33376 44140
rect 33336 43790 33364 44134
rect 32772 43784 32824 43790
rect 32772 43726 32824 43732
rect 33324 43784 33376 43790
rect 33324 43726 33376 43732
rect 32784 43314 32812 43726
rect 32956 43716 33008 43722
rect 32956 43658 33008 43664
rect 32772 43308 32824 43314
rect 32772 43250 32824 43256
rect 32784 42702 32812 43250
rect 32772 42696 32824 42702
rect 32772 42638 32824 42644
rect 32128 42628 32180 42634
rect 32128 42570 32180 42576
rect 32036 42560 32088 42566
rect 32036 42502 32088 42508
rect 28908 42356 28960 42362
rect 28908 42298 28960 42304
rect 29000 42220 29052 42226
rect 29000 42162 29052 42168
rect 29012 41818 29040 42162
rect 29000 41812 29052 41818
rect 29000 41754 29052 41760
rect 32140 41614 32168 42570
rect 30196 41608 30248 41614
rect 30196 41550 30248 41556
rect 32128 41608 32180 41614
rect 32128 41550 32180 41556
rect 29644 41540 29696 41546
rect 29644 41482 29696 41488
rect 29656 41274 29684 41482
rect 29644 41268 29696 41274
rect 29644 41210 29696 41216
rect 29000 41132 29052 41138
rect 29000 41074 29052 41080
rect 29012 40730 29040 41074
rect 30208 41070 30236 41550
rect 31116 41540 31168 41546
rect 31116 41482 31168 41488
rect 30380 41472 30432 41478
rect 30380 41414 30432 41420
rect 30196 41064 30248 41070
rect 30196 41006 30248 41012
rect 30012 40928 30064 40934
rect 30012 40870 30064 40876
rect 29000 40724 29052 40730
rect 29000 40666 29052 40672
rect 29736 40452 29788 40458
rect 29736 40394 29788 40400
rect 29748 40186 29776 40394
rect 29736 40180 29788 40186
rect 29736 40122 29788 40128
rect 29644 39636 29696 39642
rect 29644 39578 29696 39584
rect 28448 39092 28500 39098
rect 28448 39034 28500 39040
rect 27712 39024 27764 39030
rect 27712 38966 27764 38972
rect 28540 38956 28592 38962
rect 28540 38898 28592 38904
rect 27712 38276 27764 38282
rect 27712 38218 27764 38224
rect 27620 37936 27672 37942
rect 27620 37878 27672 37884
rect 27724 37466 27752 38218
rect 27804 38208 27856 38214
rect 27804 38150 27856 38156
rect 27712 37460 27764 37466
rect 27712 37402 27764 37408
rect 27344 36848 27396 36854
rect 27344 36790 27396 36796
rect 27816 36378 27844 38150
rect 28552 38010 28580 38898
rect 28540 38004 28592 38010
rect 28540 37946 28592 37952
rect 27804 36372 27856 36378
rect 27804 36314 27856 36320
rect 25780 36168 25832 36174
rect 25780 36110 25832 36116
rect 26240 36168 26292 36174
rect 26240 36110 26292 36116
rect 27068 36168 27120 36174
rect 27068 36110 27120 36116
rect 23664 35828 23716 35834
rect 23664 35770 23716 35776
rect 24400 35828 24452 35834
rect 24400 35770 24452 35776
rect 25044 35828 25096 35834
rect 25044 35770 25096 35776
rect 22100 35760 22152 35766
rect 22100 35702 22152 35708
rect 23676 35698 23704 35770
rect 20720 35692 20772 35698
rect 20720 35634 20772 35640
rect 21088 35692 21140 35698
rect 21088 35634 21140 35640
rect 23664 35692 23716 35698
rect 23664 35634 23716 35640
rect 20628 34944 20680 34950
rect 20628 34886 20680 34892
rect 20640 34678 20668 34886
rect 20628 34672 20680 34678
rect 20628 34614 20680 34620
rect 20628 34400 20680 34406
rect 20628 34342 20680 34348
rect 20640 33998 20668 34342
rect 20628 33992 20680 33998
rect 20628 33934 20680 33940
rect 20732 33930 20760 35634
rect 21100 35154 21128 35634
rect 27080 35630 27108 36110
rect 28356 35692 28408 35698
rect 28356 35634 28408 35640
rect 27068 35624 27120 35630
rect 27068 35566 27120 35572
rect 27080 35494 27108 35566
rect 27068 35488 27120 35494
rect 27068 35430 27120 35436
rect 21088 35148 21140 35154
rect 21088 35090 21140 35096
rect 21100 34202 21128 35090
rect 27080 35086 27108 35430
rect 28368 35290 28396 35634
rect 28448 35488 28500 35494
rect 28448 35430 28500 35436
rect 28356 35284 28408 35290
rect 28356 35226 28408 35232
rect 24400 35080 24452 35086
rect 24400 35022 24452 35028
rect 26240 35080 26292 35086
rect 26240 35022 26292 35028
rect 27068 35080 27120 35086
rect 27068 35022 27120 35028
rect 22836 35012 22888 35018
rect 22836 34954 22888 34960
rect 22468 34944 22520 34950
rect 22468 34886 22520 34892
rect 21088 34196 21140 34202
rect 21088 34138 21140 34144
rect 21824 34196 21876 34202
rect 21824 34138 21876 34144
rect 20720 33924 20772 33930
rect 20720 33866 20772 33872
rect 20628 33856 20680 33862
rect 20628 33798 20680 33804
rect 20640 33590 20668 33798
rect 20628 33584 20680 33590
rect 20628 33526 20680 33532
rect 21836 33522 21864 34138
rect 21824 33516 21876 33522
rect 21824 33458 21876 33464
rect 22100 33516 22152 33522
rect 22100 33458 22152 33464
rect 20536 33380 20588 33386
rect 20536 33322 20588 33328
rect 19248 32904 19300 32910
rect 19248 32846 19300 32852
rect 20168 32904 20220 32910
rect 20168 32846 20220 32852
rect 18880 32564 18932 32570
rect 18880 32506 18932 32512
rect 18052 32496 18104 32502
rect 18052 32438 18104 32444
rect 19260 32434 19288 32846
rect 21836 32842 21864 33458
rect 22112 33114 22140 33458
rect 22100 33108 22152 33114
rect 22100 33050 22152 33056
rect 21824 32836 21876 32842
rect 21824 32778 21876 32784
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 21836 32434 21864 32778
rect 22480 32502 22508 34886
rect 22848 33114 22876 34954
rect 23756 34672 23808 34678
rect 23756 34614 23808 34620
rect 23768 34542 23796 34614
rect 23848 34604 23900 34610
rect 23848 34546 23900 34552
rect 23756 34536 23808 34542
rect 23756 34478 23808 34484
rect 23768 33522 23796 34478
rect 23756 33516 23808 33522
rect 23756 33458 23808 33464
rect 23204 33312 23256 33318
rect 23204 33254 23256 33260
rect 22836 33108 22888 33114
rect 22836 33050 22888 33056
rect 23216 32910 23244 33254
rect 23204 32904 23256 32910
rect 23204 32846 23256 32852
rect 23296 32836 23348 32842
rect 23296 32778 23348 32784
rect 22468 32496 22520 32502
rect 22468 32438 22520 32444
rect 19248 32428 19300 32434
rect 19248 32370 19300 32376
rect 21824 32428 21876 32434
rect 21824 32370 21876 32376
rect 17960 32292 18012 32298
rect 17960 32234 18012 32240
rect 19260 31890 19288 32370
rect 19248 31884 19300 31890
rect 19248 31826 19300 31832
rect 19260 31278 19288 31826
rect 21272 31816 21324 31822
rect 21272 31758 21324 31764
rect 22468 31816 22520 31822
rect 22468 31758 22520 31764
rect 20996 31680 21048 31686
rect 20996 31622 21048 31628
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19340 31340 19392 31346
rect 19340 31282 19392 31288
rect 19248 31272 19300 31278
rect 19248 31214 19300 31220
rect 17316 30932 17368 30938
rect 17316 30874 17368 30880
rect 15936 30728 15988 30734
rect 15936 30670 15988 30676
rect 16212 30728 16264 30734
rect 16212 30670 16264 30676
rect 15660 30320 15712 30326
rect 15660 30262 15712 30268
rect 15948 30190 15976 30670
rect 19352 30394 19380 31282
rect 19432 31136 19484 31142
rect 19432 31078 19484 31084
rect 19340 30388 19392 30394
rect 19340 30330 19392 30336
rect 15936 30184 15988 30190
rect 15936 30126 15988 30132
rect 18052 30184 18104 30190
rect 18052 30126 18104 30132
rect 15384 30116 15436 30122
rect 15384 30058 15436 30064
rect 15948 29646 15976 30126
rect 18064 30054 18092 30126
rect 18052 30048 18104 30054
rect 18052 29990 18104 29996
rect 19248 30048 19300 30054
rect 19248 29990 19300 29996
rect 14648 29640 14700 29646
rect 14648 29582 14700 29588
rect 15936 29640 15988 29646
rect 15936 29582 15988 29588
rect 17040 29640 17092 29646
rect 17040 29582 17092 29588
rect 14660 29170 14688 29582
rect 16120 29572 16172 29578
rect 16120 29514 16172 29520
rect 16028 29504 16080 29510
rect 16028 29446 16080 29452
rect 15476 29232 15528 29238
rect 15476 29174 15528 29180
rect 14096 29164 14148 29170
rect 14096 29106 14148 29112
rect 14648 29164 14700 29170
rect 14648 29106 14700 29112
rect 14108 28082 14136 29106
rect 14280 28960 14332 28966
rect 14280 28902 14332 28908
rect 14292 28150 14320 28902
rect 14280 28144 14332 28150
rect 14280 28086 14332 28092
rect 14096 28076 14148 28082
rect 14096 28018 14148 28024
rect 14096 27872 14148 27878
rect 14096 27814 14148 27820
rect 13544 27600 13596 27606
rect 13544 27542 13596 27548
rect 14108 27470 14136 27814
rect 14096 27464 14148 27470
rect 14096 27406 14148 27412
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 12256 27056 12308 27062
rect 12256 26998 12308 27004
rect 12532 27056 12584 27062
rect 12532 26998 12584 27004
rect 11796 26988 11848 26994
rect 11796 26930 11848 26936
rect 11808 26586 11836 26930
rect 11796 26580 11848 26586
rect 11796 26522 11848 26528
rect 12268 26382 12296 26998
rect 10324 26376 10376 26382
rect 10324 26318 10376 26324
rect 12072 26376 12124 26382
rect 12072 26318 12124 26324
rect 12256 26376 12308 26382
rect 12256 26318 12308 26324
rect 10336 25906 10364 26318
rect 5172 25900 5224 25906
rect 5172 25842 5224 25848
rect 6920 25900 6972 25906
rect 6920 25842 6972 25848
rect 9588 25900 9640 25906
rect 9588 25842 9640 25848
rect 10324 25900 10376 25906
rect 10324 25842 10376 25848
rect 4620 25696 4672 25702
rect 4620 25638 4672 25644
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4632 25378 4660 25638
rect 4540 25350 4660 25378
rect 4540 25294 4568 25350
rect 4528 25288 4580 25294
rect 4528 25230 4580 25236
rect 4344 25152 4396 25158
rect 4344 25094 4396 25100
rect 4356 24818 4384 25094
rect 4540 24886 4568 25230
rect 5184 24954 5212 25842
rect 12084 25838 12112 26318
rect 12544 26234 12572 26998
rect 13636 26988 13688 26994
rect 13636 26930 13688 26936
rect 13648 26382 13676 26930
rect 13636 26376 13688 26382
rect 13636 26318 13688 26324
rect 14096 26376 14148 26382
rect 14096 26318 14148 26324
rect 12452 26206 12572 26234
rect 8944 25832 8996 25838
rect 8944 25774 8996 25780
rect 12072 25832 12124 25838
rect 12072 25774 12124 25780
rect 5816 25696 5868 25702
rect 5816 25638 5868 25644
rect 5172 24948 5224 24954
rect 5172 24890 5224 24896
rect 4528 24880 4580 24886
rect 4528 24822 4580 24828
rect 4344 24812 4396 24818
rect 4344 24754 4396 24760
rect 1860 24744 1912 24750
rect 1860 24686 1912 24692
rect 1872 24274 1900 24686
rect 5828 24614 5856 25638
rect 6368 25288 6420 25294
rect 6368 25230 6420 25236
rect 6092 25220 6144 25226
rect 6092 25162 6144 25168
rect 3332 24608 3384 24614
rect 3332 24550 3384 24556
rect 5816 24608 5868 24614
rect 5816 24550 5868 24556
rect 1860 24268 1912 24274
rect 1860 24210 1912 24216
rect 3344 24206 3372 24550
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 3332 24200 3384 24206
rect 3332 24142 3384 24148
rect 5264 24132 5316 24138
rect 5264 24074 5316 24080
rect 3240 24064 3292 24070
rect 3240 24006 3292 24012
rect 3252 23798 3280 24006
rect 3240 23792 3292 23798
rect 3240 23734 3292 23740
rect 2228 23724 2280 23730
rect 2228 23666 2280 23672
rect 2240 23050 2268 23666
rect 3700 23520 3752 23526
rect 3700 23462 3752 23468
rect 5172 23520 5224 23526
rect 5172 23462 5224 23468
rect 3712 23118 3740 23462
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 5184 23186 5212 23462
rect 5172 23180 5224 23186
rect 5172 23122 5224 23128
rect 3700 23112 3752 23118
rect 3700 23054 3752 23060
rect 2228 23044 2280 23050
rect 2228 22986 2280 22992
rect 2240 22642 2268 22986
rect 3240 22976 3292 22982
rect 3240 22918 3292 22924
rect 3252 22710 3280 22918
rect 3240 22704 3292 22710
rect 3240 22646 3292 22652
rect 2228 22636 2280 22642
rect 2228 22578 2280 22584
rect 2240 21962 2268 22578
rect 3608 22432 3660 22438
rect 3608 22374 3660 22380
rect 3620 22030 3648 22374
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 5184 22030 5212 23122
rect 3608 22024 3660 22030
rect 3608 21966 3660 21972
rect 4436 22024 4488 22030
rect 4436 21966 4488 21972
rect 5172 22024 5224 22030
rect 5172 21966 5224 21972
rect 2228 21956 2280 21962
rect 2228 21898 2280 21904
rect 3424 21956 3476 21962
rect 3424 21898 3476 21904
rect 2136 21548 2188 21554
rect 2240 21536 2268 21898
rect 3240 21888 3292 21894
rect 3240 21830 3292 21836
rect 3252 21622 3280 21830
rect 3436 21690 3464 21898
rect 3424 21684 3476 21690
rect 3424 21626 3476 21632
rect 3240 21616 3292 21622
rect 3240 21558 3292 21564
rect 4448 21554 4476 21966
rect 5172 21888 5224 21894
rect 5172 21830 5224 21836
rect 5184 21622 5212 21830
rect 5172 21616 5224 21622
rect 5172 21558 5224 21564
rect 2188 21508 2268 21536
rect 4436 21548 4488 21554
rect 2136 21490 2188 21496
rect 4436 21490 4488 21496
rect 4896 21344 4948 21350
rect 4896 21286 4948 21292
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4344 21072 4396 21078
rect 4344 21014 4396 21020
rect 4356 20398 4384 21014
rect 4908 20466 4936 21286
rect 5276 20874 5304 24074
rect 6104 23866 6132 25162
rect 6380 24818 6408 25230
rect 8956 24886 8984 25774
rect 10324 25696 10376 25702
rect 10324 25638 10376 25644
rect 10336 25294 10364 25638
rect 10324 25288 10376 25294
rect 10324 25230 10376 25236
rect 12084 25226 12112 25774
rect 12072 25220 12124 25226
rect 12072 25162 12124 25168
rect 10324 25152 10376 25158
rect 10324 25094 10376 25100
rect 8944 24880 8996 24886
rect 8944 24822 8996 24828
rect 10336 24818 10364 25094
rect 12084 24818 12112 25162
rect 6368 24812 6420 24818
rect 6368 24754 6420 24760
rect 8024 24812 8076 24818
rect 8024 24754 8076 24760
rect 10324 24812 10376 24818
rect 10324 24754 10376 24760
rect 12072 24812 12124 24818
rect 12072 24754 12124 24760
rect 6184 24608 6236 24614
rect 6184 24550 6236 24556
rect 6092 23860 6144 23866
rect 6092 23802 6144 23808
rect 6196 23118 6224 24550
rect 6380 24410 6408 24754
rect 6368 24404 6420 24410
rect 6368 24346 6420 24352
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 6564 23322 6592 23666
rect 7012 23656 7064 23662
rect 7012 23598 7064 23604
rect 6552 23316 6604 23322
rect 6552 23258 6604 23264
rect 7024 23118 7052 23598
rect 8036 23322 8064 24754
rect 10416 24608 10468 24614
rect 10416 24550 10468 24556
rect 10428 24206 10456 24550
rect 12452 24410 12480 26206
rect 14108 25906 14136 26318
rect 14188 26308 14240 26314
rect 14188 26250 14240 26256
rect 13544 25900 13596 25906
rect 13544 25842 13596 25848
rect 14096 25900 14148 25906
rect 14096 25842 14148 25848
rect 13556 25498 13584 25842
rect 14200 25498 14228 26250
rect 13544 25492 13596 25498
rect 13544 25434 13596 25440
rect 14188 25492 14240 25498
rect 14188 25434 14240 25440
rect 14752 25362 14780 27406
rect 15108 26784 15160 26790
rect 15108 26726 15160 26732
rect 15120 26382 15148 26726
rect 15488 26518 15516 29174
rect 15476 26512 15528 26518
rect 15476 26454 15528 26460
rect 15108 26376 15160 26382
rect 15108 26318 15160 26324
rect 15936 26376 15988 26382
rect 15936 26318 15988 26324
rect 15948 25906 15976 26318
rect 16040 26314 16068 29446
rect 16132 29306 16160 29514
rect 16120 29300 16172 29306
rect 16120 29242 16172 29248
rect 16396 29164 16448 29170
rect 16396 29106 16448 29112
rect 16120 27872 16172 27878
rect 16120 27814 16172 27820
rect 16132 27470 16160 27814
rect 16408 27606 16436 29106
rect 17052 29102 17080 29582
rect 17316 29572 17368 29578
rect 17316 29514 17368 29520
rect 16672 29096 16724 29102
rect 16672 29038 16724 29044
rect 17040 29096 17092 29102
rect 17040 29038 17092 29044
rect 16684 28558 16712 29038
rect 16672 28552 16724 28558
rect 16672 28494 16724 28500
rect 16684 28014 16712 28494
rect 16856 28416 16908 28422
rect 16856 28358 16908 28364
rect 16868 28150 16896 28358
rect 16856 28144 16908 28150
rect 16856 28086 16908 28092
rect 16672 28008 16724 28014
rect 16672 27950 16724 27956
rect 16396 27600 16448 27606
rect 16396 27542 16448 27548
rect 16684 27470 16712 27950
rect 16120 27464 16172 27470
rect 16120 27406 16172 27412
rect 16672 27464 16724 27470
rect 16672 27406 16724 27412
rect 16684 26926 16712 27406
rect 16672 26920 16724 26926
rect 16672 26862 16724 26868
rect 16028 26308 16080 26314
rect 16028 26250 16080 26256
rect 15476 25900 15528 25906
rect 15476 25842 15528 25848
rect 15936 25900 15988 25906
rect 15936 25842 15988 25848
rect 15384 25696 15436 25702
rect 15384 25638 15436 25644
rect 14740 25356 14792 25362
rect 14740 25298 14792 25304
rect 13452 25220 13504 25226
rect 13452 25162 13504 25168
rect 13464 24954 13492 25162
rect 13452 24948 13504 24954
rect 13452 24890 13504 24896
rect 14752 24818 14780 25298
rect 15396 25294 15424 25638
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 14740 24812 14792 24818
rect 14740 24754 14792 24760
rect 13464 24410 13492 24754
rect 11520 24404 11572 24410
rect 11520 24346 11572 24352
rect 12440 24404 12492 24410
rect 12440 24346 12492 24352
rect 13452 24404 13504 24410
rect 13452 24346 13504 24352
rect 9220 24200 9272 24206
rect 9220 24142 9272 24148
rect 10416 24200 10468 24206
rect 10416 24142 10468 24148
rect 9232 23662 9260 24142
rect 11532 24070 11560 24346
rect 15488 24274 15516 25842
rect 16684 25294 16712 26862
rect 17328 26586 17356 29514
rect 17960 29504 18012 29510
rect 17960 29446 18012 29452
rect 17972 26994 18000 29446
rect 18064 28558 18092 29990
rect 19260 29714 19288 29990
rect 19248 29708 19300 29714
rect 19248 29650 19300 29656
rect 18696 29164 18748 29170
rect 18696 29106 18748 29112
rect 18708 28762 18736 29106
rect 18788 28960 18840 28966
rect 18788 28902 18840 28908
rect 18696 28756 18748 28762
rect 18696 28698 18748 28704
rect 18052 28552 18104 28558
rect 18052 28494 18104 28500
rect 18052 28416 18104 28422
rect 18052 28358 18104 28364
rect 18064 27130 18092 28358
rect 18800 28150 18828 28902
rect 19248 28552 19300 28558
rect 19248 28494 19300 28500
rect 18788 28144 18840 28150
rect 18788 28086 18840 28092
rect 19260 28082 19288 28494
rect 19444 28150 19472 31078
rect 20628 30728 20680 30734
rect 20628 30670 20680 30676
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19984 30252 20036 30258
rect 19984 30194 20036 30200
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19996 28762 20024 30194
rect 20640 29714 20668 30670
rect 20628 29708 20680 29714
rect 20628 29650 20680 29656
rect 20640 29578 20668 29650
rect 20628 29572 20680 29578
rect 20628 29514 20680 29520
rect 20640 29306 20668 29514
rect 20628 29300 20680 29306
rect 20628 29242 20680 29248
rect 20076 29164 20128 29170
rect 20076 29106 20128 29112
rect 19984 28756 20036 28762
rect 19984 28698 20036 28704
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19432 28144 19484 28150
rect 19432 28086 19484 28092
rect 19248 28076 19300 28082
rect 19248 28018 19300 28024
rect 18420 27872 18472 27878
rect 18420 27814 18472 27820
rect 18432 27470 18460 27814
rect 19260 27538 19288 28018
rect 19248 27532 19300 27538
rect 19248 27474 19300 27480
rect 18420 27464 18472 27470
rect 18420 27406 18472 27412
rect 18236 27328 18288 27334
rect 18236 27270 18288 27276
rect 18052 27124 18104 27130
rect 18052 27066 18104 27072
rect 18248 27062 18276 27270
rect 18236 27056 18288 27062
rect 18236 26998 18288 27004
rect 19260 26994 19288 27474
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 17960 26988 18012 26994
rect 17960 26930 18012 26936
rect 19248 26988 19300 26994
rect 19248 26930 19300 26936
rect 16856 26580 16908 26586
rect 16856 26522 16908 26528
rect 17316 26580 17368 26586
rect 17316 26522 17368 26528
rect 16868 26042 16896 26522
rect 19260 26450 19288 26930
rect 19248 26444 19300 26450
rect 19248 26386 19300 26392
rect 17868 26308 17920 26314
rect 17868 26250 17920 26256
rect 19984 26308 20036 26314
rect 19984 26250 20036 26256
rect 17880 26042 17908 26250
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 16856 26036 16908 26042
rect 16856 25978 16908 25984
rect 17868 26036 17920 26042
rect 17868 25978 17920 25984
rect 19892 25832 19944 25838
rect 19892 25774 19944 25780
rect 19904 25362 19932 25774
rect 19892 25356 19944 25362
rect 19892 25298 19944 25304
rect 16672 25288 16724 25294
rect 16672 25230 16724 25236
rect 17316 25288 17368 25294
rect 17316 25230 17368 25236
rect 17328 24750 17356 25230
rect 19248 25220 19300 25226
rect 19248 25162 19300 25168
rect 18696 25152 18748 25158
rect 18696 25094 18748 25100
rect 18708 24818 18736 25094
rect 18696 24812 18748 24818
rect 18696 24754 18748 24760
rect 17316 24744 17368 24750
rect 17316 24686 17368 24692
rect 16120 24608 16172 24614
rect 16120 24550 16172 24556
rect 15476 24268 15528 24274
rect 15476 24210 15528 24216
rect 16132 24206 16160 24550
rect 17328 24206 17356 24686
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18696 24608 18748 24614
rect 18696 24550 18748 24556
rect 12072 24200 12124 24206
rect 12072 24142 12124 24148
rect 16120 24200 16172 24206
rect 16120 24142 16172 24148
rect 17316 24200 17368 24206
rect 17316 24142 17368 24148
rect 10692 24064 10744 24070
rect 10692 24006 10744 24012
rect 11520 24064 11572 24070
rect 11520 24006 11572 24012
rect 10704 23798 10732 24006
rect 10692 23792 10744 23798
rect 10692 23734 10744 23740
rect 9312 23724 9364 23730
rect 9312 23666 9364 23672
rect 9220 23656 9272 23662
rect 9220 23598 9272 23604
rect 8944 23520 8996 23526
rect 8944 23462 8996 23468
rect 8024 23316 8076 23322
rect 8024 23258 8076 23264
rect 8956 23118 8984 23462
rect 9232 23118 9260 23598
rect 6184 23112 6236 23118
rect 6184 23054 6236 23060
rect 7012 23112 7064 23118
rect 7012 23054 7064 23060
rect 8944 23112 8996 23118
rect 8944 23054 8996 23060
rect 9220 23112 9272 23118
rect 9220 23054 9272 23060
rect 5448 22024 5500 22030
rect 5448 21966 5500 21972
rect 5460 21146 5488 21966
rect 7024 21486 7052 23054
rect 9232 22642 9260 23054
rect 9324 22778 9352 23666
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 10796 23118 10824 23462
rect 10784 23112 10836 23118
rect 10784 23054 10836 23060
rect 11532 23050 11560 24006
rect 12084 23526 12112 24142
rect 13268 24132 13320 24138
rect 13268 24074 13320 24080
rect 13280 23866 13308 24074
rect 14096 24064 14148 24070
rect 14096 24006 14148 24012
rect 16856 24064 16908 24070
rect 16856 24006 16908 24012
rect 14108 23866 14136 24006
rect 13268 23860 13320 23866
rect 13268 23802 13320 23808
rect 14096 23860 14148 23866
rect 14096 23802 14148 23808
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 15752 23724 15804 23730
rect 15752 23666 15804 23672
rect 12072 23520 12124 23526
rect 12072 23462 12124 23468
rect 12256 23520 12308 23526
rect 12256 23462 12308 23468
rect 12268 23186 12296 23462
rect 12256 23180 12308 23186
rect 12256 23122 12308 23128
rect 11520 23044 11572 23050
rect 11520 22986 11572 22992
rect 10692 22976 10744 22982
rect 10692 22918 10744 22924
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 10704 22710 10732 22918
rect 10692 22704 10744 22710
rect 10692 22646 10744 22652
rect 9220 22636 9272 22642
rect 9220 22578 9272 22584
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 7012 21480 7064 21486
rect 7012 21422 7064 21428
rect 5448 21140 5500 21146
rect 5448 21082 5500 21088
rect 7024 20942 7052 21422
rect 8484 21344 8536 21350
rect 8484 21286 8536 21292
rect 6368 20936 6420 20942
rect 6368 20878 6420 20884
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 8208 20936 8260 20942
rect 8208 20878 8260 20884
rect 5264 20868 5316 20874
rect 5264 20810 5316 20816
rect 5816 20868 5868 20874
rect 5816 20810 5868 20816
rect 4896 20460 4948 20466
rect 4896 20402 4948 20408
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 4344 20392 4396 20398
rect 4344 20334 4396 20340
rect 4080 20262 4108 20334
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 4080 19378 4108 20198
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4620 19712 4672 19718
rect 4620 19654 4672 19660
rect 1584 19372 1636 19378
rect 1584 19314 1636 19320
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 1596 18834 1624 19314
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 1584 18828 1636 18834
rect 1584 18770 1636 18776
rect 1596 18290 1624 18770
rect 2976 18766 3004 19110
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 2964 18760 3016 18766
rect 2964 18702 3016 18708
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 2976 18358 3004 18566
rect 2964 18352 3016 18358
rect 2964 18294 3016 18300
rect 4632 18290 4660 19654
rect 5552 19378 5580 20402
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 5736 19854 5764 20198
rect 5828 19854 5856 20810
rect 6380 20398 6408 20878
rect 7656 20868 7708 20874
rect 7656 20810 7708 20816
rect 7668 20602 7696 20810
rect 7748 20800 7800 20806
rect 7748 20742 7800 20748
rect 7656 20596 7708 20602
rect 7656 20538 7708 20544
rect 6368 20392 6420 20398
rect 6368 20334 6420 20340
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 5816 19848 5868 19854
rect 5816 19790 5868 19796
rect 5724 19712 5776 19718
rect 5724 19654 5776 19660
rect 5736 19446 5764 19654
rect 5724 19440 5776 19446
rect 5724 19382 5776 19388
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 6380 19310 6408 20334
rect 7760 19446 7788 20742
rect 8220 19786 8248 20878
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 8208 19780 8260 19786
rect 8208 19722 8260 19728
rect 7748 19440 7800 19446
rect 7748 19382 7800 19388
rect 8220 19378 8248 19722
rect 8208 19372 8260 19378
rect 8208 19314 8260 19320
rect 6368 19304 6420 19310
rect 6368 19246 6420 19252
rect 6380 18766 6408 19246
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7760 18766 7788 19110
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 7748 18760 7800 18766
rect 7748 18702 7800 18708
rect 6380 18290 6408 18702
rect 7748 18624 7800 18630
rect 7748 18566 7800 18572
rect 7760 18358 7788 18566
rect 7748 18352 7800 18358
rect 7748 18294 7800 18300
rect 8312 18290 8340 20402
rect 8496 19378 8524 21286
rect 8944 20936 8996 20942
rect 8944 20878 8996 20884
rect 8956 20534 8984 20878
rect 9600 20602 9628 21490
rect 10232 20868 10284 20874
rect 10232 20810 10284 20816
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9588 20596 9640 20602
rect 9588 20538 9640 20544
rect 8944 20528 8996 20534
rect 8944 20470 8996 20476
rect 8956 19854 8984 20470
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 8484 19372 8536 19378
rect 8484 19314 8536 19320
rect 8956 18766 8984 19790
rect 9588 19780 9640 19786
rect 9588 19722 9640 19728
rect 9600 19514 9628 19722
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9692 19446 9720 20742
rect 9680 19440 9732 19446
rect 9680 19382 9732 19388
rect 10244 18970 10272 20810
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 10232 18964 10284 18970
rect 10232 18906 10284 18912
rect 10336 18766 10364 19654
rect 11532 18766 11560 22986
rect 12268 22710 12296 23122
rect 13096 22778 13124 23666
rect 13820 23656 13872 23662
rect 13820 23598 13872 23604
rect 14740 23656 14792 23662
rect 14740 23598 14792 23604
rect 13832 23202 13860 23598
rect 13740 23186 13860 23202
rect 13728 23180 13860 23186
rect 13780 23174 13860 23180
rect 13728 23122 13780 23128
rect 13084 22772 13136 22778
rect 13084 22714 13136 22720
rect 12256 22704 12308 22710
rect 12256 22646 12308 22652
rect 12268 22030 12296 22646
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 12256 22024 12308 22030
rect 12256 21966 12308 21972
rect 12268 21554 12296 21966
rect 12256 21548 12308 21554
rect 12256 21490 12308 21496
rect 12268 21146 12296 21490
rect 12256 21140 12308 21146
rect 12256 21082 12308 21088
rect 11612 20392 11664 20398
rect 11612 20334 11664 20340
rect 11624 19854 11652 20334
rect 12912 20330 12940 22578
rect 13268 21956 13320 21962
rect 13268 21898 13320 21904
rect 12992 21888 13044 21894
rect 12992 21830 13044 21836
rect 13004 20534 13032 21830
rect 13280 21146 13308 21898
rect 14752 21554 14780 23598
rect 15476 23520 15528 23526
rect 15476 23462 15528 23468
rect 15488 23186 15516 23462
rect 15764 23322 15792 23666
rect 16028 23520 16080 23526
rect 16028 23462 16080 23468
rect 15752 23316 15804 23322
rect 15752 23258 15804 23264
rect 15476 23180 15528 23186
rect 15476 23122 15528 23128
rect 15488 22710 15516 23122
rect 15476 22704 15528 22710
rect 15476 22646 15528 22652
rect 15488 22098 15516 22646
rect 15752 22636 15804 22642
rect 15752 22578 15804 22584
rect 15476 22092 15528 22098
rect 15476 22034 15528 22040
rect 15764 21894 15792 22578
rect 16040 22030 16068 23462
rect 16868 23118 16896 24006
rect 17328 23186 17356 24142
rect 18052 23520 18104 23526
rect 18052 23462 18104 23468
rect 17316 23180 17368 23186
rect 17316 23122 17368 23128
rect 16856 23112 16908 23118
rect 16856 23054 16908 23060
rect 18064 23050 18092 23462
rect 18524 23322 18552 24550
rect 18708 24206 18736 24550
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 18696 24064 18748 24070
rect 18696 24006 18748 24012
rect 18708 23798 18736 24006
rect 19260 23866 19288 25162
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19996 24886 20024 26250
rect 20088 25906 20116 29106
rect 21008 28558 21036 31622
rect 21284 31482 21312 31758
rect 21272 31476 21324 31482
rect 21272 31418 21324 31424
rect 22480 31346 22508 31758
rect 23308 31346 23336 32778
rect 23860 32570 23888 34546
rect 24412 33998 24440 35022
rect 24492 34740 24544 34746
rect 24492 34682 24544 34688
rect 24676 34740 24728 34746
rect 24676 34682 24728 34688
rect 24400 33992 24452 33998
rect 24400 33934 24452 33940
rect 24412 33522 24440 33934
rect 24400 33516 24452 33522
rect 24400 33458 24452 33464
rect 24412 32910 24440 33458
rect 24400 32904 24452 32910
rect 24400 32846 24452 32852
rect 23848 32564 23900 32570
rect 23848 32506 23900 32512
rect 24504 32434 24532 34682
rect 24688 32910 24716 34682
rect 25044 34604 25096 34610
rect 25044 34546 25096 34552
rect 24860 33856 24912 33862
rect 24860 33798 24912 33804
rect 24676 32904 24728 32910
rect 24676 32846 24728 32852
rect 24492 32428 24544 32434
rect 24492 32370 24544 32376
rect 24872 31822 24900 33798
rect 25056 33658 25084 34546
rect 26252 34066 26280 35022
rect 26976 35012 27028 35018
rect 26976 34954 27028 34960
rect 28356 35012 28408 35018
rect 28356 34954 28408 34960
rect 26608 34944 26660 34950
rect 26608 34886 26660 34892
rect 26240 34060 26292 34066
rect 26240 34002 26292 34008
rect 25688 33924 25740 33930
rect 25688 33866 25740 33872
rect 26332 33924 26384 33930
rect 26332 33866 26384 33872
rect 25044 33652 25096 33658
rect 25044 33594 25096 33600
rect 25044 32836 25096 32842
rect 25044 32778 25096 32784
rect 23664 31816 23716 31822
rect 23664 31758 23716 31764
rect 24860 31816 24912 31822
rect 24860 31758 24912 31764
rect 21272 31340 21324 31346
rect 21272 31282 21324 31288
rect 22468 31340 22520 31346
rect 22468 31282 22520 31288
rect 23296 31340 23348 31346
rect 23296 31282 23348 31288
rect 21284 30394 21312 31282
rect 22480 30802 22508 31282
rect 22468 30796 22520 30802
rect 22468 30738 22520 30744
rect 22008 30592 22060 30598
rect 22008 30534 22060 30540
rect 21272 30388 21324 30394
rect 21272 30330 21324 30336
rect 21916 30252 21968 30258
rect 21916 30194 21968 30200
rect 21928 29850 21956 30194
rect 21916 29844 21968 29850
rect 21916 29786 21968 29792
rect 22020 29646 22048 30534
rect 23204 30184 23256 30190
rect 23204 30126 23256 30132
rect 22008 29640 22060 29646
rect 22008 29582 22060 29588
rect 23216 29170 23244 30126
rect 23204 29164 23256 29170
rect 23204 29106 23256 29112
rect 22468 29096 22520 29102
rect 22468 29038 22520 29044
rect 22480 28558 22508 29038
rect 23676 29034 23704 31758
rect 23756 31680 23808 31686
rect 23756 31622 23808 31628
rect 23768 30734 23796 31622
rect 25056 31278 25084 32778
rect 25700 32570 25728 33866
rect 25780 33856 25832 33862
rect 25780 33798 25832 33804
rect 25792 33590 25820 33798
rect 25780 33584 25832 33590
rect 25780 33526 25832 33532
rect 26344 33114 26372 33866
rect 26620 33590 26648 34886
rect 26884 34536 26936 34542
rect 26884 34478 26936 34484
rect 26896 34082 26924 34478
rect 26988 34202 27016 34954
rect 28368 34746 28396 34954
rect 28356 34740 28408 34746
rect 28356 34682 28408 34688
rect 28460 34678 28488 35430
rect 28448 34672 28500 34678
rect 28448 34614 28500 34620
rect 28356 34604 28408 34610
rect 28356 34546 28408 34552
rect 26976 34196 27028 34202
rect 26976 34138 27028 34144
rect 26896 34054 27016 34082
rect 26608 33584 26660 33590
rect 26608 33526 26660 33532
rect 26988 33454 27016 34054
rect 28368 33658 28396 34546
rect 28356 33652 28408 33658
rect 28356 33594 28408 33600
rect 26976 33448 27028 33454
rect 26976 33390 27028 33396
rect 26332 33108 26384 33114
rect 26332 33050 26384 33056
rect 26988 32910 27016 33390
rect 26976 32904 27028 32910
rect 26976 32846 27028 32852
rect 27528 32904 27580 32910
rect 27528 32846 27580 32852
rect 25688 32564 25740 32570
rect 25688 32506 25740 32512
rect 27540 32366 27568 32846
rect 28356 32768 28408 32774
rect 28356 32710 28408 32716
rect 27528 32360 27580 32366
rect 27528 32302 27580 32308
rect 27540 32026 27568 32302
rect 27528 32020 27580 32026
rect 27528 31962 27580 31968
rect 27068 31340 27120 31346
rect 27068 31282 27120 31288
rect 25044 31272 25096 31278
rect 25044 31214 25096 31220
rect 24584 31136 24636 31142
rect 24584 31078 24636 31084
rect 23756 30728 23808 30734
rect 23756 30670 23808 30676
rect 24492 30660 24544 30666
rect 24492 30602 24544 30608
rect 23848 30592 23900 30598
rect 23848 30534 23900 30540
rect 23860 29646 23888 30534
rect 24504 30394 24532 30602
rect 24492 30388 24544 30394
rect 24492 30330 24544 30336
rect 23848 29640 23900 29646
rect 23848 29582 23900 29588
rect 23848 29504 23900 29510
rect 23848 29446 23900 29452
rect 23860 29238 23888 29446
rect 24596 29238 24624 31078
rect 24952 30728 25004 30734
rect 24952 30670 25004 30676
rect 24964 30190 24992 30670
rect 24952 30184 25004 30190
rect 24952 30126 25004 30132
rect 24964 29238 24992 30126
rect 25056 29646 25084 31214
rect 26240 31136 26292 31142
rect 26240 31078 26292 31084
rect 26424 31136 26476 31142
rect 26424 31078 26476 31084
rect 25872 30252 25924 30258
rect 25872 30194 25924 30200
rect 25044 29640 25096 29646
rect 25044 29582 25096 29588
rect 25884 29306 25912 30194
rect 26252 30122 26280 31078
rect 26436 30326 26464 31078
rect 26424 30320 26476 30326
rect 26424 30262 26476 30268
rect 26240 30116 26292 30122
rect 26240 30058 26292 30064
rect 27080 29850 27108 31282
rect 27528 31272 27580 31278
rect 27528 31214 27580 31220
rect 27540 30734 27568 31214
rect 27528 30728 27580 30734
rect 27528 30670 27580 30676
rect 27160 30592 27212 30598
rect 27160 30534 27212 30540
rect 27068 29844 27120 29850
rect 27068 29786 27120 29792
rect 25872 29300 25924 29306
rect 25872 29242 25924 29248
rect 27172 29238 27200 30534
rect 27540 29646 27568 30670
rect 27528 29640 27580 29646
rect 27528 29582 27580 29588
rect 28368 29578 28396 32710
rect 28356 29572 28408 29578
rect 28356 29514 28408 29520
rect 23848 29232 23900 29238
rect 23848 29174 23900 29180
rect 24584 29232 24636 29238
rect 24584 29174 24636 29180
rect 24952 29232 25004 29238
rect 24952 29174 25004 29180
rect 27160 29232 27212 29238
rect 27160 29174 27212 29180
rect 25872 29164 25924 29170
rect 25872 29106 25924 29112
rect 23664 29028 23716 29034
rect 23664 28970 23716 28976
rect 20996 28552 21048 28558
rect 20996 28494 21048 28500
rect 22468 28552 22520 28558
rect 22468 28494 22520 28500
rect 25136 28552 25188 28558
rect 25136 28494 25188 28500
rect 20536 28416 20588 28422
rect 20536 28358 20588 28364
rect 20548 27606 20576 28358
rect 22480 28014 22508 28494
rect 23480 28484 23532 28490
rect 23480 28426 23532 28432
rect 23204 28416 23256 28422
rect 23204 28358 23256 28364
rect 22468 28008 22520 28014
rect 22468 27950 22520 27956
rect 20628 27872 20680 27878
rect 20628 27814 20680 27820
rect 20536 27600 20588 27606
rect 20536 27542 20588 27548
rect 20640 27470 20668 27814
rect 22480 27470 22508 27950
rect 20628 27464 20680 27470
rect 20628 27406 20680 27412
rect 22468 27464 22520 27470
rect 22468 27406 22520 27412
rect 21272 26784 21324 26790
rect 21272 26726 21324 26732
rect 21284 26382 21312 26726
rect 21272 26376 21324 26382
rect 21272 26318 21324 26324
rect 22480 26314 22508 27406
rect 23112 26988 23164 26994
rect 23112 26930 23164 26936
rect 23124 26586 23152 26930
rect 23112 26580 23164 26586
rect 23112 26522 23164 26528
rect 23216 26382 23244 28358
rect 23388 27396 23440 27402
rect 23388 27338 23440 27344
rect 23400 26926 23428 27338
rect 23492 27130 23520 28426
rect 24492 28076 24544 28082
rect 24492 28018 24544 28024
rect 24768 28076 24820 28082
rect 24768 28018 24820 28024
rect 24124 27872 24176 27878
rect 24124 27814 24176 27820
rect 24136 27470 24164 27814
rect 24124 27464 24176 27470
rect 24124 27406 24176 27412
rect 24504 27334 24532 28018
rect 23848 27328 23900 27334
rect 23848 27270 23900 27276
rect 24492 27328 24544 27334
rect 24492 27270 24544 27276
rect 23480 27124 23532 27130
rect 23480 27066 23532 27072
rect 23860 27062 23888 27270
rect 24780 27062 24808 28018
rect 25148 27470 25176 28494
rect 25884 28218 25912 29106
rect 27620 28552 27672 28558
rect 27620 28494 27672 28500
rect 27068 28484 27120 28490
rect 27068 28426 27120 28432
rect 27080 28218 27108 28426
rect 25872 28212 25924 28218
rect 25872 28154 25924 28160
rect 27068 28212 27120 28218
rect 27068 28154 27120 28160
rect 25884 27878 25912 28154
rect 27632 28150 27660 28494
rect 28080 28484 28132 28490
rect 28080 28426 28132 28432
rect 27620 28144 27672 28150
rect 27620 28086 27672 28092
rect 25872 27872 25924 27878
rect 25872 27814 25924 27820
rect 27632 27470 27660 28086
rect 28092 27946 28120 28426
rect 28356 28416 28408 28422
rect 28356 28358 28408 28364
rect 28368 28150 28396 28358
rect 28356 28144 28408 28150
rect 28356 28086 28408 28092
rect 28172 28076 28224 28082
rect 28172 28018 28224 28024
rect 28080 27940 28132 27946
rect 28080 27882 28132 27888
rect 28184 27606 28212 28018
rect 28172 27600 28224 27606
rect 28172 27542 28224 27548
rect 25136 27464 25188 27470
rect 25136 27406 25188 27412
rect 27620 27464 27672 27470
rect 27620 27406 27672 27412
rect 23848 27056 23900 27062
rect 23848 26998 23900 27004
rect 24768 27056 24820 27062
rect 24768 26998 24820 27004
rect 23388 26920 23440 26926
rect 23388 26862 23440 26868
rect 23204 26376 23256 26382
rect 23204 26318 23256 26324
rect 23400 26330 23428 26862
rect 25148 26382 25176 27406
rect 25320 27396 25372 27402
rect 25320 27338 25372 27344
rect 25332 27130 25360 27338
rect 25320 27124 25372 27130
rect 25320 27066 25372 27072
rect 25780 26988 25832 26994
rect 25780 26930 25832 26936
rect 25792 26586 25820 26930
rect 25780 26580 25832 26586
rect 25780 26522 25832 26528
rect 27632 26382 27660 27406
rect 27896 27328 27948 27334
rect 27896 27270 27948 27276
rect 27804 26988 27856 26994
rect 27804 26930 27856 26936
rect 25136 26376 25188 26382
rect 23400 26314 23520 26330
rect 25136 26318 25188 26324
rect 27620 26376 27672 26382
rect 27620 26318 27672 26324
rect 22468 26308 22520 26314
rect 22468 26250 22520 26256
rect 23388 26308 23520 26314
rect 23440 26302 23520 26308
rect 23388 26250 23440 26256
rect 21272 26240 21324 26246
rect 21272 26182 21324 26188
rect 20076 25900 20128 25906
rect 20076 25842 20128 25848
rect 20904 25900 20956 25906
rect 20904 25842 20956 25848
rect 19984 24880 20036 24886
rect 19984 24822 20036 24828
rect 19340 24132 19392 24138
rect 19340 24074 19392 24080
rect 19248 23860 19300 23866
rect 19248 23802 19300 23808
rect 18696 23792 18748 23798
rect 18696 23734 18748 23740
rect 19352 23730 19380 24074
rect 20812 24064 20864 24070
rect 20812 24006 20864 24012
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 20824 23798 20852 24006
rect 20812 23792 20864 23798
rect 20812 23734 20864 23740
rect 19340 23724 19392 23730
rect 19340 23666 19392 23672
rect 18788 23520 18840 23526
rect 18788 23462 18840 23468
rect 18512 23316 18564 23322
rect 18512 23258 18564 23264
rect 18800 23118 18828 23462
rect 18788 23112 18840 23118
rect 18788 23054 18840 23060
rect 18052 23044 18104 23050
rect 18052 22986 18104 22992
rect 18064 22642 18092 22986
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 18052 22636 18104 22642
rect 18052 22578 18104 22584
rect 20628 22636 20680 22642
rect 20628 22578 20680 22584
rect 16120 22432 16172 22438
rect 16120 22374 16172 22380
rect 15844 22024 15896 22030
rect 15844 21966 15896 21972
rect 16028 22024 16080 22030
rect 16028 21966 16080 21972
rect 15752 21888 15804 21894
rect 15752 21830 15804 21836
rect 14464 21548 14516 21554
rect 14464 21490 14516 21496
rect 14740 21548 14792 21554
rect 14740 21490 14792 21496
rect 13636 21344 13688 21350
rect 13636 21286 13688 21292
rect 13268 21140 13320 21146
rect 13268 21082 13320 21088
rect 13648 20942 13676 21286
rect 13636 20936 13688 20942
rect 13636 20878 13688 20884
rect 12992 20528 13044 20534
rect 12992 20470 13044 20476
rect 12900 20324 12952 20330
rect 12900 20266 12952 20272
rect 14476 20058 14504 21490
rect 15856 21486 15884 21966
rect 15844 21480 15896 21486
rect 15844 21422 15896 21428
rect 15856 21146 15884 21422
rect 15844 21140 15896 21146
rect 15844 21082 15896 21088
rect 14740 21004 14792 21010
rect 14740 20946 14792 20952
rect 14752 20466 14780 20946
rect 16132 20942 16160 22374
rect 18064 21554 18092 22578
rect 20640 22234 20668 22578
rect 20916 22438 20944 25842
rect 21284 25294 21312 26182
rect 23492 25974 23520 26302
rect 25504 26308 25556 26314
rect 25504 26250 25556 26256
rect 26976 26308 27028 26314
rect 26976 26250 27028 26256
rect 25516 26042 25544 26250
rect 25504 26036 25556 26042
rect 25504 25978 25556 25984
rect 23480 25968 23532 25974
rect 23480 25910 23532 25916
rect 24952 25968 25004 25974
rect 24952 25910 25004 25916
rect 23112 25900 23164 25906
rect 23112 25842 23164 25848
rect 21824 25832 21876 25838
rect 21824 25774 21876 25780
rect 21272 25288 21324 25294
rect 21272 25230 21324 25236
rect 21732 25288 21784 25294
rect 21732 25230 21784 25236
rect 21272 25152 21324 25158
rect 21272 25094 21324 25100
rect 21284 24818 21312 25094
rect 21744 24818 21772 25230
rect 21272 24812 21324 24818
rect 21272 24754 21324 24760
rect 21732 24812 21784 24818
rect 21732 24754 21784 24760
rect 21180 24608 21232 24614
rect 21180 24550 21232 24556
rect 21192 24206 21220 24550
rect 21180 24200 21232 24206
rect 21180 24142 21232 24148
rect 20996 23724 21048 23730
rect 20996 23666 21048 23672
rect 21008 22642 21036 23666
rect 21088 23112 21140 23118
rect 21088 23054 21140 23060
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 20812 22432 20864 22438
rect 20812 22374 20864 22380
rect 20904 22432 20956 22438
rect 20904 22374 20956 22380
rect 20628 22228 20680 22234
rect 20628 22170 20680 22176
rect 19156 22024 19208 22030
rect 19156 21966 19208 21972
rect 16488 21548 16540 21554
rect 16488 21490 16540 21496
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 18420 21548 18472 21554
rect 18420 21490 18472 21496
rect 16500 21146 16528 21490
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 16488 21140 16540 21146
rect 16488 21082 16540 21088
rect 16120 20936 16172 20942
rect 16120 20878 16172 20884
rect 18064 20534 18092 21286
rect 18432 21146 18460 21490
rect 18420 21140 18472 21146
rect 18420 21082 18472 21088
rect 18052 20528 18104 20534
rect 18052 20470 18104 20476
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 14464 20052 14516 20058
rect 14464 19994 14516 20000
rect 14752 19922 14780 20402
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 14740 19916 14792 19922
rect 14740 19858 14792 19864
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11624 19378 11652 19790
rect 12808 19780 12860 19786
rect 12808 19722 12860 19728
rect 12820 19378 12848 19722
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12912 19446 12940 19654
rect 12900 19440 12952 19446
rect 12900 19382 12952 19388
rect 11612 19372 11664 19378
rect 11612 19314 11664 19320
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12808 19372 12860 19378
rect 12808 19314 12860 19320
rect 13912 19372 13964 19378
rect 13912 19314 13964 19320
rect 11624 18766 11652 19314
rect 8944 18760 8996 18766
rect 8944 18702 8996 18708
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 1596 17746 1624 18226
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4632 17762 4660 18226
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 1584 17740 1636 17746
rect 1584 17682 1636 17688
rect 2504 17740 2556 17746
rect 2504 17682 2556 17688
rect 4540 17734 4660 17762
rect 2516 17202 2544 17682
rect 4540 17678 4568 17734
rect 4528 17672 4580 17678
rect 4528 17614 4580 17620
rect 3884 17604 3936 17610
rect 3884 17546 3936 17552
rect 3896 17338 3924 17546
rect 3884 17332 3936 17338
rect 3884 17274 3936 17280
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 4436 17196 4488 17202
rect 4540 17184 4568 17614
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 4488 17156 4568 17184
rect 4436 17138 4488 17144
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4632 16590 4660 17478
rect 5000 17270 5028 18022
rect 8956 17678 8984 18702
rect 11624 18290 11652 18702
rect 12728 18426 12756 19314
rect 13924 18766 13952 19314
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 11612 18284 11664 18290
rect 11612 18226 11664 18232
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 4988 17264 5040 17270
rect 4988 17206 5040 17212
rect 5460 17202 5488 17614
rect 7748 17604 7800 17610
rect 7748 17546 7800 17552
rect 7760 17338 7788 17546
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 5172 17196 5224 17202
rect 5172 17138 5224 17144
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 2688 16584 2740 16590
rect 2688 16526 2740 16532
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 2700 16046 2728 16526
rect 4724 16182 4752 16934
rect 5184 16794 5212 17138
rect 7024 16794 7052 17138
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 5552 16046 5580 16526
rect 7748 16516 7800 16522
rect 7748 16458 7800 16464
rect 7760 16250 7788 16458
rect 8404 16250 8432 17478
rect 8956 17270 8984 17614
rect 9416 17338 9444 18226
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 8944 17264 8996 17270
rect 8944 17206 8996 17212
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9324 16522 9352 16730
rect 9312 16516 9364 16522
rect 9312 16458 9364 16464
rect 9416 16250 9444 17138
rect 9600 16590 9628 18022
rect 11624 17678 11652 18226
rect 11612 17672 11664 17678
rect 11612 17614 11664 17620
rect 10232 17604 10284 17610
rect 10232 17546 10284 17552
rect 10244 16794 10272 17546
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 11348 16590 11376 17478
rect 11624 17202 11652 17614
rect 12912 17338 12940 18226
rect 13924 18170 13952 18702
rect 14016 18358 14044 19110
rect 14004 18352 14056 18358
rect 14004 18294 14056 18300
rect 14108 18290 14136 19858
rect 16132 19854 16160 20198
rect 18708 20058 18736 20402
rect 19168 20330 19196 21966
rect 20536 21956 20588 21962
rect 20536 21898 20588 21904
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19892 21344 19944 21350
rect 19892 21286 19944 21292
rect 19248 21004 19300 21010
rect 19248 20946 19300 20952
rect 19260 20482 19288 20946
rect 19904 20942 19932 21286
rect 20548 21146 20576 21898
rect 20628 21548 20680 21554
rect 20628 21490 20680 21496
rect 20536 21140 20588 21146
rect 20536 21082 20588 21088
rect 19892 20936 19944 20942
rect 19892 20878 19944 20884
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 20640 20602 20668 21490
rect 20824 20874 20852 22374
rect 20812 20868 20864 20874
rect 20812 20810 20864 20816
rect 20916 20806 20944 22374
rect 20904 20800 20956 20806
rect 20904 20742 20956 20748
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 19260 20466 19380 20482
rect 19260 20460 19392 20466
rect 19260 20454 19340 20460
rect 19340 20402 19392 20408
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 19156 20324 19208 20330
rect 19156 20266 19208 20272
rect 18696 20052 18748 20058
rect 18696 19994 18748 20000
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 17316 19848 17368 19854
rect 19168 19836 19196 20266
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19352 19854 19380 20198
rect 20640 20058 20668 20402
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 19248 19848 19300 19854
rect 19168 19808 19248 19836
rect 17316 19790 17368 19796
rect 19248 19790 19300 19796
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 17328 19378 17356 19790
rect 18696 19780 18748 19786
rect 18696 19722 18748 19728
rect 18708 19514 18736 19722
rect 19260 19514 19288 19790
rect 20916 19786 20944 20742
rect 20904 19780 20956 19786
rect 20904 19722 20956 19728
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 20720 19440 20772 19446
rect 20720 19382 20772 19388
rect 17316 19372 17368 19378
rect 17316 19314 17368 19320
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 14740 18692 14792 18698
rect 14740 18634 14792 18640
rect 14752 18426 14780 18634
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 14740 18420 14792 18426
rect 14740 18362 14792 18368
rect 14096 18284 14148 18290
rect 14096 18226 14148 18232
rect 13924 18142 14044 18170
rect 12900 17332 12952 17338
rect 12900 17274 12952 17280
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 12176 16794 12204 17138
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 14016 16658 14044 18142
rect 14108 17746 14136 18226
rect 14096 17740 14148 17746
rect 14096 17682 14148 17688
rect 14108 17202 14136 17682
rect 15580 17678 15608 18566
rect 17328 18222 17356 19314
rect 19260 18426 19288 19314
rect 20732 18766 20760 19382
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 20536 18352 20588 18358
rect 20536 18294 20588 18300
rect 17316 18216 17368 18222
rect 17316 18158 17368 18164
rect 17328 17678 17356 18158
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 15844 17604 15896 17610
rect 15844 17546 15896 17552
rect 15476 17536 15528 17542
rect 15476 17478 15528 17484
rect 15752 17536 15804 17542
rect 15752 17478 15804 17484
rect 15488 17270 15516 17478
rect 15476 17264 15528 17270
rect 15476 17206 15528 17212
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 14004 16652 14056 16658
rect 14004 16594 14056 16600
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 11336 16584 11388 16590
rect 11336 16526 11388 16532
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 2688 16040 2740 16046
rect 2688 15982 2740 15988
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 2872 15904 2924 15910
rect 2872 15846 2924 15852
rect 1780 15502 1808 15846
rect 2884 15502 2912 15846
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 5552 15502 5580 15982
rect 6932 15706 6960 16050
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 10428 15502 10456 16526
rect 14016 15570 14044 16594
rect 15488 16590 15516 16934
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 15764 16182 15792 17478
rect 15856 16794 15884 17546
rect 17328 17202 17356 17614
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 15752 16176 15804 16182
rect 15752 16118 15804 16124
rect 16684 16114 16712 16526
rect 17328 16114 17356 17138
rect 18524 16794 18552 17138
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 19156 16584 19208 16590
rect 19156 16526 19208 16532
rect 19168 16114 19196 16526
rect 19248 16516 19300 16522
rect 19248 16458 19300 16464
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 17316 16108 17368 16114
rect 17316 16050 17368 16056
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 14004 15564 14056 15570
rect 14004 15506 14056 15512
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 1780 15026 1808 15438
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3252 15094 3280 15302
rect 3240 15088 3292 15094
rect 3240 15030 3292 15036
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1780 14414 1808 14962
rect 3056 14816 3108 14822
rect 3056 14758 3108 14764
rect 3068 14414 3096 14758
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 1768 14408 1820 14414
rect 1768 14350 1820 14356
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 1780 13938 1808 14350
rect 5552 14278 5580 15438
rect 7932 15428 7984 15434
rect 7932 15370 7984 15376
rect 7944 15162 7972 15370
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 9784 15094 9812 15438
rect 12164 15428 12216 15434
rect 12164 15370 12216 15376
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 9772 15088 9824 15094
rect 9772 15030 9824 15036
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6288 14414 6316 14894
rect 8128 14618 8156 14962
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 3056 14272 3108 14278
rect 3056 14214 3108 14220
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 3068 14006 3096 14214
rect 3056 14000 3108 14006
rect 3056 13942 3108 13948
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 1780 13818 1808 13874
rect 1780 13790 1900 13818
rect 1872 13326 1900 13790
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 3068 13326 3096 13670
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 5552 13326 5580 14214
rect 6288 13870 6316 14350
rect 7932 14340 7984 14346
rect 7932 14282 7984 14288
rect 7944 14074 7972 14282
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 6276 13864 6328 13870
rect 6276 13806 6328 13812
rect 6288 13326 6316 13806
rect 8220 13530 8248 13874
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 1872 12850 1900 13262
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 3252 12918 3280 13126
rect 3240 12912 3292 12918
rect 3240 12854 3292 12860
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3896 12238 3924 12718
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3896 11762 3924 12174
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 4264 11898 4292 12106
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 5368 11830 5396 12582
rect 5552 12238 5580 13262
rect 5816 13252 5868 13258
rect 5816 13194 5868 13200
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 5644 12306 5672 12718
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5356 11824 5408 11830
rect 5356 11766 5408 11772
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 5828 11354 5856 13194
rect 6288 12782 6316 13262
rect 7748 13252 7800 13258
rect 7748 13194 7800 13200
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6276 12776 6328 12782
rect 6276 12718 6328 12724
rect 6092 12164 6144 12170
rect 6092 12106 6144 12112
rect 6104 11694 6132 12106
rect 6380 11830 6408 13126
rect 7760 12986 7788 13194
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 6104 11082 6132 11630
rect 7024 11150 7052 12038
rect 7760 11898 7788 12786
rect 9692 12238 9720 14758
rect 9784 13734 9812 15030
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10796 13870 10824 14214
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9784 13326 9812 13670
rect 10796 13326 10824 13806
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 9784 12986 9812 13262
rect 10324 13184 10376 13190
rect 10324 13126 10376 13132
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9784 12442 9812 12922
rect 10336 12918 10364 13126
rect 10980 12986 11008 14962
rect 11060 14408 11112 14414
rect 11112 14368 11192 14396
rect 11060 14350 11112 14356
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 11072 13326 11100 13670
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10324 12912 10376 12918
rect 10324 12854 10376 12860
rect 11164 12442 11192 14368
rect 11808 13258 11836 15302
rect 12176 13530 12204 15370
rect 14292 15026 14320 16050
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15764 15502 15792 15846
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15764 15094 15792 15302
rect 15752 15088 15804 15094
rect 15752 15030 15804 15036
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 12268 14414 12296 14894
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 13648 13938 13676 14758
rect 14188 14408 14240 14414
rect 14108 14368 14188 14396
rect 14108 13938 14136 14368
rect 14292 14396 14320 14962
rect 14240 14368 14320 14396
rect 14188 14350 14240 14356
rect 14556 14340 14608 14346
rect 14556 14282 14608 14288
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 13636 13932 13688 13938
rect 13636 13874 13688 13880
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9784 11898 9812 12378
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 10796 11830 10824 12038
rect 10784 11824 10836 11830
rect 10784 11766 10836 11772
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10796 11150 10824 11494
rect 11164 11354 11192 12378
rect 13832 12238 13860 12718
rect 14200 12238 14228 14214
rect 14568 12986 14596 14282
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 15304 12442 15332 13194
rect 15396 12442 15424 14962
rect 16684 14958 16712 16050
rect 18708 15706 18736 16050
rect 18696 15700 18748 15706
rect 18696 15642 18748 15648
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17328 14958 17356 15438
rect 18788 15428 18840 15434
rect 18788 15370 18840 15376
rect 18800 15162 18828 15370
rect 18788 15156 18840 15162
rect 18788 15098 18840 15104
rect 19168 15026 19196 16050
rect 19260 15162 19288 16458
rect 19352 16250 19380 16934
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 20548 16250 20576 18294
rect 20732 17270 20760 18566
rect 20904 18080 20956 18086
rect 20904 18022 20956 18028
rect 20916 17678 20944 18022
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20916 17202 20944 17614
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20916 16046 20944 16526
rect 20904 16040 20956 16046
rect 20904 15982 20956 15988
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19248 15156 19300 15162
rect 19248 15098 19300 15104
rect 19352 15026 19380 15846
rect 20916 15706 20944 15982
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 19432 15428 19484 15434
rect 19432 15370 19484 15376
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 19156 15020 19208 15026
rect 19156 14962 19208 14968
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 16672 14952 16724 14958
rect 16672 14894 16724 14900
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15672 14414 15700 14758
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15488 14006 15516 14214
rect 15476 14000 15528 14006
rect 15476 13942 15528 13948
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 12918 15516 13670
rect 16684 13190 16712 14894
rect 18524 14618 18552 14962
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 19168 14482 19196 14962
rect 19156 14476 19208 14482
rect 19156 14418 19208 14424
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16776 13938 16804 14350
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16672 13184 16724 13190
rect 16672 13126 16724 13132
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 16684 12238 16712 13126
rect 16776 12850 16804 13874
rect 19168 13870 19196 14418
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 19156 13864 19208 13870
rect 19156 13806 19208 13812
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 14188 12232 14240 12238
rect 14188 12174 14240 12180
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12176 11354 12204 11630
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12072 11280 12124 11286
rect 12072 11222 12124 11228
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10980 11082 11008 11154
rect 12084 11098 12112 11222
rect 13832 11218 13860 12174
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 14016 11354 14044 11630
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 6092 11076 6144 11082
rect 6092 11018 6144 11024
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 10968 11076 11020 11082
rect 12084 11070 12480 11098
rect 10968 11018 11020 11024
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 6104 10130 6132 11018
rect 9876 10674 9904 11018
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10796 10742 10824 10950
rect 10784 10736 10836 10742
rect 10784 10678 10836 10684
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 9876 10266 9904 10610
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 5920 9042 5948 9454
rect 7300 9178 7328 9930
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 5368 8514 5396 8978
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5460 8566 5488 8774
rect 5276 8498 5396 8514
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5264 8492 5396 8498
rect 5316 8486 5396 8492
rect 5264 8434 5316 8440
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 5368 7886 5396 8486
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 1872 7410 1900 7822
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3252 7478 3280 7686
rect 3240 7472 3292 7478
rect 3240 7414 3292 7420
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1872 6914 1900 7346
rect 4172 7290 4200 7822
rect 5368 7546 5396 7822
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 3988 7262 4200 7290
rect 1872 6886 1992 6914
rect 1964 6798 1992 6886
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 1964 6322 1992 6734
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3252 6390 3280 6598
rect 3240 6384 3292 6390
rect 3240 6326 3292 6332
rect 3988 6322 4016 7262
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 4080 6914 4108 7142
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4080 6886 4200 6914
rect 4172 6390 4200 6886
rect 5460 6798 5488 8298
rect 5644 8090 5672 8842
rect 7484 8566 7512 9862
rect 9048 9518 9076 10066
rect 10704 10062 10732 10406
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10520 9654 10548 9862
rect 10508 9648 10560 9654
rect 10508 9590 10560 9596
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 7760 8974 7788 9318
rect 9232 8974 9260 9318
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 7472 8560 7524 8566
rect 7472 8502 7524 8508
rect 8680 8430 8708 8910
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10428 8634 10456 8842
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10612 8566 10640 9862
rect 10796 8786 10824 10542
rect 10980 10130 11008 11018
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10980 9058 11008 10066
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 11072 9178 11100 9930
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 10888 9030 11008 9058
rect 10888 8974 10916 9030
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10704 8758 10824 8786
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5920 7886 5948 8366
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7760 7886 7788 8230
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 5920 7342 5948 7822
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 6564 7002 6592 7754
rect 7196 7472 7248 7478
rect 7196 7414 7248 7420
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6748 6798 6776 7278
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 5264 6724 5316 6730
rect 5264 6666 5316 6672
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5276 6458 5304 6666
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 1964 5234 1992 6258
rect 3988 5778 4016 6258
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 3988 5166 4016 5714
rect 4080 5710 4108 6054
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 5828 5778 5856 6666
rect 7208 6322 7236 7414
rect 8680 7410 8708 8366
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8404 7002 8432 7346
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8680 6798 8708 7346
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 7748 6724 7800 6730
rect 7748 6666 7800 6672
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5368 5234 5396 5510
rect 5828 5234 5856 5714
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 3988 4282 4016 5102
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4622 4108 4966
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 5828 4706 5856 5170
rect 5736 4678 5856 4706
rect 5736 4622 5764 4678
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 5184 4146 5212 4422
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5552 4010 5580 4490
rect 5736 4146 5764 4558
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 5736 3738 5764 4082
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 6012 3534 6040 4422
rect 6104 3738 6132 5578
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 7208 5302 7236 5510
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7392 4146 7420 4966
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7760 4010 7788 6666
rect 8680 6458 8708 6734
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8864 6390 8892 7142
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 8852 6384 8904 6390
rect 8852 6326 8904 6332
rect 8956 6254 8984 6734
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8956 5778 8984 6190
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 8956 5234 8984 5714
rect 9968 5710 9996 7142
rect 10704 6798 10732 8758
rect 11808 8090 11836 10610
rect 12452 9654 12480 11070
rect 13832 10606 13860 11154
rect 13912 11076 13964 11082
rect 13912 11018 13964 11024
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13924 10266 13952 11018
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 14016 10044 14044 11290
rect 14096 11280 14148 11286
rect 14096 11222 14148 11228
rect 14108 10742 14136 11222
rect 15396 11150 15424 11494
rect 15488 11354 15516 11698
rect 16684 11694 16712 12174
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 16684 11354 16712 11630
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15212 10810 15240 11018
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 16776 10674 16804 12786
rect 17224 12164 17276 12170
rect 17224 12106 17276 12112
rect 17236 11354 17264 12106
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17328 11830 17356 12038
rect 17316 11824 17368 11830
rect 17316 11766 17368 11772
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14096 10056 14148 10062
rect 14016 10016 14096 10044
rect 14096 9998 14148 10004
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12176 8566 12204 8774
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 12176 7886 12204 8366
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 10244 5914 10272 6666
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 10336 5302 10364 6598
rect 10704 5778 10732 6734
rect 10796 6458 10824 7346
rect 12176 7206 12204 7822
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12176 6798 12204 7142
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 12164 6792 12216 6798
rect 12164 6734 12216 6740
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 11900 6322 11928 6734
rect 12268 6458 12296 7754
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12452 6322 12480 9590
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12820 8634 12848 9522
rect 14108 9382 14136 9998
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14108 8974 14136 9318
rect 14384 8974 14412 10406
rect 16672 10056 16724 10062
rect 16776 10044 16804 10610
rect 17972 10266 18000 12786
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 18064 10742 18092 11494
rect 18052 10736 18104 10742
rect 18052 10678 18104 10684
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 18064 10062 18092 10406
rect 16724 10016 16804 10044
rect 18052 10056 18104 10062
rect 16672 9998 16724 10004
rect 18052 9998 18104 10004
rect 15476 9988 15528 9994
rect 15476 9930 15528 9936
rect 15488 9178 15516 9930
rect 16684 9586 16712 9998
rect 18156 9654 18184 12582
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 14108 8430 14136 8910
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13084 7812 13136 7818
rect 13084 7754 13136 7760
rect 13096 7002 13124 7754
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 13556 6390 13584 7686
rect 13832 7478 13860 8230
rect 13820 7472 13872 7478
rect 13820 7414 13872 7420
rect 14108 7206 14136 8366
rect 14832 7812 14884 7818
rect 14832 7754 14884 7760
rect 14844 7410 14872 7754
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14108 6866 14136 7142
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14292 6798 14320 7142
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 13544 6384 13596 6390
rect 13544 6326 13596 6332
rect 14752 6322 14780 6802
rect 15856 6390 15884 7686
rect 16040 6458 16068 8434
rect 16684 7970 16712 9522
rect 18248 9450 18276 13806
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19248 11076 19300 11082
rect 19248 11018 19300 11024
rect 19260 10742 19288 11018
rect 19248 10736 19300 10742
rect 19248 10678 19300 10684
rect 19352 10606 19380 11086
rect 19340 10600 19392 10606
rect 19340 10542 19392 10548
rect 18604 10464 18656 10470
rect 18604 10406 18656 10412
rect 18616 10062 18644 10406
rect 19352 10266 19380 10542
rect 19340 10260 19392 10266
rect 19340 10202 19392 10208
rect 18604 10056 18656 10062
rect 18604 9998 18656 10004
rect 18236 9444 18288 9450
rect 18236 9386 18288 9392
rect 17316 8424 17368 8430
rect 17316 8366 17368 8372
rect 16684 7942 16896 7970
rect 16868 7886 16896 7942
rect 17328 7886 17356 8366
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 16212 7812 16264 7818
rect 16212 7754 16264 7760
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 16132 6798 16160 7142
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 15844 6384 15896 6390
rect 15844 6326 15896 6332
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10324 5296 10376 5302
rect 10324 5238 10376 5244
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9784 4690 9812 5170
rect 10704 5030 10732 5714
rect 11060 5636 11112 5642
rect 11060 5578 11112 5584
rect 11072 5370 11100 5578
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10704 4706 10732 4966
rect 10704 4690 10824 4706
rect 9772 4684 9824 4690
rect 10704 4684 10836 4690
rect 10704 4678 10784 4684
rect 9772 4626 9824 4632
rect 10784 4626 10836 4632
rect 10796 4146 10824 4626
rect 11164 4622 11192 5510
rect 12452 5302 12480 6258
rect 16224 5914 16252 7754
rect 17328 7410 17356 7822
rect 18328 7812 18380 7818
rect 18328 7754 18380 7760
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17696 7478 17724 7686
rect 17684 7472 17736 7478
rect 17684 7414 17736 7420
rect 17316 7404 17368 7410
rect 17316 7346 17368 7352
rect 17328 6866 17356 7346
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 16304 6248 16356 6254
rect 16304 6190 16356 6196
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 16316 5778 16344 6190
rect 16304 5772 16356 5778
rect 16304 5714 16356 5720
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 13740 5166 13768 5646
rect 15476 5636 15528 5642
rect 15476 5578 15528 5584
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 7748 4004 7800 4010
rect 7748 3946 7800 3952
rect 10796 3738 10824 4082
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 10796 3058 10824 3674
rect 11256 3534 11284 4422
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 11808 3738 11836 4082
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 12912 3126 12940 3878
rect 12900 3120 12952 3126
rect 12900 3062 12952 3068
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 11532 2514 11560 2994
rect 12900 2848 12952 2854
rect 12900 2790 12952 2796
rect 11520 2508 11572 2514
rect 11520 2450 11572 2456
rect 12912 2446 12940 2790
rect 13096 2582 13124 4082
rect 13372 4078 13400 4558
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 13372 3602 13400 4014
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 13372 3058 13400 3538
rect 13832 3126 13860 4966
rect 14752 4282 14780 5170
rect 15488 4826 15516 5578
rect 16316 4826 16344 5714
rect 16592 5710 16620 6598
rect 18340 6458 18368 7754
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 15476 4548 15528 4554
rect 15476 4490 15528 4496
rect 14740 4276 14792 4282
rect 14740 4218 14792 4224
rect 15488 3738 15516 4490
rect 16316 4146 16344 4762
rect 16776 4146 16804 5510
rect 18616 5234 18644 9998
rect 19352 9518 19380 10202
rect 19444 10062 19472 15370
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 20812 13728 20864 13734
rect 20812 13670 20864 13676
rect 20824 13326 20852 13670
rect 20812 13320 20864 13326
rect 20732 13280 20812 13308
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 20732 12850 20760 13280
rect 20812 13262 20864 13268
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 21008 11914 21036 22578
rect 21100 22030 21128 23054
rect 21180 23044 21232 23050
rect 21180 22986 21232 22992
rect 21088 22024 21140 22030
rect 21088 21966 21140 21972
rect 21100 20942 21128 21966
rect 21192 21894 21220 22986
rect 21744 22642 21772 24754
rect 21836 24206 21864 25774
rect 23124 25498 23152 25842
rect 24492 25696 24544 25702
rect 24492 25638 24544 25644
rect 23112 25492 23164 25498
rect 23112 25434 23164 25440
rect 23204 25220 23256 25226
rect 23204 25162 23256 25168
rect 23216 24954 23244 25162
rect 23204 24948 23256 24954
rect 23204 24890 23256 24896
rect 23204 24812 23256 24818
rect 23204 24754 23256 24760
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 21836 23730 21864 24142
rect 23112 24132 23164 24138
rect 23112 24074 23164 24080
rect 22652 24064 22704 24070
rect 22652 24006 22704 24012
rect 22664 23798 22692 24006
rect 22652 23792 22704 23798
rect 22652 23734 22704 23740
rect 21824 23724 21876 23730
rect 21824 23666 21876 23672
rect 22836 23044 22888 23050
rect 22836 22986 22888 22992
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22468 22976 22520 22982
rect 22468 22918 22520 22924
rect 21732 22636 21784 22642
rect 21732 22578 21784 22584
rect 21744 22030 21772 22578
rect 21732 22024 21784 22030
rect 21732 21966 21784 21972
rect 21180 21888 21232 21894
rect 21180 21830 21232 21836
rect 21744 21554 21772 21966
rect 22112 21622 22140 22918
rect 22480 22710 22508 22918
rect 22468 22704 22520 22710
rect 22468 22646 22520 22652
rect 22848 21690 22876 22986
rect 23124 22778 23152 24074
rect 23216 23866 23244 24754
rect 24124 24744 24176 24750
rect 24124 24686 24176 24692
rect 23204 23860 23256 23866
rect 23204 23802 23256 23808
rect 24136 23662 24164 24686
rect 24504 24206 24532 25638
rect 24964 25294 24992 25910
rect 26988 25906 27016 26250
rect 25504 25900 25556 25906
rect 25504 25842 25556 25848
rect 26976 25900 27028 25906
rect 26976 25842 27028 25848
rect 27712 25900 27764 25906
rect 27712 25842 27764 25848
rect 24952 25288 25004 25294
rect 24952 25230 25004 25236
rect 25320 25220 25372 25226
rect 25320 25162 25372 25168
rect 25332 24410 25360 25162
rect 25516 24954 25544 25842
rect 27620 25152 27672 25158
rect 27620 25094 27672 25100
rect 25504 24948 25556 24954
rect 25504 24890 25556 24896
rect 25504 24812 25556 24818
rect 25504 24754 25556 24760
rect 25320 24404 25372 24410
rect 25320 24346 25372 24352
rect 24492 24200 24544 24206
rect 24492 24142 24544 24148
rect 25516 23866 25544 24754
rect 26240 24744 26292 24750
rect 26240 24686 26292 24692
rect 26252 24206 26280 24686
rect 27632 24206 27660 25094
rect 26240 24200 26292 24206
rect 26240 24142 26292 24148
rect 27620 24200 27672 24206
rect 27620 24142 27672 24148
rect 25504 23860 25556 23866
rect 25504 23802 25556 23808
rect 25780 23724 25832 23730
rect 25780 23666 25832 23672
rect 24124 23656 24176 23662
rect 24124 23598 24176 23604
rect 24136 23118 24164 23598
rect 25792 23322 25820 23666
rect 26252 23662 26280 24142
rect 27620 24064 27672 24070
rect 27620 24006 27672 24012
rect 27632 23798 27660 24006
rect 27620 23792 27672 23798
rect 27620 23734 27672 23740
rect 26240 23656 26292 23662
rect 26240 23598 26292 23604
rect 27620 23520 27672 23526
rect 27620 23462 27672 23468
rect 25780 23316 25832 23322
rect 25780 23258 25832 23264
rect 24124 23112 24176 23118
rect 24124 23054 24176 23060
rect 23112 22772 23164 22778
rect 23112 22714 23164 22720
rect 24136 22710 24164 23054
rect 27632 23050 27660 23462
rect 27724 23322 27752 25842
rect 27712 23316 27764 23322
rect 27712 23258 27764 23264
rect 25136 23044 25188 23050
rect 25136 22986 25188 22992
rect 27620 23044 27672 23050
rect 27620 22986 27672 22992
rect 25148 22778 25176 22986
rect 25136 22772 25188 22778
rect 25136 22714 25188 22720
rect 24124 22704 24176 22710
rect 24124 22646 24176 22652
rect 25780 22636 25832 22642
rect 25780 22578 25832 22584
rect 25792 22234 25820 22578
rect 25964 22568 26016 22574
rect 25964 22510 26016 22516
rect 25780 22228 25832 22234
rect 25780 22170 25832 22176
rect 23204 21956 23256 21962
rect 23204 21898 23256 21904
rect 25136 21956 25188 21962
rect 25136 21898 25188 21904
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 22100 21616 22152 21622
rect 22100 21558 22152 21564
rect 21732 21548 21784 21554
rect 21732 21490 21784 21496
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 21100 20534 21128 20878
rect 21088 20528 21140 20534
rect 21088 20470 21140 20476
rect 21744 20466 21772 21490
rect 22468 20800 22520 20806
rect 22468 20742 22520 20748
rect 22480 20534 22508 20742
rect 23216 20602 23244 21898
rect 25148 21690 25176 21898
rect 25136 21684 25188 21690
rect 25136 21626 25188 21632
rect 25780 21548 25832 21554
rect 25780 21490 25832 21496
rect 24492 21344 24544 21350
rect 24492 21286 24544 21292
rect 24504 20942 24532 21286
rect 25792 21146 25820 21490
rect 25780 21140 25832 21146
rect 25780 21082 25832 21088
rect 24492 20936 24544 20942
rect 24492 20878 24544 20884
rect 23204 20596 23256 20602
rect 23204 20538 23256 20544
rect 22468 20528 22520 20534
rect 22468 20470 22520 20476
rect 21732 20460 21784 20466
rect 21732 20402 21784 20408
rect 21744 20058 21772 20402
rect 24504 20398 24532 20878
rect 25688 20868 25740 20874
rect 25688 20810 25740 20816
rect 24492 20392 24544 20398
rect 24492 20334 24544 20340
rect 21732 20052 21784 20058
rect 21732 19994 21784 20000
rect 21272 19372 21324 19378
rect 21272 19314 21324 19320
rect 21284 18426 21312 19314
rect 21744 18766 21772 19994
rect 24504 19854 24532 20334
rect 25700 20058 25728 20810
rect 25872 20256 25924 20262
rect 25872 20198 25924 20204
rect 25688 20052 25740 20058
rect 25688 19994 25740 20000
rect 25884 19854 25912 20198
rect 23664 19848 23716 19854
rect 23664 19790 23716 19796
rect 24492 19848 24544 19854
rect 24492 19790 24544 19796
rect 25872 19848 25924 19854
rect 25872 19790 25924 19796
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 23480 19372 23532 19378
rect 23480 19314 23532 19320
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 21744 18290 21772 18702
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 21732 18284 21784 18290
rect 21732 18226 21784 18232
rect 21284 17338 21312 18226
rect 21744 17678 21772 18226
rect 21732 17672 21784 17678
rect 21732 17614 21784 17620
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21836 17202 21864 19314
rect 23204 19168 23256 19174
rect 23204 19110 23256 19116
rect 22284 18692 22336 18698
rect 22284 18634 22336 18640
rect 22296 17882 22324 18634
rect 23216 18358 23244 19110
rect 23204 18352 23256 18358
rect 23204 18294 23256 18300
rect 23492 18154 23520 19314
rect 23676 19310 23704 19790
rect 25976 19786 26004 22510
rect 27632 22438 27660 22986
rect 27816 22710 27844 26930
rect 27908 26382 27936 27270
rect 27896 26376 27948 26382
rect 27896 26318 27948 26324
rect 28552 26234 28580 37946
rect 29092 37800 29144 37806
rect 29092 37742 29144 37748
rect 29104 36786 29132 37742
rect 29656 37262 29684 39578
rect 30024 38350 30052 40870
rect 30208 40730 30236 41006
rect 30196 40724 30248 40730
rect 30196 40666 30248 40672
rect 30392 40066 30420 41414
rect 30300 40050 30420 40066
rect 30288 40044 30420 40050
rect 30340 40038 30420 40044
rect 30288 39986 30340 39992
rect 30196 39976 30248 39982
rect 30196 39918 30248 39924
rect 30208 39438 30236 39918
rect 30196 39432 30248 39438
rect 30196 39374 30248 39380
rect 30208 38962 30236 39374
rect 30288 39364 30340 39370
rect 30288 39306 30340 39312
rect 30196 38956 30248 38962
rect 30196 38898 30248 38904
rect 30012 38344 30064 38350
rect 30012 38286 30064 38292
rect 30208 38282 30236 38898
rect 30196 38276 30248 38282
rect 30196 38218 30248 38224
rect 30300 38010 30328 39306
rect 30840 38752 30892 38758
rect 30840 38694 30892 38700
rect 30288 38004 30340 38010
rect 30288 37946 30340 37952
rect 29552 37256 29604 37262
rect 29552 37198 29604 37204
rect 29644 37256 29696 37262
rect 29644 37198 29696 37204
rect 29092 36780 29144 36786
rect 29092 36722 29144 36728
rect 28908 36576 28960 36582
rect 28908 36518 28960 36524
rect 28920 35834 28948 36518
rect 29104 36242 29132 36722
rect 29092 36236 29144 36242
rect 29092 36178 29144 36184
rect 29564 35834 29592 37198
rect 29828 36576 29880 36582
rect 29828 36518 29880 36524
rect 28908 35828 28960 35834
rect 28908 35770 28960 35776
rect 29552 35828 29604 35834
rect 29552 35770 29604 35776
rect 28920 35630 28948 35770
rect 28908 35624 28960 35630
rect 28908 35566 28960 35572
rect 28920 35154 28948 35566
rect 28908 35148 28960 35154
rect 28908 35090 28960 35096
rect 28920 34066 28948 35090
rect 28908 34060 28960 34066
rect 28908 34002 28960 34008
rect 29840 33998 29868 36518
rect 29920 36032 29972 36038
rect 29920 35974 29972 35980
rect 29932 35834 29960 35974
rect 29920 35828 29972 35834
rect 29920 35770 29972 35776
rect 29932 34610 29960 35770
rect 30196 35692 30248 35698
rect 30196 35634 30248 35640
rect 30208 34746 30236 35634
rect 30288 35488 30340 35494
rect 30288 35430 30340 35436
rect 30300 35086 30328 35430
rect 30288 35080 30340 35086
rect 30288 35022 30340 35028
rect 30380 34944 30432 34950
rect 30380 34886 30432 34892
rect 30196 34740 30248 34746
rect 30196 34682 30248 34688
rect 29920 34604 29972 34610
rect 29920 34546 29972 34552
rect 29828 33992 29880 33998
rect 29828 33934 29880 33940
rect 29932 33522 29960 34546
rect 30392 33590 30420 34886
rect 30380 33584 30432 33590
rect 30380 33526 30432 33532
rect 29920 33516 29972 33522
rect 29920 33458 29972 33464
rect 29932 32978 29960 33458
rect 29920 32972 29972 32978
rect 29920 32914 29972 32920
rect 28632 32836 28684 32842
rect 28632 32778 28684 32784
rect 28644 29306 28672 32778
rect 29932 32434 29960 32914
rect 29092 32428 29144 32434
rect 29092 32370 29144 32376
rect 29920 32428 29972 32434
rect 29920 32370 29972 32376
rect 29000 30592 29052 30598
rect 29000 30534 29052 30540
rect 28908 30252 28960 30258
rect 28828 30212 28908 30240
rect 28828 29714 28856 30212
rect 28908 30194 28960 30200
rect 28816 29708 28868 29714
rect 28816 29650 28868 29656
rect 28632 29300 28684 29306
rect 28632 29242 28684 29248
rect 28828 29102 28856 29650
rect 29012 29646 29040 30534
rect 29104 29850 29132 32370
rect 29276 32224 29328 32230
rect 29276 32166 29328 32172
rect 29288 30666 29316 32166
rect 30852 31482 30880 38694
rect 31128 38554 31156 41482
rect 32036 41472 32088 41478
rect 32036 41414 32088 41420
rect 31576 41132 31628 41138
rect 31576 41074 31628 41080
rect 31588 40186 31616 41074
rect 31760 40928 31812 40934
rect 31760 40870 31812 40876
rect 31576 40180 31628 40186
rect 31576 40122 31628 40128
rect 31576 40044 31628 40050
rect 31576 39986 31628 39992
rect 31588 39098 31616 39986
rect 31772 39438 31800 40870
rect 32048 40526 32076 41414
rect 32140 41070 32168 41550
rect 32404 41540 32456 41546
rect 32404 41482 32456 41488
rect 32128 41064 32180 41070
rect 32128 41006 32180 41012
rect 32140 40730 32168 41006
rect 32128 40724 32180 40730
rect 32128 40666 32180 40672
rect 32036 40520 32088 40526
rect 32036 40462 32088 40468
rect 32312 40452 32364 40458
rect 32312 40394 32364 40400
rect 31944 40384 31996 40390
rect 31944 40326 31996 40332
rect 31760 39432 31812 39438
rect 31760 39374 31812 39380
rect 31576 39092 31628 39098
rect 31576 39034 31628 39040
rect 31956 39030 31984 40326
rect 31944 39024 31996 39030
rect 31944 38966 31996 38972
rect 31116 38548 31168 38554
rect 31116 38490 31168 38496
rect 31760 38344 31812 38350
rect 31760 38286 31812 38292
rect 30932 37868 30984 37874
rect 30932 37810 30984 37816
rect 30944 37466 30972 37810
rect 31772 37806 31800 38286
rect 31760 37800 31812 37806
rect 31760 37742 31812 37748
rect 30932 37460 30984 37466
rect 30932 37402 30984 37408
rect 31772 37262 31800 37742
rect 31760 37256 31812 37262
rect 31760 37198 31812 37204
rect 30932 36780 30984 36786
rect 30932 36722 30984 36728
rect 30944 36378 30972 36722
rect 31772 36718 31800 37198
rect 31760 36712 31812 36718
rect 31760 36654 31812 36660
rect 31772 36378 31800 36654
rect 30932 36372 30984 36378
rect 30932 36314 30984 36320
rect 31760 36372 31812 36378
rect 31760 36314 31812 36320
rect 31024 36100 31076 36106
rect 31024 36042 31076 36048
rect 31036 35290 31064 36042
rect 31772 35834 31800 36314
rect 32324 36106 32352 40394
rect 32416 39642 32444 41482
rect 32496 41064 32548 41070
rect 32496 41006 32548 41012
rect 32508 40118 32536 41006
rect 32968 40458 32996 43658
rect 34072 42566 34100 44746
rect 34152 43648 34204 43654
rect 34152 43590 34204 43596
rect 34164 42702 34192 43590
rect 34808 43450 34836 45426
rect 35348 45280 35400 45286
rect 35348 45222 35400 45228
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 35360 43450 35388 45222
rect 35440 44396 35492 44402
rect 35440 44338 35492 44344
rect 35452 43994 35480 44338
rect 36360 44192 36412 44198
rect 36360 44134 36412 44140
rect 35440 43988 35492 43994
rect 35440 43930 35492 43936
rect 34796 43444 34848 43450
rect 34796 43386 34848 43392
rect 35348 43444 35400 43450
rect 35348 43386 35400 43392
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 36372 42702 36400 44134
rect 34152 42696 34204 42702
rect 34152 42638 34204 42644
rect 36360 42696 36412 42702
rect 36360 42638 36412 42644
rect 34704 42628 34756 42634
rect 34704 42570 34756 42576
rect 34060 42560 34112 42566
rect 34060 42502 34112 42508
rect 34244 42220 34296 42226
rect 34244 42162 34296 42168
rect 34060 41132 34112 41138
rect 34060 41074 34112 41080
rect 32956 40452 33008 40458
rect 32956 40394 33008 40400
rect 32496 40112 32548 40118
rect 32496 40054 32548 40060
rect 32772 40044 32824 40050
rect 32772 39986 32824 39992
rect 32404 39636 32456 39642
rect 32404 39578 32456 39584
rect 32784 39506 32812 39986
rect 34072 39642 34100 41074
rect 34152 39840 34204 39846
rect 34152 39782 34204 39788
rect 34060 39636 34112 39642
rect 34060 39578 34112 39584
rect 32772 39500 32824 39506
rect 32772 39442 32824 39448
rect 32784 39370 32812 39442
rect 34164 39438 34192 39782
rect 34152 39432 34204 39438
rect 34152 39374 34204 39380
rect 32772 39364 32824 39370
rect 32772 39306 32824 39312
rect 32784 38962 32812 39306
rect 34256 39098 34284 42162
rect 34716 42158 34744 42570
rect 36556 42566 36584 45426
rect 37924 45416 37976 45422
rect 37924 45358 37976 45364
rect 37936 44878 37964 45358
rect 37924 44872 37976 44878
rect 37924 44814 37976 44820
rect 36728 44736 36780 44742
rect 36728 44678 36780 44684
rect 36636 44396 36688 44402
rect 36636 44338 36688 44344
rect 36648 43178 36676 44338
rect 36740 43382 36768 44678
rect 37936 44334 37964 44814
rect 38016 44804 38068 44810
rect 38016 44746 38068 44752
rect 39120 44804 39172 44810
rect 39120 44746 39172 44752
rect 37924 44328 37976 44334
rect 37924 44270 37976 44276
rect 37936 43790 37964 44270
rect 37372 43784 37424 43790
rect 37372 43726 37424 43732
rect 37924 43784 37976 43790
rect 37924 43726 37976 43732
rect 36728 43376 36780 43382
rect 36728 43318 36780 43324
rect 37384 43246 37412 43726
rect 38028 43450 38056 44746
rect 38016 43444 38068 43450
rect 38016 43386 38068 43392
rect 37372 43240 37424 43246
rect 37372 43182 37424 43188
rect 36636 43172 36688 43178
rect 36636 43114 36688 43120
rect 37384 42702 37412 43182
rect 37372 42696 37424 42702
rect 37372 42638 37424 42644
rect 37832 42696 37884 42702
rect 37832 42638 37884 42644
rect 36544 42560 36596 42566
rect 36544 42502 36596 42508
rect 37844 42226 37872 42638
rect 39132 42566 39160 44746
rect 39224 43994 39252 45426
rect 39396 45280 39448 45286
rect 39396 45222 39448 45228
rect 39304 44736 39356 44742
rect 39304 44678 39356 44684
rect 39212 43988 39264 43994
rect 39212 43930 39264 43936
rect 39316 43790 39344 44678
rect 39304 43784 39356 43790
rect 39304 43726 39356 43732
rect 39212 43716 39264 43722
rect 39212 43658 39264 43664
rect 39224 43314 39252 43658
rect 39408 43382 39436 45222
rect 40408 44872 40460 44878
rect 40408 44814 40460 44820
rect 40420 44334 40448 44814
rect 40408 44328 40460 44334
rect 40408 44270 40460 44276
rect 40040 44192 40092 44198
rect 40040 44134 40092 44140
rect 39396 43376 39448 43382
rect 39396 43318 39448 43324
rect 39212 43308 39264 43314
rect 39212 43250 39264 43256
rect 40052 42702 40080 44134
rect 40316 43308 40368 43314
rect 40316 43250 40368 43256
rect 40040 42696 40092 42702
rect 40040 42638 40092 42644
rect 39120 42560 39172 42566
rect 39120 42502 39172 42508
rect 40040 42560 40092 42566
rect 40040 42502 40092 42508
rect 40052 42242 40080 42502
rect 37832 42220 37884 42226
rect 37832 42162 37884 42168
rect 39960 42214 40080 42242
rect 40224 42220 40276 42226
rect 34704 42152 34756 42158
rect 34704 42094 34756 42100
rect 34716 41682 34744 42094
rect 36084 42016 36136 42022
rect 36084 41958 36136 41964
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34704 41676 34756 41682
rect 34704 41618 34756 41624
rect 35348 41676 35400 41682
rect 35348 41618 35400 41624
rect 35360 41138 35388 41618
rect 35348 41132 35400 41138
rect 35348 41074 35400 41080
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 35992 40520 36044 40526
rect 35992 40462 36044 40468
rect 34336 40452 34388 40458
rect 34336 40394 34388 40400
rect 34348 40118 34376 40394
rect 36004 40118 36032 40462
rect 34336 40112 34388 40118
rect 34336 40054 34388 40060
rect 35992 40112 36044 40118
rect 35992 40054 36044 40060
rect 34348 39506 34376 40054
rect 36096 39846 36124 41958
rect 37844 41614 37872 42162
rect 37832 41608 37884 41614
rect 37832 41550 37884 41556
rect 36544 41540 36596 41546
rect 36544 41482 36596 41488
rect 36268 41472 36320 41478
rect 36268 41414 36320 41420
rect 36084 39840 36136 39846
rect 36084 39782 36136 39788
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34336 39500 34388 39506
rect 34336 39442 34388 39448
rect 34244 39092 34296 39098
rect 34244 39034 34296 39040
rect 36280 39030 36308 41414
rect 36556 41274 36584 41482
rect 37740 41472 37792 41478
rect 37740 41414 37792 41420
rect 36544 41268 36596 41274
rect 36544 41210 36596 41216
rect 36728 41132 36780 41138
rect 36728 41074 36780 41080
rect 36740 40186 36768 41074
rect 37752 40526 37780 41414
rect 37740 40520 37792 40526
rect 37740 40462 37792 40468
rect 37844 40458 37872 41550
rect 39120 41540 39172 41546
rect 39120 41482 39172 41488
rect 37832 40452 37884 40458
rect 37832 40394 37884 40400
rect 37464 40384 37516 40390
rect 37464 40326 37516 40332
rect 36728 40180 36780 40186
rect 36728 40122 36780 40128
rect 37372 40044 37424 40050
rect 37372 39986 37424 39992
rect 37384 39642 37412 39986
rect 37372 39636 37424 39642
rect 37372 39578 37424 39584
rect 37476 39438 37504 40326
rect 37844 39506 37872 40394
rect 38752 39840 38804 39846
rect 38752 39782 38804 39788
rect 38936 39840 38988 39846
rect 38936 39782 38988 39788
rect 37832 39500 37884 39506
rect 37832 39442 37884 39448
rect 37464 39432 37516 39438
rect 37464 39374 37516 39380
rect 36268 39024 36320 39030
rect 36268 38966 36320 38972
rect 38764 38962 38792 39782
rect 38948 39438 38976 39782
rect 39132 39642 39160 41482
rect 39960 41070 39988 42214
rect 40224 42162 40276 42168
rect 39948 41064 40000 41070
rect 39948 41006 40000 41012
rect 39396 40928 39448 40934
rect 39396 40870 39448 40876
rect 39408 40594 39436 40870
rect 39960 40594 39988 41006
rect 40040 40928 40092 40934
rect 40040 40870 40092 40876
rect 40132 40928 40184 40934
rect 40132 40870 40184 40876
rect 39396 40588 39448 40594
rect 39396 40530 39448 40536
rect 39948 40588 40000 40594
rect 39948 40530 40000 40536
rect 39304 40384 39356 40390
rect 39304 40326 39356 40332
rect 39120 39636 39172 39642
rect 39120 39578 39172 39584
rect 38936 39432 38988 39438
rect 38936 39374 38988 39380
rect 39316 39030 39344 40326
rect 39408 40050 39436 40530
rect 40052 40526 40080 40870
rect 40040 40520 40092 40526
rect 40040 40462 40092 40468
rect 40144 40050 40172 40870
rect 39396 40044 39448 40050
rect 39396 39986 39448 39992
rect 40132 40044 40184 40050
rect 40132 39986 40184 39992
rect 40236 39098 40264 42162
rect 40328 42106 40356 43250
rect 40420 42702 40448 44270
rect 40776 44192 40828 44198
rect 40776 44134 40828 44140
rect 40500 43784 40552 43790
rect 40500 43726 40552 43732
rect 40512 43110 40540 43726
rect 40500 43104 40552 43110
rect 40500 43046 40552 43052
rect 40408 42696 40460 42702
rect 40408 42638 40460 42644
rect 40408 42220 40460 42226
rect 40408 42162 40460 42168
rect 40420 42106 40448 42162
rect 40328 42078 40448 42106
rect 40316 42016 40368 42022
rect 40316 41958 40368 41964
rect 40328 39846 40356 41958
rect 40316 39840 40368 39846
rect 40316 39782 40368 39788
rect 40420 39642 40448 42078
rect 40512 41614 40540 43046
rect 40788 42702 40816 44134
rect 40776 42696 40828 42702
rect 40776 42638 40828 42644
rect 40500 41608 40552 41614
rect 40500 41550 40552 41556
rect 40592 41132 40644 41138
rect 40592 41074 40644 41080
rect 40604 40186 40632 41074
rect 40592 40180 40644 40186
rect 40592 40122 40644 40128
rect 40408 39636 40460 39642
rect 40408 39578 40460 39584
rect 40316 39432 40368 39438
rect 40316 39374 40368 39380
rect 40224 39092 40276 39098
rect 40224 39034 40276 39040
rect 39304 39024 39356 39030
rect 39304 38966 39356 38972
rect 32772 38956 32824 38962
rect 32772 38898 32824 38904
rect 36084 38956 36136 38962
rect 36084 38898 36136 38904
rect 38752 38956 38804 38962
rect 38752 38898 38804 38904
rect 34704 38888 34756 38894
rect 34704 38830 34756 38836
rect 34716 38350 34744 38830
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 36096 38554 36124 38898
rect 36636 38752 36688 38758
rect 36636 38694 36688 38700
rect 36084 38548 36136 38554
rect 36084 38490 36136 38496
rect 34704 38344 34756 38350
rect 34704 38286 34756 38292
rect 33508 38276 33560 38282
rect 33508 38218 33560 38224
rect 33520 38010 33548 38218
rect 33508 38004 33560 38010
rect 33508 37946 33560 37952
rect 34716 37942 34744 38286
rect 35348 38276 35400 38282
rect 35348 38218 35400 38224
rect 34796 38208 34848 38214
rect 34796 38150 34848 38156
rect 34704 37936 34756 37942
rect 34704 37878 34756 37884
rect 33140 37868 33192 37874
rect 33140 37810 33192 37816
rect 33152 37466 33180 37810
rect 33140 37460 33192 37466
rect 33140 37402 33192 37408
rect 34716 37330 34744 37878
rect 34704 37324 34756 37330
rect 34704 37266 34756 37272
rect 34808 37262 34836 38150
rect 35360 38010 35388 38218
rect 35348 38004 35400 38010
rect 35348 37946 35400 37952
rect 35348 37868 35400 37874
rect 35348 37810 35400 37816
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34796 37256 34848 37262
rect 34796 37198 34848 37204
rect 33508 37188 33560 37194
rect 33508 37130 33560 37136
rect 33520 36922 33548 37130
rect 35360 37126 35388 37810
rect 36648 37262 36676 38694
rect 38764 38350 38792 38898
rect 38752 38344 38804 38350
rect 38752 38286 38804 38292
rect 37556 38276 37608 38282
rect 37556 38218 37608 38224
rect 37568 37466 37596 38218
rect 37924 38208 37976 38214
rect 37924 38150 37976 38156
rect 37556 37460 37608 37466
rect 37556 37402 37608 37408
rect 35440 37256 35492 37262
rect 35440 37198 35492 37204
rect 36636 37256 36688 37262
rect 36636 37198 36688 37204
rect 35348 37120 35400 37126
rect 35348 37062 35400 37068
rect 33508 36916 33560 36922
rect 33508 36858 33560 36864
rect 35452 36786 35480 37198
rect 37936 36854 37964 38150
rect 38764 37942 38792 38286
rect 38752 37936 38804 37942
rect 38752 37878 38804 37884
rect 38660 37868 38712 37874
rect 38660 37810 38712 37816
rect 39120 37868 39172 37874
rect 39120 37810 39172 37816
rect 39396 37868 39448 37874
rect 39396 37810 39448 37816
rect 38672 36922 38700 37810
rect 38752 37664 38804 37670
rect 38752 37606 38804 37612
rect 38660 36916 38712 36922
rect 38660 36858 38712 36864
rect 37924 36848 37976 36854
rect 37924 36790 37976 36796
rect 33508 36780 33560 36786
rect 33508 36722 33560 36728
rect 35440 36780 35492 36786
rect 35440 36722 35492 36728
rect 38660 36780 38712 36786
rect 38660 36722 38712 36728
rect 32312 36100 32364 36106
rect 32312 36042 32364 36048
rect 33520 35834 33548 36722
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 35452 36174 35480 36722
rect 36728 36576 36780 36582
rect 36728 36518 36780 36524
rect 34612 36168 34664 36174
rect 34612 36110 34664 36116
rect 35440 36168 35492 36174
rect 35440 36110 35492 36116
rect 31760 35828 31812 35834
rect 31760 35770 31812 35776
rect 33508 35828 33560 35834
rect 33508 35770 33560 35776
rect 31772 35290 31800 35770
rect 34624 35630 34652 36110
rect 36084 36100 36136 36106
rect 36084 36042 36136 36048
rect 35992 36032 36044 36038
rect 35992 35974 36044 35980
rect 34612 35624 34664 35630
rect 34612 35566 34664 35572
rect 31024 35284 31076 35290
rect 31024 35226 31076 35232
rect 31760 35284 31812 35290
rect 31760 35226 31812 35232
rect 31772 34610 31800 35226
rect 31852 35012 31904 35018
rect 31852 34954 31904 34960
rect 31760 34604 31812 34610
rect 31760 34546 31812 34552
rect 31864 34202 31892 34954
rect 32128 34604 32180 34610
rect 32128 34546 32180 34552
rect 31852 34196 31904 34202
rect 31852 34138 31904 34144
rect 31668 33992 31720 33998
rect 31668 33934 31720 33940
rect 31680 33318 31708 33934
rect 31760 33516 31812 33522
rect 31760 33458 31812 33464
rect 31208 33312 31260 33318
rect 31208 33254 31260 33260
rect 31668 33312 31720 33318
rect 31668 33254 31720 33260
rect 31220 32910 31248 33254
rect 31208 32904 31260 32910
rect 31208 32846 31260 32852
rect 31300 32768 31352 32774
rect 31300 32710 31352 32716
rect 31312 32502 31340 32710
rect 31300 32496 31352 32502
rect 31300 32438 31352 32444
rect 31680 32434 31708 33254
rect 31772 32570 31800 33458
rect 32140 33454 32168 34546
rect 34624 34542 34652 35566
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 36004 35018 36032 35974
rect 36096 35834 36124 36042
rect 36084 35828 36136 35834
rect 36084 35770 36136 35776
rect 36740 35766 36768 36518
rect 38672 36378 38700 36722
rect 38660 36372 38712 36378
rect 38660 36314 38712 36320
rect 38764 36174 38792 37606
rect 39132 36718 39160 37810
rect 38844 36712 38896 36718
rect 38844 36654 38896 36660
rect 39120 36712 39172 36718
rect 39120 36654 39172 36660
rect 38752 36168 38804 36174
rect 38752 36110 38804 36116
rect 37372 36032 37424 36038
rect 37372 35974 37424 35980
rect 36728 35760 36780 35766
rect 36728 35702 36780 35708
rect 36360 35692 36412 35698
rect 36360 35634 36412 35640
rect 35992 35012 36044 35018
rect 35992 34954 36044 34960
rect 36372 34746 36400 35634
rect 36360 34740 36412 34746
rect 36360 34682 36412 34688
rect 37384 34678 37412 35974
rect 37740 35624 37792 35630
rect 37740 35566 37792 35572
rect 37752 35154 37780 35566
rect 37740 35148 37792 35154
rect 37740 35090 37792 35096
rect 37752 34678 37780 35090
rect 38856 34746 38884 36654
rect 39132 36242 39160 36654
rect 39120 36236 39172 36242
rect 39120 36178 39172 36184
rect 39408 35834 39436 37810
rect 39488 36576 39540 36582
rect 39488 36518 39540 36524
rect 39396 35828 39448 35834
rect 39396 35770 39448 35776
rect 39500 35766 39528 36518
rect 39948 36168 40000 36174
rect 39948 36110 40000 36116
rect 39488 35760 39540 35766
rect 39488 35702 39540 35708
rect 39856 35624 39908 35630
rect 39856 35566 39908 35572
rect 38844 34740 38896 34746
rect 38844 34682 38896 34688
rect 39120 34740 39172 34746
rect 39120 34682 39172 34688
rect 37372 34672 37424 34678
rect 37372 34614 37424 34620
rect 37740 34672 37792 34678
rect 37740 34614 37792 34620
rect 34704 34604 34756 34610
rect 34704 34546 34756 34552
rect 36084 34604 36136 34610
rect 36084 34546 36136 34552
rect 34612 34536 34664 34542
rect 34612 34478 34664 34484
rect 34624 33998 34652 34478
rect 34612 33992 34664 33998
rect 34612 33934 34664 33940
rect 33508 33924 33560 33930
rect 33508 33866 33560 33872
rect 33048 33856 33100 33862
rect 33048 33798 33100 33804
rect 32128 33448 32180 33454
rect 32128 33390 32180 33396
rect 33060 32910 33088 33798
rect 33520 33658 33548 33866
rect 33508 33652 33560 33658
rect 33508 33594 33560 33600
rect 34624 33538 34652 33934
rect 34716 33658 34744 34546
rect 34796 34400 34848 34406
rect 34796 34342 34848 34348
rect 34808 33998 34836 34342
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 36096 34202 36124 34546
rect 37924 34400 37976 34406
rect 37924 34342 37976 34348
rect 36084 34196 36136 34202
rect 36084 34138 36136 34144
rect 37936 33998 37964 34342
rect 39132 33998 39160 34682
rect 39868 34406 39896 35566
rect 39960 35154 39988 36110
rect 40328 35894 40356 39374
rect 40420 37262 40448 39578
rect 40972 39438 41000 51954
rect 41144 51332 41196 51338
rect 41144 51274 41196 51280
rect 41156 49434 41184 51274
rect 41788 51264 41840 51270
rect 41788 51206 41840 51212
rect 41696 50856 41748 50862
rect 41696 50798 41748 50804
rect 41708 50318 41736 50798
rect 41800 50318 41828 51206
rect 41696 50312 41748 50318
rect 41696 50254 41748 50260
rect 41788 50312 41840 50318
rect 41788 50254 41840 50260
rect 41236 50176 41288 50182
rect 41236 50118 41288 50124
rect 41420 50176 41472 50182
rect 41420 50118 41472 50124
rect 41248 49910 41276 50118
rect 41236 49904 41288 49910
rect 41236 49846 41288 49852
rect 41144 49428 41196 49434
rect 41144 49370 41196 49376
rect 41432 48822 41460 50118
rect 41708 49230 41736 50254
rect 43088 49910 43116 52090
rect 44468 52086 44496 53382
rect 44560 52154 44588 54538
rect 45296 54262 45324 54606
rect 45284 54256 45336 54262
rect 45284 54198 45336 54204
rect 44824 54188 44876 54194
rect 44824 54130 44876 54136
rect 44836 53242 44864 54130
rect 45296 54126 45324 54198
rect 45284 54120 45336 54126
rect 45284 54062 45336 54068
rect 45192 53984 45244 53990
rect 45192 53926 45244 53932
rect 44824 53236 44876 53242
rect 44824 53178 44876 53184
rect 45204 52494 45232 53926
rect 45296 53582 45324 54062
rect 47032 53984 47084 53990
rect 47032 53926 47084 53932
rect 47044 53582 47072 53926
rect 47136 53582 47164 58482
rect 47320 58138 47348 58890
rect 47768 58880 47820 58886
rect 47768 58822 47820 58828
rect 48320 58880 48372 58886
rect 48320 58822 48372 58828
rect 47780 58614 47808 58822
rect 47768 58608 47820 58614
rect 47768 58550 47820 58556
rect 47308 58132 47360 58138
rect 47308 58074 47360 58080
rect 48332 55758 48360 58822
rect 48516 56846 48544 59366
rect 48792 57934 48820 59910
rect 48976 59634 49004 60046
rect 49332 60036 49384 60042
rect 49332 59978 49384 59984
rect 50620 60036 50672 60042
rect 50620 59978 50672 59984
rect 48964 59628 49016 59634
rect 48964 59570 49016 59576
rect 48976 59022 49004 59570
rect 48964 59016 49016 59022
rect 48964 58958 49016 58964
rect 48976 58342 49004 58958
rect 48964 58336 49016 58342
rect 48964 58278 49016 58284
rect 48976 58138 49004 58278
rect 48964 58132 49016 58138
rect 48964 58074 49016 58080
rect 48780 57928 48832 57934
rect 48780 57870 48832 57876
rect 48976 57390 49004 58074
rect 48964 57384 49016 57390
rect 48964 57326 49016 57332
rect 48504 56840 48556 56846
rect 48504 56782 48556 56788
rect 48976 56778 49004 57326
rect 48964 56772 49016 56778
rect 48964 56714 49016 56720
rect 48976 56370 49004 56714
rect 48964 56364 49016 56370
rect 48964 56306 49016 56312
rect 49344 55962 49372 59978
rect 50294 59868 50602 59888
rect 50294 59866 50300 59868
rect 50356 59866 50380 59868
rect 50436 59866 50460 59868
rect 50516 59866 50540 59868
rect 50596 59866 50602 59868
rect 50356 59814 50358 59866
rect 50538 59814 50540 59866
rect 50294 59812 50300 59814
rect 50356 59812 50380 59814
rect 50436 59812 50460 59814
rect 50516 59812 50540 59814
rect 50596 59812 50602 59814
rect 50294 59792 50602 59812
rect 49516 59628 49568 59634
rect 49516 59570 49568 59576
rect 49424 58948 49476 58954
rect 49424 58890 49476 58896
rect 49436 57050 49464 58890
rect 49528 57594 49556 59570
rect 50294 58780 50602 58800
rect 50294 58778 50300 58780
rect 50356 58778 50380 58780
rect 50436 58778 50460 58780
rect 50516 58778 50540 58780
rect 50596 58778 50602 58780
rect 50356 58726 50358 58778
rect 50538 58726 50540 58778
rect 50294 58724 50300 58726
rect 50356 58724 50380 58726
rect 50436 58724 50460 58726
rect 50516 58724 50540 58726
rect 50596 58724 50602 58726
rect 50294 58704 50602 58724
rect 49608 57792 49660 57798
rect 49608 57734 49660 57740
rect 49516 57588 49568 57594
rect 49516 57530 49568 57536
rect 49424 57044 49476 57050
rect 49424 56986 49476 56992
rect 49620 56438 49648 57734
rect 50294 57692 50602 57712
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57616 50602 57636
rect 50160 57384 50212 57390
rect 50160 57326 50212 57332
rect 50172 56914 50200 57326
rect 50160 56908 50212 56914
rect 50160 56850 50212 56856
rect 49608 56432 49660 56438
rect 49608 56374 49660 56380
rect 49332 55956 49384 55962
rect 49332 55898 49384 55904
rect 50172 55758 50200 56850
rect 50294 56604 50602 56624
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56528 50602 56548
rect 50632 56506 50660 59978
rect 50816 59566 50844 60046
rect 51540 59968 51592 59974
rect 51540 59910 51592 59916
rect 53196 59968 53248 59974
rect 53196 59910 53248 59916
rect 50804 59560 50856 59566
rect 50804 59502 50856 59508
rect 50816 59022 50844 59502
rect 51080 59424 51132 59430
rect 51080 59366 51132 59372
rect 50804 59016 50856 59022
rect 50804 58958 50856 58964
rect 50816 58478 50844 58958
rect 50804 58472 50856 58478
rect 50804 58414 50856 58420
rect 50816 57934 50844 58414
rect 50804 57928 50856 57934
rect 50804 57870 50856 57876
rect 50816 57390 50844 57870
rect 51092 57866 51120 59366
rect 51080 57860 51132 57866
rect 51080 57802 51132 57808
rect 51552 57458 51580 59910
rect 51908 59628 51960 59634
rect 51908 59570 51960 59576
rect 51540 57452 51592 57458
rect 51540 57394 51592 57400
rect 50804 57384 50856 57390
rect 50804 57326 50856 57332
rect 50620 56500 50672 56506
rect 50620 56442 50672 56448
rect 51920 56234 51948 59570
rect 53208 59022 53236 59910
rect 53380 59560 53432 59566
rect 53380 59502 53432 59508
rect 53392 59022 53420 59502
rect 53196 59016 53248 59022
rect 53196 58958 53248 58964
rect 53380 59016 53432 59022
rect 53380 58958 53432 58964
rect 52552 58880 52604 58886
rect 52552 58822 52604 58828
rect 52184 58336 52236 58342
rect 52184 58278 52236 58284
rect 52196 57526 52224 58278
rect 52184 57520 52236 57526
rect 52184 57462 52236 57468
rect 52184 57248 52236 57254
rect 52184 57190 52236 57196
rect 52196 56438 52224 57190
rect 52564 56846 52592 58822
rect 53104 58608 53156 58614
rect 53104 58550 53156 58556
rect 52920 58540 52972 58546
rect 52920 58482 52972 58488
rect 52932 58138 52960 58482
rect 52920 58132 52972 58138
rect 52920 58074 52972 58080
rect 52828 57860 52880 57866
rect 52828 57802 52880 57808
rect 52840 57050 52868 57802
rect 53116 57526 53144 58550
rect 53392 57934 53420 58958
rect 54128 58546 54156 60046
rect 54944 60036 54996 60042
rect 54944 59978 54996 59984
rect 58440 60036 58492 60042
rect 58440 59978 58492 59984
rect 54956 59770 54984 59978
rect 54944 59764 54996 59770
rect 54944 59706 54996 59712
rect 55404 59696 55456 59702
rect 55404 59638 55456 59644
rect 54760 59628 54812 59634
rect 54760 59570 54812 59576
rect 54852 59628 54904 59634
rect 54852 59570 54904 59576
rect 54772 59226 54800 59570
rect 54760 59220 54812 59226
rect 54760 59162 54812 59168
rect 54760 58948 54812 58954
rect 54760 58890 54812 58896
rect 54116 58540 54168 58546
rect 54116 58482 54168 58488
rect 54392 58336 54444 58342
rect 54392 58278 54444 58284
rect 54404 57934 54432 58278
rect 54772 58138 54800 58890
rect 54760 58132 54812 58138
rect 54760 58074 54812 58080
rect 53380 57928 53432 57934
rect 53380 57870 53432 57876
rect 54392 57928 54444 57934
rect 54392 57870 54444 57876
rect 53392 57594 53420 57870
rect 53380 57588 53432 57594
rect 53380 57530 53432 57536
rect 53104 57520 53156 57526
rect 53104 57462 53156 57468
rect 52828 57044 52880 57050
rect 52828 56986 52880 56992
rect 53392 56846 53420 57530
rect 54864 57050 54892 59570
rect 55416 59022 55444 59638
rect 55864 59560 55916 59566
rect 55864 59502 55916 59508
rect 55404 59016 55456 59022
rect 55404 58958 55456 58964
rect 55876 58546 55904 59502
rect 55956 59424 56008 59430
rect 55956 59366 56008 59372
rect 55968 58614 55996 59366
rect 58452 59226 58480 59978
rect 57520 59220 57572 59226
rect 57520 59162 57572 59168
rect 58440 59220 58492 59226
rect 58440 59162 58492 59168
rect 57060 59016 57112 59022
rect 57060 58958 57112 58964
rect 56784 58948 56836 58954
rect 56784 58890 56836 58896
rect 55956 58608 56008 58614
rect 55956 58550 56008 58556
rect 55220 58540 55272 58546
rect 55220 58482 55272 58488
rect 55864 58540 55916 58546
rect 55864 58482 55916 58488
rect 55232 57934 55260 58482
rect 55220 57928 55272 57934
rect 55220 57870 55272 57876
rect 55232 57458 55260 57870
rect 56600 57792 56652 57798
rect 56600 57734 56652 57740
rect 56140 57520 56192 57526
rect 56140 57462 56192 57468
rect 55220 57452 55272 57458
rect 55220 57394 55272 57400
rect 54852 57044 54904 57050
rect 54852 56986 54904 56992
rect 55232 56914 55260 57394
rect 55220 56908 55272 56914
rect 55220 56850 55272 56856
rect 52552 56840 52604 56846
rect 52552 56782 52604 56788
rect 53380 56840 53432 56846
rect 53380 56782 53432 56788
rect 52644 56772 52696 56778
rect 52644 56714 52696 56720
rect 52184 56432 52236 56438
rect 52184 56374 52236 56380
rect 51908 56228 51960 56234
rect 51908 56170 51960 56176
rect 48320 55752 48372 55758
rect 48320 55694 48372 55700
rect 50160 55752 50212 55758
rect 50160 55694 50212 55700
rect 49700 55412 49752 55418
rect 49700 55354 49752 55360
rect 49056 55276 49108 55282
rect 49056 55218 49108 55224
rect 47584 55208 47636 55214
rect 47584 55150 47636 55156
rect 47596 54670 47624 55150
rect 49068 54874 49096 55218
rect 49056 54868 49108 54874
rect 49056 54810 49108 54816
rect 47584 54664 47636 54670
rect 47584 54606 47636 54612
rect 47216 54528 47268 54534
rect 47216 54470 47268 54476
rect 47228 54262 47256 54470
rect 47216 54256 47268 54262
rect 47216 54198 47268 54204
rect 47596 54126 47624 54606
rect 48964 54596 49016 54602
rect 48964 54538 49016 54544
rect 48976 54330 49004 54538
rect 49712 54330 49740 55354
rect 50172 54670 50200 55694
rect 51172 55684 51224 55690
rect 51172 55626 51224 55632
rect 50294 55516 50602 55536
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55440 50602 55460
rect 50896 55276 50948 55282
rect 50896 55218 50948 55224
rect 50160 54664 50212 54670
rect 50160 54606 50212 54612
rect 48964 54324 49016 54330
rect 48964 54266 49016 54272
rect 49700 54324 49752 54330
rect 49700 54266 49752 54272
rect 50172 54194 50200 54606
rect 50294 54428 50602 54448
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54352 50602 54372
rect 50908 54330 50936 55218
rect 51184 54874 51212 55626
rect 51540 55616 51592 55622
rect 51540 55558 51592 55564
rect 51552 55350 51580 55558
rect 52552 55412 52604 55418
rect 52552 55354 52604 55360
rect 51540 55344 51592 55350
rect 51540 55286 51592 55292
rect 51264 55072 51316 55078
rect 51264 55014 51316 55020
rect 51172 54868 51224 54874
rect 51172 54810 51224 54816
rect 51276 54670 51304 55014
rect 52564 54670 52592 55354
rect 52656 55282 52684 56714
rect 55232 56522 55260 56850
rect 55680 56772 55732 56778
rect 55680 56714 55732 56720
rect 55140 56494 55260 56522
rect 55692 56506 55720 56714
rect 55680 56500 55732 56506
rect 55140 56438 55168 56494
rect 55680 56442 55732 56448
rect 55128 56432 55180 56438
rect 55128 56374 55180 56380
rect 55956 56364 56008 56370
rect 55956 56306 56008 56312
rect 53380 56296 53432 56302
rect 53380 56238 53432 56244
rect 53392 55758 53420 56238
rect 52736 55752 52788 55758
rect 52736 55694 52788 55700
rect 53380 55752 53432 55758
rect 53380 55694 53432 55700
rect 52644 55276 52696 55282
rect 52644 55218 52696 55224
rect 51264 54664 51316 54670
rect 51264 54606 51316 54612
rect 52552 54664 52604 54670
rect 52552 54606 52604 54612
rect 52748 54602 52776 55694
rect 55968 55418 55996 56306
rect 56152 55690 56180 57462
rect 56612 55758 56640 57734
rect 56692 57452 56744 57458
rect 56692 57394 56744 57400
rect 56704 57050 56732 57394
rect 56692 57044 56744 57050
rect 56692 56986 56744 56992
rect 56796 55962 56824 58890
rect 57072 58546 57100 58958
rect 57060 58540 57112 58546
rect 57060 58482 57112 58488
rect 56876 58336 56928 58342
rect 56876 58278 56928 58284
rect 56888 56846 56916 58278
rect 57072 57934 57100 58482
rect 57060 57928 57112 57934
rect 57060 57870 57112 57876
rect 57072 56846 57100 57870
rect 57244 57248 57296 57254
rect 57244 57190 57296 57196
rect 57256 56846 57284 57190
rect 56876 56840 56928 56846
rect 56876 56782 56928 56788
rect 57060 56840 57112 56846
rect 57060 56782 57112 56788
rect 57244 56840 57296 56846
rect 57244 56782 57296 56788
rect 56784 55956 56836 55962
rect 56784 55898 56836 55904
rect 56600 55752 56652 55758
rect 56600 55694 56652 55700
rect 56140 55684 56192 55690
rect 56140 55626 56192 55632
rect 56152 55570 56180 55626
rect 57072 55622 57100 56782
rect 56060 55542 56180 55570
rect 57060 55616 57112 55622
rect 57060 55558 57112 55564
rect 55956 55412 56008 55418
rect 55956 55354 56008 55360
rect 55496 55072 55548 55078
rect 55496 55014 55548 55020
rect 52736 54596 52788 54602
rect 52736 54538 52788 54544
rect 52552 54528 52604 54534
rect 52552 54470 52604 54476
rect 50896 54324 50948 54330
rect 50896 54266 50948 54272
rect 48964 54188 49016 54194
rect 48964 54130 49016 54136
rect 50160 54188 50212 54194
rect 50160 54130 50212 54136
rect 52460 54188 52512 54194
rect 52460 54130 52512 54136
rect 47584 54120 47636 54126
rect 47584 54062 47636 54068
rect 45284 53576 45336 53582
rect 45284 53518 45336 53524
rect 47032 53576 47084 53582
rect 47032 53518 47084 53524
rect 47124 53576 47176 53582
rect 47124 53518 47176 53524
rect 45296 53038 45324 53518
rect 46664 53440 46716 53446
rect 46664 53382 46716 53388
rect 46676 53174 46704 53382
rect 46664 53168 46716 53174
rect 46664 53110 46716 53116
rect 45284 53032 45336 53038
rect 45284 52974 45336 52980
rect 45468 52896 45520 52902
rect 45468 52838 45520 52844
rect 45480 52494 45508 52838
rect 45192 52488 45244 52494
rect 45192 52430 45244 52436
rect 45468 52488 45520 52494
rect 45468 52430 45520 52436
rect 44548 52148 44600 52154
rect 44548 52090 44600 52096
rect 44456 52080 44508 52086
rect 44456 52022 44508 52028
rect 43168 51944 43220 51950
rect 43168 51886 43220 51892
rect 43180 50998 43208 51886
rect 45480 51490 45508 52430
rect 47136 52154 47164 53518
rect 47596 53446 47624 54062
rect 47584 53440 47636 53446
rect 47584 53382 47636 53388
rect 47596 53038 47624 53382
rect 48976 53242 49004 54130
rect 50172 53650 50200 54130
rect 52472 53786 52500 54130
rect 52460 53780 52512 53786
rect 52460 53722 52512 53728
rect 50160 53644 50212 53650
rect 50160 53586 50212 53592
rect 52564 53582 52592 54470
rect 52748 54126 52776 54538
rect 55404 54188 55456 54194
rect 55404 54130 55456 54136
rect 52736 54120 52788 54126
rect 52736 54062 52788 54068
rect 52920 53984 52972 53990
rect 52920 53926 52972 53932
rect 54116 53984 54168 53990
rect 54116 53926 54168 53932
rect 52932 53582 52960 53926
rect 54128 53582 54156 53926
rect 52552 53576 52604 53582
rect 52552 53518 52604 53524
rect 52920 53576 52972 53582
rect 52920 53518 52972 53524
rect 54116 53576 54168 53582
rect 54116 53518 54168 53524
rect 51356 53440 51408 53446
rect 51356 53382 51408 53388
rect 50294 53340 50602 53360
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53264 50602 53284
rect 48964 53236 49016 53242
rect 48964 53178 49016 53184
rect 48320 53100 48372 53106
rect 48320 53042 48372 53048
rect 47584 53032 47636 53038
rect 47584 52974 47636 52980
rect 47596 52426 47624 52974
rect 48332 52698 48360 53042
rect 48320 52692 48372 52698
rect 48320 52634 48372 52640
rect 51368 52494 51396 53382
rect 52932 53106 52960 53518
rect 55416 53242 55444 54130
rect 55508 54126 55536 55014
rect 55496 54120 55548 54126
rect 55496 54062 55548 54068
rect 55956 53576 56008 53582
rect 55956 53518 56008 53524
rect 55404 53236 55456 53242
rect 55404 53178 55456 53184
rect 55968 53106 55996 53518
rect 52920 53100 52972 53106
rect 52920 53042 52972 53048
rect 54760 53100 54812 53106
rect 54760 53042 54812 53048
rect 55956 53100 56008 53106
rect 55956 53042 56008 53048
rect 54772 52698 54800 53042
rect 54760 52692 54812 52698
rect 54760 52634 54812 52640
rect 55968 52562 55996 53042
rect 55956 52556 56008 52562
rect 55956 52498 56008 52504
rect 48964 52488 49016 52494
rect 48964 52430 49016 52436
rect 51356 52488 51408 52494
rect 51356 52430 51408 52436
rect 53104 52488 53156 52494
rect 53104 52430 53156 52436
rect 54484 52488 54536 52494
rect 54484 52430 54536 52436
rect 47584 52420 47636 52426
rect 47584 52362 47636 52368
rect 47124 52148 47176 52154
rect 47124 52090 47176 52096
rect 47596 51950 47624 52362
rect 48976 52154 49004 52430
rect 52460 52352 52512 52358
rect 52460 52294 52512 52300
rect 50294 52252 50602 52272
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52176 50602 52196
rect 48964 52148 49016 52154
rect 48964 52090 49016 52096
rect 52472 52086 52500 52294
rect 52460 52080 52512 52086
rect 52460 52022 52512 52028
rect 53116 52018 53144 52430
rect 54496 52154 54524 52430
rect 54484 52148 54536 52154
rect 54484 52090 54536 52096
rect 55968 52018 55996 52498
rect 49056 52012 49108 52018
rect 49056 51954 49108 51960
rect 53104 52012 53156 52018
rect 53104 51954 53156 51960
rect 54300 52012 54352 52018
rect 54300 51954 54352 51960
rect 55956 52012 56008 52018
rect 55956 51954 56008 51960
rect 47584 51944 47636 51950
rect 47584 51886 47636 51892
rect 48780 51944 48832 51950
rect 48780 51886 48832 51892
rect 45480 51474 45600 51490
rect 45480 51468 45612 51474
rect 45480 51462 45560 51468
rect 45560 51410 45612 51416
rect 47596 51406 47624 51886
rect 47584 51400 47636 51406
rect 47584 51342 47636 51348
rect 47216 51264 47268 51270
rect 47216 51206 47268 51212
rect 47228 50998 47256 51206
rect 43168 50992 43220 50998
rect 43168 50934 43220 50940
rect 47216 50992 47268 50998
rect 47216 50934 47268 50940
rect 43720 50924 43772 50930
rect 43720 50866 43772 50872
rect 44272 50924 44324 50930
rect 44272 50866 44324 50872
rect 46388 50924 46440 50930
rect 46388 50866 46440 50872
rect 43076 49904 43128 49910
rect 43076 49846 43128 49852
rect 41696 49224 41748 49230
rect 41696 49166 41748 49172
rect 41420 48816 41472 48822
rect 41420 48758 41472 48764
rect 41708 48754 41736 49166
rect 41788 49156 41840 49162
rect 41788 49098 41840 49104
rect 41800 48890 41828 49098
rect 43076 49088 43128 49094
rect 43076 49030 43128 49036
rect 41788 48884 41840 48890
rect 41788 48826 41840 48832
rect 43088 48822 43116 49030
rect 43076 48816 43128 48822
rect 43076 48758 43128 48764
rect 41696 48748 41748 48754
rect 41696 48690 41748 48696
rect 42432 48748 42484 48754
rect 42432 48690 42484 48696
rect 42444 48210 42472 48690
rect 42984 48544 43036 48550
rect 42984 48486 43036 48492
rect 42432 48204 42484 48210
rect 42432 48146 42484 48152
rect 41144 48068 41196 48074
rect 41144 48010 41196 48016
rect 41156 45354 41184 48010
rect 41788 48000 41840 48006
rect 41788 47942 41840 47948
rect 41328 47592 41380 47598
rect 41328 47534 41380 47540
rect 41340 47054 41368 47534
rect 41800 47054 41828 47942
rect 42444 47666 42472 48146
rect 42996 48142 43024 48486
rect 43732 48278 43760 50866
rect 43812 50720 43864 50726
rect 43812 50662 43864 50668
rect 43824 49910 43852 50662
rect 44284 50318 44312 50866
rect 45652 50720 45704 50726
rect 45652 50662 45704 50668
rect 44272 50312 44324 50318
rect 44272 50254 44324 50260
rect 44284 49978 44312 50254
rect 44272 49972 44324 49978
rect 44272 49914 44324 49920
rect 43812 49904 43864 49910
rect 43812 49846 43864 49852
rect 45008 49768 45060 49774
rect 45008 49710 45060 49716
rect 45020 49230 45048 49710
rect 45664 49230 45692 50662
rect 46296 50244 46348 50250
rect 46296 50186 46348 50192
rect 46308 49434 46336 50186
rect 46296 49428 46348 49434
rect 46296 49370 46348 49376
rect 45008 49224 45060 49230
rect 45008 49166 45060 49172
rect 45652 49224 45704 49230
rect 45652 49166 45704 49172
rect 44456 48748 44508 48754
rect 44456 48690 44508 48696
rect 43720 48272 43772 48278
rect 43720 48214 43772 48220
rect 42984 48136 43036 48142
rect 42984 48078 43036 48084
rect 44468 47802 44496 48690
rect 45020 48686 45048 49166
rect 46400 48890 46428 50866
rect 47596 50862 47624 51342
rect 47768 51332 47820 51338
rect 47768 51274 47820 51280
rect 47584 50856 47636 50862
rect 47584 50798 47636 50804
rect 47596 50318 47624 50798
rect 47780 50522 47808 51274
rect 47768 50516 47820 50522
rect 47768 50458 47820 50464
rect 47584 50312 47636 50318
rect 47584 50254 47636 50260
rect 48792 49842 48820 51886
rect 49068 51610 49096 51954
rect 52184 51808 52236 51814
rect 52184 51750 52236 51756
rect 49056 51604 49108 51610
rect 49056 51546 49108 51552
rect 52196 51406 52224 51750
rect 53116 51490 53144 51954
rect 54312 51610 54340 51954
rect 55968 51610 55996 51954
rect 54300 51604 54352 51610
rect 54300 51546 54352 51552
rect 55956 51604 56008 51610
rect 55956 51546 56008 51552
rect 53024 51462 53144 51490
rect 53024 51406 53052 51462
rect 50620 51400 50672 51406
rect 50620 51342 50672 51348
rect 52184 51400 52236 51406
rect 52184 51342 52236 51348
rect 53012 51400 53064 51406
rect 53012 51342 53064 51348
rect 48964 51332 49016 51338
rect 48964 51274 49016 51280
rect 48976 51066 49004 51274
rect 50294 51164 50602 51184
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51088 50602 51108
rect 48964 51060 49016 51066
rect 48964 51002 49016 51008
rect 50632 50862 50660 51342
rect 52276 51264 52328 51270
rect 52276 51206 52328 51212
rect 52288 50998 52316 51206
rect 55968 50998 55996 51546
rect 56060 51338 56088 55542
rect 56140 55276 56192 55282
rect 56140 55218 56192 55224
rect 56152 54330 56180 55218
rect 57072 55078 57100 55558
rect 57060 55072 57112 55078
rect 57060 55014 57112 55020
rect 57072 54738 57100 55014
rect 57060 54732 57112 54738
rect 57060 54674 57112 54680
rect 57336 54596 57388 54602
rect 57336 54538 57388 54544
rect 56140 54324 56192 54330
rect 56140 54266 56192 54272
rect 57348 53242 57376 54538
rect 57336 53236 57388 53242
rect 57336 53178 57388 53184
rect 57336 52420 57388 52426
rect 57336 52362 57388 52368
rect 57348 52154 57376 52362
rect 57336 52148 57388 52154
rect 57336 52090 57388 52096
rect 57152 52012 57204 52018
rect 57152 51954 57204 51960
rect 56048 51332 56100 51338
rect 56048 51274 56100 51280
rect 52276 50992 52328 50998
rect 52276 50934 52328 50940
rect 55956 50992 56008 50998
rect 55956 50934 56008 50940
rect 50620 50856 50672 50862
rect 50620 50798 50672 50804
rect 50632 50318 50660 50798
rect 52184 50720 52236 50726
rect 52184 50662 52236 50668
rect 52196 50318 52224 50662
rect 55968 50386 55996 50934
rect 55956 50380 56008 50386
rect 55956 50322 56008 50328
rect 50620 50312 50672 50318
rect 50620 50254 50672 50260
rect 52184 50312 52236 50318
rect 52184 50254 52236 50260
rect 50294 50076 50602 50096
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50000 50602 50020
rect 48780 49836 48832 49842
rect 48780 49778 48832 49784
rect 46756 49632 46808 49638
rect 46756 49574 46808 49580
rect 46388 48884 46440 48890
rect 46388 48826 46440 48832
rect 45008 48680 45060 48686
rect 45008 48622 45060 48628
rect 45020 48210 45048 48622
rect 45008 48204 45060 48210
rect 45008 48146 45060 48152
rect 46388 48068 46440 48074
rect 46388 48010 46440 48016
rect 44456 47796 44508 47802
rect 44456 47738 44508 47744
rect 42432 47660 42484 47666
rect 42432 47602 42484 47608
rect 45652 47660 45704 47666
rect 45652 47602 45704 47608
rect 41328 47048 41380 47054
rect 41328 46990 41380 46996
rect 41788 47048 41840 47054
rect 41788 46990 41840 46996
rect 41236 46912 41288 46918
rect 41236 46854 41288 46860
rect 41248 46646 41276 46854
rect 41236 46640 41288 46646
rect 41236 46582 41288 46588
rect 41340 45966 41368 46990
rect 42444 46578 42472 47602
rect 44548 47456 44600 47462
rect 44548 47398 44600 47404
rect 43076 46912 43128 46918
rect 43076 46854 43128 46860
rect 42432 46572 42484 46578
rect 42432 46514 42484 46520
rect 42800 46368 42852 46374
rect 42800 46310 42852 46316
rect 41328 45960 41380 45966
rect 41328 45902 41380 45908
rect 42432 45960 42484 45966
rect 42432 45902 42484 45908
rect 41972 45824 42024 45830
rect 41972 45766 42024 45772
rect 41984 45490 42012 45766
rect 42444 45490 42472 45902
rect 42812 45558 42840 46310
rect 43088 45966 43116 46854
rect 43812 46572 43864 46578
rect 43812 46514 43864 46520
rect 44180 46572 44232 46578
rect 44180 46514 44232 46520
rect 43824 46170 43852 46514
rect 43812 46164 43864 46170
rect 43812 46106 43864 46112
rect 43076 45960 43128 45966
rect 43076 45902 43128 45908
rect 42800 45552 42852 45558
rect 42800 45494 42852 45500
rect 41972 45484 42024 45490
rect 41972 45426 42024 45432
rect 42432 45484 42484 45490
rect 42432 45426 42484 45432
rect 42524 45484 42576 45490
rect 42524 45426 42576 45432
rect 42536 45370 42564 45426
rect 41144 45348 41196 45354
rect 41144 45290 41196 45296
rect 42444 45342 42564 45370
rect 44192 45354 44220 46514
rect 44272 46504 44324 46510
rect 44272 46446 44324 46452
rect 44284 46034 44312 46446
rect 44272 46028 44324 46034
rect 44272 45970 44324 45976
rect 44560 45558 44588 47398
rect 45664 46714 45692 47602
rect 46400 47258 46428 48010
rect 46768 47734 46796 49574
rect 48228 49292 48280 49298
rect 48228 49234 48280 49240
rect 48240 48346 48268 49234
rect 48792 49162 48820 49778
rect 50632 49774 50660 50254
rect 52092 50176 52144 50182
rect 52092 50118 52144 50124
rect 52104 49910 52132 50118
rect 55404 49972 55456 49978
rect 55404 49914 55456 49920
rect 52092 49904 52144 49910
rect 52092 49846 52144 49852
rect 53932 49836 53984 49842
rect 53932 49778 53984 49784
rect 50620 49768 50672 49774
rect 50620 49710 50672 49716
rect 52736 49768 52788 49774
rect 52736 49710 52788 49716
rect 50160 49632 50212 49638
rect 50160 49574 50212 49580
rect 50068 49224 50120 49230
rect 50068 49166 50120 49172
rect 48780 49156 48832 49162
rect 48780 49098 48832 49104
rect 48792 48754 48820 49098
rect 49792 49088 49844 49094
rect 49792 49030 49844 49036
rect 48780 48748 48832 48754
rect 48780 48690 48832 48696
rect 48228 48340 48280 48346
rect 48228 48282 48280 48288
rect 48240 48210 48268 48282
rect 48228 48204 48280 48210
rect 48228 48146 48280 48152
rect 47860 48000 47912 48006
rect 47860 47942 47912 47948
rect 46756 47728 46808 47734
rect 46756 47670 46808 47676
rect 46388 47252 46440 47258
rect 46388 47194 46440 47200
rect 46940 47048 46992 47054
rect 46940 46990 46992 46996
rect 46204 46980 46256 46986
rect 46204 46922 46256 46928
rect 45652 46708 45704 46714
rect 45652 46650 45704 46656
rect 46216 46170 46244 46922
rect 46952 46578 46980 46990
rect 47872 46646 47900 47942
rect 48240 47122 48268 48146
rect 49804 48142 49832 49030
rect 50080 48618 50108 49166
rect 50172 48822 50200 49574
rect 50632 49162 50660 49710
rect 52748 49230 52776 49710
rect 52736 49224 52788 49230
rect 52736 49166 52788 49172
rect 50620 49156 50672 49162
rect 50620 49098 50672 49104
rect 50294 48988 50602 49008
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48912 50602 48932
rect 50160 48816 50212 48822
rect 50160 48758 50212 48764
rect 50068 48612 50120 48618
rect 50068 48554 50120 48560
rect 50068 48272 50120 48278
rect 50068 48214 50120 48220
rect 49792 48136 49844 48142
rect 49792 48078 49844 48084
rect 49700 48068 49752 48074
rect 49700 48010 49752 48016
rect 49608 48000 49660 48006
rect 49608 47942 49660 47948
rect 48228 47116 48280 47122
rect 48228 47058 48280 47064
rect 47860 46640 47912 46646
rect 47860 46582 47912 46588
rect 48240 46578 48268 47058
rect 49620 47054 49648 47942
rect 49712 47258 49740 48010
rect 50080 47802 50108 48214
rect 50294 47900 50602 47920
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47824 50602 47844
rect 50068 47796 50120 47802
rect 50068 47738 50120 47744
rect 49700 47252 49752 47258
rect 49700 47194 49752 47200
rect 49608 47048 49660 47054
rect 49608 46990 49660 46996
rect 46940 46572 46992 46578
rect 46940 46514 46992 46520
rect 48228 46572 48280 46578
rect 48228 46514 48280 46520
rect 46204 46164 46256 46170
rect 46204 46106 46256 46112
rect 46952 45966 46980 46514
rect 48964 46368 49016 46374
rect 48964 46310 49016 46316
rect 48976 45966 49004 46310
rect 50080 46034 50108 47738
rect 50632 47054 50660 49098
rect 52748 48550 52776 49166
rect 53380 49156 53432 49162
rect 53380 49098 53432 49104
rect 53196 48748 53248 48754
rect 53196 48690 53248 48696
rect 52736 48544 52788 48550
rect 52736 48486 52788 48492
rect 52748 48142 52776 48486
rect 52736 48136 52788 48142
rect 52736 48078 52788 48084
rect 50896 48000 50948 48006
rect 50896 47942 50948 47948
rect 50908 47054 50936 47942
rect 52552 47660 52604 47666
rect 52552 47602 52604 47608
rect 50620 47048 50672 47054
rect 50620 46990 50672 46996
rect 50896 47048 50948 47054
rect 50896 46990 50948 46996
rect 50294 46812 50602 46832
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46736 50602 46756
rect 50632 46714 50660 46990
rect 52460 46980 52512 46986
rect 52460 46922 52512 46928
rect 52000 46912 52052 46918
rect 52000 46854 52052 46860
rect 50620 46708 50672 46714
rect 50620 46650 50672 46656
rect 52012 46646 52040 46854
rect 52000 46640 52052 46646
rect 52000 46582 52052 46588
rect 51540 46368 51592 46374
rect 51540 46310 51592 46316
rect 50068 46028 50120 46034
rect 50068 45970 50120 45976
rect 51552 45966 51580 46310
rect 52472 45966 52500 46922
rect 52564 46170 52592 47602
rect 52748 47598 52776 48078
rect 53208 47734 53236 48690
rect 53392 48346 53420 49098
rect 53840 49088 53892 49094
rect 53840 49030 53892 49036
rect 53380 48340 53432 48346
rect 53380 48282 53432 48288
rect 53196 47728 53248 47734
rect 53196 47670 53248 47676
rect 52736 47592 52788 47598
rect 52736 47534 52788 47540
rect 52748 46986 52776 47534
rect 53852 47054 53880 49030
rect 53944 47258 53972 49778
rect 55312 49292 55364 49298
rect 55312 49234 55364 49240
rect 55324 48686 55352 49234
rect 55416 48822 55444 49914
rect 55968 49434 55996 50322
rect 55956 49428 56008 49434
rect 55956 49370 56008 49376
rect 55404 48816 55456 48822
rect 55404 48758 55456 48764
rect 56060 48754 56088 51274
rect 57164 51066 57192 51954
rect 57152 51060 57204 51066
rect 57152 51002 57204 51008
rect 57428 50924 57480 50930
rect 57428 50866 57480 50872
rect 57440 50522 57468 50866
rect 57428 50516 57480 50522
rect 57428 50458 57480 50464
rect 56600 50244 56652 50250
rect 56600 50186 56652 50192
rect 56324 49632 56376 49638
rect 56324 49574 56376 49580
rect 56336 49230 56364 49574
rect 56324 49224 56376 49230
rect 56324 49166 56376 49172
rect 56048 48748 56100 48754
rect 56048 48690 56100 48696
rect 55312 48680 55364 48686
rect 55312 48622 55364 48628
rect 56612 48278 56640 50186
rect 56784 49836 56836 49842
rect 56784 49778 56836 49784
rect 56692 49088 56744 49094
rect 56692 49030 56744 49036
rect 56600 48272 56652 48278
rect 56600 48214 56652 48220
rect 56704 48142 56732 49030
rect 56796 48890 56824 49778
rect 56784 48884 56836 48890
rect 56784 48826 56836 48832
rect 55312 48136 55364 48142
rect 55312 48078 55364 48084
rect 56692 48136 56744 48142
rect 56692 48078 56744 48084
rect 54116 48068 54168 48074
rect 54116 48010 54168 48016
rect 54128 47802 54156 48010
rect 54116 47796 54168 47802
rect 54116 47738 54168 47744
rect 53932 47252 53984 47258
rect 53932 47194 53984 47200
rect 53840 47048 53892 47054
rect 53840 46990 53892 46996
rect 55324 46986 55352 48078
rect 52736 46980 52788 46986
rect 52736 46922 52788 46928
rect 53656 46980 53708 46986
rect 53656 46922 53708 46928
rect 55312 46980 55364 46986
rect 55312 46922 55364 46928
rect 53668 46578 53696 46922
rect 53656 46572 53708 46578
rect 53656 46514 53708 46520
rect 55324 46510 55352 46922
rect 55496 46572 55548 46578
rect 55496 46514 55548 46520
rect 56692 46572 56744 46578
rect 56692 46514 56744 46520
rect 55312 46504 55364 46510
rect 55312 46446 55364 46452
rect 55036 46368 55088 46374
rect 55036 46310 55088 46316
rect 52552 46164 52604 46170
rect 52552 46106 52604 46112
rect 45744 45960 45796 45966
rect 45744 45902 45796 45908
rect 46940 45960 46992 45966
rect 46940 45902 46992 45908
rect 48964 45960 49016 45966
rect 48964 45902 49016 45908
rect 51540 45960 51592 45966
rect 51540 45902 51592 45908
rect 52460 45960 52512 45966
rect 52460 45902 52512 45908
rect 45652 45892 45704 45898
rect 45652 45834 45704 45840
rect 45664 45626 45692 45834
rect 45652 45620 45704 45626
rect 45652 45562 45704 45568
rect 44548 45552 44600 45558
rect 44548 45494 44600 45500
rect 44180 45348 44232 45354
rect 42444 44878 42472 45342
rect 44180 45290 44232 45296
rect 45756 44946 45784 45902
rect 46952 45490 46980 45902
rect 53380 45892 53432 45898
rect 53380 45834 53432 45840
rect 48228 45824 48280 45830
rect 48228 45766 48280 45772
rect 48240 45558 48268 45766
rect 50294 45724 50602 45744
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45648 50602 45668
rect 48228 45552 48280 45558
rect 48228 45494 48280 45500
rect 46940 45484 46992 45490
rect 46940 45426 46992 45432
rect 47584 45484 47636 45490
rect 47584 45426 47636 45432
rect 51540 45484 51592 45490
rect 51540 45426 51592 45432
rect 47596 44946 47624 45426
rect 49424 45416 49476 45422
rect 49424 45358 49476 45364
rect 48964 45280 49016 45286
rect 48964 45222 49016 45228
rect 45744 44940 45796 44946
rect 45744 44882 45796 44888
rect 47584 44940 47636 44946
rect 47584 44882 47636 44888
rect 42432 44872 42484 44878
rect 42432 44814 42484 44820
rect 41880 44804 41932 44810
rect 41880 44746 41932 44752
rect 41052 44736 41104 44742
rect 41052 44678 41104 44684
rect 41064 41614 41092 44678
rect 41788 44396 41840 44402
rect 41788 44338 41840 44344
rect 41800 41818 41828 44338
rect 41892 42566 41920 44746
rect 42444 44402 42472 44814
rect 42708 44804 42760 44810
rect 42708 44746 42760 44752
rect 42432 44396 42484 44402
rect 42432 44338 42484 44344
rect 42720 43994 42748 44746
rect 43812 44736 43864 44742
rect 43812 44678 43864 44684
rect 43824 44470 43852 44678
rect 45756 44470 45784 44882
rect 48976 44878 49004 45222
rect 48964 44872 49016 44878
rect 48964 44814 49016 44820
rect 48872 44804 48924 44810
rect 48872 44746 48924 44752
rect 47124 44736 47176 44742
rect 47124 44678 47176 44684
rect 43812 44464 43864 44470
rect 43812 44406 43864 44412
rect 45744 44464 45796 44470
rect 45744 44406 45796 44412
rect 44456 44396 44508 44402
rect 44456 44338 44508 44344
rect 42800 44192 42852 44198
rect 42800 44134 42852 44140
rect 42708 43988 42760 43994
rect 42708 43930 42760 43936
rect 42812 43790 42840 44134
rect 44468 43926 44496 44338
rect 45284 44328 45336 44334
rect 45756 44282 45784 44406
rect 46664 44396 46716 44402
rect 46664 44338 46716 44344
rect 45284 44270 45336 44276
rect 44456 43920 44508 43926
rect 44456 43862 44508 43868
rect 45296 43790 45324 44270
rect 45664 44254 45784 44282
rect 45664 43994 45692 44254
rect 46676 43994 46704 44338
rect 45652 43988 45704 43994
rect 45652 43930 45704 43936
rect 46664 43988 46716 43994
rect 46664 43930 46716 43936
rect 47136 43790 47164 44678
rect 48320 44396 48372 44402
rect 48320 44338 48372 44344
rect 47860 44192 47912 44198
rect 47860 44134 47912 44140
rect 42800 43784 42852 43790
rect 42800 43726 42852 43732
rect 44456 43784 44508 43790
rect 44456 43726 44508 43732
rect 45284 43784 45336 43790
rect 45284 43726 45336 43732
rect 47124 43784 47176 43790
rect 47124 43726 47176 43732
rect 42432 43240 42484 43246
rect 42432 43182 42484 43188
rect 42444 42922 42472 43182
rect 43076 43104 43128 43110
rect 43076 43046 43128 43052
rect 42444 42906 42564 42922
rect 42444 42900 42576 42906
rect 42444 42894 42524 42900
rect 42444 42702 42472 42894
rect 42524 42842 42576 42848
rect 42432 42696 42484 42702
rect 42432 42638 42484 42644
rect 41880 42560 41932 42566
rect 41880 42502 41932 42508
rect 41788 41812 41840 41818
rect 41788 41754 41840 41760
rect 41052 41608 41104 41614
rect 41052 41550 41104 41556
rect 42432 41608 42484 41614
rect 42432 41550 42484 41556
rect 41788 41132 41840 41138
rect 41788 41074 41840 41080
rect 41800 40730 41828 41074
rect 42444 41070 42472 41550
rect 42432 41064 42484 41070
rect 42432 41006 42484 41012
rect 41788 40724 41840 40730
rect 41788 40666 41840 40672
rect 42444 40526 42472 41006
rect 43088 40526 43116 43046
rect 44468 42906 44496 43726
rect 46480 43716 46532 43722
rect 46480 43658 46532 43664
rect 46492 43450 46520 43658
rect 46480 43444 46532 43450
rect 46480 43386 46532 43392
rect 46204 43376 46256 43382
rect 46204 43318 46256 43324
rect 45192 43308 45244 43314
rect 45192 43250 45244 43256
rect 44456 42900 44508 42906
rect 44456 42842 44508 42848
rect 44468 42702 44496 42842
rect 44456 42696 44508 42702
rect 44456 42638 44508 42644
rect 43812 42628 43864 42634
rect 43812 42570 43864 42576
rect 43824 41818 43852 42570
rect 44468 42362 44496 42638
rect 45100 42560 45152 42566
rect 45100 42502 45152 42508
rect 44456 42356 44508 42362
rect 44456 42298 44508 42304
rect 43812 41812 43864 41818
rect 43812 41754 43864 41760
rect 43720 41540 43772 41546
rect 43720 41482 43772 41488
rect 43732 41274 43760 41482
rect 43720 41268 43772 41274
rect 43720 41210 43772 41216
rect 43812 41132 43864 41138
rect 43812 41074 43864 41080
rect 43824 40730 43852 41074
rect 43812 40724 43864 40730
rect 43812 40666 43864 40672
rect 45112 40526 45140 42502
rect 45204 42226 45232 43250
rect 45192 42220 45244 42226
rect 45192 42162 45244 42168
rect 45204 41818 45232 42162
rect 45192 41812 45244 41818
rect 45192 41754 45244 41760
rect 45204 41138 45232 41754
rect 45192 41132 45244 41138
rect 45192 41074 45244 41080
rect 45204 40730 45232 41074
rect 46216 40730 46244 43318
rect 46388 43308 46440 43314
rect 46388 43250 46440 43256
rect 46400 42906 46428 43250
rect 46388 42900 46440 42906
rect 46388 42842 46440 42848
rect 47872 42702 47900 44134
rect 47952 43716 48004 43722
rect 47952 43658 48004 43664
rect 47860 42696 47912 42702
rect 47860 42638 47912 42644
rect 46756 42628 46808 42634
rect 46756 42570 46808 42576
rect 46768 42362 46796 42570
rect 46756 42356 46808 42362
rect 46756 42298 46808 42304
rect 46388 42220 46440 42226
rect 46388 42162 46440 42168
rect 46400 41818 46428 42162
rect 46388 41812 46440 41818
rect 46388 41754 46440 41760
rect 46572 41540 46624 41546
rect 46572 41482 46624 41488
rect 46584 41274 46612 41482
rect 46572 41268 46624 41274
rect 46572 41210 46624 41216
rect 46848 41132 46900 41138
rect 46848 41074 46900 41080
rect 45192 40724 45244 40730
rect 45192 40666 45244 40672
rect 46204 40724 46256 40730
rect 46204 40666 46256 40672
rect 42432 40520 42484 40526
rect 42432 40462 42484 40468
rect 43076 40520 43128 40526
rect 43076 40462 43128 40468
rect 45100 40520 45152 40526
rect 45100 40462 45152 40468
rect 42444 40050 42472 40462
rect 43720 40452 43772 40458
rect 43720 40394 43772 40400
rect 43732 40186 43760 40394
rect 43720 40180 43772 40186
rect 43720 40122 43772 40128
rect 45204 40050 45232 40666
rect 42432 40044 42484 40050
rect 42432 39986 42484 39992
rect 43812 40044 43864 40050
rect 43812 39986 43864 39992
rect 45192 40044 45244 40050
rect 45192 39986 45244 39992
rect 42444 39506 42472 39986
rect 43824 39642 43852 39986
rect 43812 39636 43864 39642
rect 43812 39578 43864 39584
rect 42432 39500 42484 39506
rect 42432 39442 42484 39448
rect 40960 39432 41012 39438
rect 40960 39374 41012 39380
rect 43720 39364 43772 39370
rect 43720 39306 43772 39312
rect 43732 39098 43760 39306
rect 43720 39092 43772 39098
rect 43720 39034 43772 39040
rect 45204 38962 45232 39986
rect 46204 39432 46256 39438
rect 46204 39374 46256 39380
rect 46216 38962 46244 39374
rect 43996 38956 44048 38962
rect 43996 38898 44048 38904
rect 45192 38956 45244 38962
rect 45192 38898 45244 38904
rect 46204 38956 46256 38962
rect 46204 38898 46256 38904
rect 42432 38888 42484 38894
rect 42432 38830 42484 38836
rect 42444 38350 42472 38830
rect 42432 38344 42484 38350
rect 42432 38286 42484 38292
rect 40500 37664 40552 37670
rect 40500 37606 40552 37612
rect 40408 37256 40460 37262
rect 40408 37198 40460 37204
rect 40512 36174 40540 37606
rect 42444 37466 42472 38286
rect 42432 37460 42484 37466
rect 42432 37402 42484 37408
rect 42444 36786 42472 37402
rect 42432 36780 42484 36786
rect 42432 36722 42484 36728
rect 42444 36174 42472 36722
rect 40500 36168 40552 36174
rect 40500 36110 40552 36116
rect 42432 36168 42484 36174
rect 42432 36110 42484 36116
rect 41420 36032 41472 36038
rect 41420 35974 41472 35980
rect 40328 35866 40540 35894
rect 39948 35148 40000 35154
rect 39948 35090 40000 35096
rect 40132 35012 40184 35018
rect 40132 34954 40184 34960
rect 39856 34400 39908 34406
rect 39856 34342 39908 34348
rect 39868 34066 39896 34342
rect 39856 34060 39908 34066
rect 39856 34002 39908 34008
rect 34796 33992 34848 33998
rect 34796 33934 34848 33940
rect 37924 33992 37976 33998
rect 37924 33934 37976 33940
rect 39120 33992 39172 33998
rect 39120 33934 39172 33940
rect 34704 33652 34756 33658
rect 34704 33594 34756 33600
rect 33876 33516 33928 33522
rect 34624 33510 34744 33538
rect 33876 33458 33928 33464
rect 33048 32904 33100 32910
rect 33048 32846 33100 32852
rect 32128 32836 32180 32842
rect 32128 32778 32180 32784
rect 31760 32564 31812 32570
rect 31760 32506 31812 32512
rect 31668 32428 31720 32434
rect 31668 32370 31720 32376
rect 31208 31952 31260 31958
rect 31208 31894 31260 31900
rect 30840 31476 30892 31482
rect 30840 31418 30892 31424
rect 31116 31476 31168 31482
rect 31116 31418 31168 31424
rect 29736 31340 29788 31346
rect 29736 31282 29788 31288
rect 29368 31136 29420 31142
rect 29368 31078 29420 31084
rect 29380 30734 29408 31078
rect 29368 30728 29420 30734
rect 29368 30670 29420 30676
rect 29276 30660 29328 30666
rect 29276 30602 29328 30608
rect 29748 30394 29776 31282
rect 29736 30388 29788 30394
rect 29736 30330 29788 30336
rect 29092 29844 29144 29850
rect 29092 29786 29144 29792
rect 29000 29640 29052 29646
rect 29000 29582 29052 29588
rect 30472 29504 30524 29510
rect 30472 29446 30524 29452
rect 30484 29238 30512 29446
rect 30472 29232 30524 29238
rect 30472 29174 30524 29180
rect 28816 29096 28868 29102
rect 28816 29038 28868 29044
rect 28828 28082 28856 29038
rect 29552 28552 29604 28558
rect 29552 28494 29604 28500
rect 28816 28076 28868 28082
rect 28816 28018 28868 28024
rect 29564 27878 29592 28494
rect 29552 27872 29604 27878
rect 29552 27814 29604 27820
rect 30104 27464 30156 27470
rect 30104 27406 30156 27412
rect 29000 27396 29052 27402
rect 29000 27338 29052 27344
rect 29012 26586 29040 27338
rect 30116 26994 30144 27406
rect 30104 26988 30156 26994
rect 30104 26930 30156 26936
rect 29000 26580 29052 26586
rect 29000 26522 29052 26528
rect 28908 26376 28960 26382
rect 28908 26318 28960 26324
rect 29552 26376 29604 26382
rect 29552 26318 29604 26324
rect 28460 26206 28580 26234
rect 28356 24812 28408 24818
rect 28356 24754 28408 24760
rect 27896 24608 27948 24614
rect 27896 24550 27948 24556
rect 27908 23118 27936 24550
rect 28368 23866 28396 24754
rect 28356 23860 28408 23866
rect 28356 23802 28408 23808
rect 27896 23112 27948 23118
rect 27896 23054 27948 23060
rect 27804 22704 27856 22710
rect 27804 22646 27856 22652
rect 27620 22432 27672 22438
rect 27620 22374 27672 22380
rect 27632 22030 27660 22374
rect 27620 22024 27672 22030
rect 27620 21966 27672 21972
rect 27632 21486 27660 21966
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 27632 21146 27660 21422
rect 27620 21140 27672 21146
rect 27620 21082 27672 21088
rect 26976 20936 27028 20942
rect 26976 20878 27028 20884
rect 26988 20398 27016 20878
rect 26976 20392 27028 20398
rect 26976 20334 27028 20340
rect 26988 19854 27016 20334
rect 26976 19848 27028 19854
rect 26976 19790 27028 19796
rect 25964 19780 26016 19786
rect 25964 19722 26016 19728
rect 23664 19304 23716 19310
rect 23664 19246 23716 19252
rect 23676 18290 23704 19246
rect 25044 19168 25096 19174
rect 25044 19110 25096 19116
rect 25056 18358 25084 19110
rect 25976 18766 26004 19722
rect 26988 19378 27016 19790
rect 28356 19780 28408 19786
rect 28356 19722 28408 19728
rect 28368 19514 28396 19722
rect 28356 19508 28408 19514
rect 28356 19450 28408 19456
rect 26976 19372 27028 19378
rect 26976 19314 27028 19320
rect 25964 18760 26016 18766
rect 25964 18702 26016 18708
rect 27620 18692 27672 18698
rect 27620 18634 27672 18640
rect 25044 18352 25096 18358
rect 25044 18294 25096 18300
rect 27632 18290 27660 18634
rect 23664 18284 23716 18290
rect 23664 18226 23716 18232
rect 27620 18284 27672 18290
rect 27620 18226 27672 18232
rect 23480 18148 23532 18154
rect 23480 18090 23532 18096
rect 22284 17876 22336 17882
rect 22284 17818 22336 17824
rect 23204 17604 23256 17610
rect 23204 17546 23256 17552
rect 23216 17338 23244 17546
rect 23204 17332 23256 17338
rect 23204 17274 23256 17280
rect 23676 17202 23704 18226
rect 25228 18080 25280 18086
rect 25228 18022 25280 18028
rect 25240 17678 25268 18022
rect 27632 17678 27660 18226
rect 24400 17672 24452 17678
rect 24400 17614 24452 17620
rect 25228 17672 25280 17678
rect 25228 17614 25280 17620
rect 27620 17672 27672 17678
rect 27620 17614 27672 17620
rect 24412 17202 24440 17614
rect 26516 17536 26568 17542
rect 26516 17478 26568 17484
rect 26528 17270 26556 17478
rect 26516 17264 26568 17270
rect 26516 17206 26568 17212
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 23204 17196 23256 17202
rect 23204 17138 23256 17144
rect 23664 17196 23716 17202
rect 23664 17138 23716 17144
rect 24400 17196 24452 17202
rect 24400 17138 24452 17144
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 22296 16182 22324 16390
rect 23216 16250 23244 17138
rect 24412 16658 24440 17138
rect 27632 17134 27660 17614
rect 27620 17128 27672 17134
rect 27620 17070 27672 17076
rect 25780 16992 25832 16998
rect 25780 16934 25832 16940
rect 24400 16652 24452 16658
rect 24400 16594 24452 16600
rect 25792 16590 25820 16934
rect 25780 16584 25832 16590
rect 25780 16526 25832 16532
rect 26240 16584 26292 16590
rect 26240 16526 26292 16532
rect 23480 16516 23532 16522
rect 23480 16458 23532 16464
rect 25872 16516 25924 16522
rect 25872 16458 25924 16464
rect 23204 16244 23256 16250
rect 23204 16186 23256 16192
rect 22284 16176 22336 16182
rect 22284 16118 22336 16124
rect 23492 15706 23520 16458
rect 25780 16448 25832 16454
rect 25780 16390 25832 16396
rect 25792 16182 25820 16390
rect 25780 16176 25832 16182
rect 25780 16118 25832 16124
rect 24400 16108 24452 16114
rect 24400 16050 24452 16056
rect 23480 15700 23532 15706
rect 23480 15642 23532 15648
rect 24412 15570 24440 16050
rect 25780 15904 25832 15910
rect 25780 15846 25832 15852
rect 24400 15564 24452 15570
rect 24400 15506 24452 15512
rect 23664 15428 23716 15434
rect 23664 15370 23716 15376
rect 23676 14618 23704 15370
rect 24412 15026 24440 15506
rect 25792 15502 25820 15846
rect 25884 15706 25912 16458
rect 26252 16250 26280 16526
rect 27068 16448 27120 16454
rect 27068 16390 27120 16396
rect 26240 16244 26292 16250
rect 26240 16186 26292 16192
rect 26792 16244 26844 16250
rect 26792 16186 26844 16192
rect 26332 16108 26384 16114
rect 26332 16050 26384 16056
rect 25872 15700 25924 15706
rect 25872 15642 25924 15648
rect 25780 15496 25832 15502
rect 25780 15438 25832 15444
rect 26344 15162 26372 16050
rect 26804 16046 26832 16186
rect 26792 16040 26844 16046
rect 26792 15982 26844 15988
rect 26804 15502 26832 15982
rect 26792 15496 26844 15502
rect 26792 15438 26844 15444
rect 26332 15156 26384 15162
rect 26332 15098 26384 15104
rect 26804 15026 26832 15438
rect 27080 15094 27108 16390
rect 28356 15904 28408 15910
rect 28356 15846 28408 15852
rect 28368 15502 28396 15846
rect 28356 15496 28408 15502
rect 28356 15438 28408 15444
rect 28172 15360 28224 15366
rect 28172 15302 28224 15308
rect 28184 15094 28212 15302
rect 27068 15088 27120 15094
rect 27068 15030 27120 15036
rect 28172 15088 28224 15094
rect 28172 15030 28224 15036
rect 24400 15020 24452 15026
rect 24400 14962 24452 14968
rect 26792 15020 26844 15026
rect 26792 14962 26844 14968
rect 23664 14612 23716 14618
rect 23664 14554 23716 14560
rect 24412 14414 24440 14962
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 26700 14816 26752 14822
rect 26700 14758 26752 14764
rect 28356 14816 28408 14822
rect 28356 14758 28408 14764
rect 24400 14408 24452 14414
rect 24400 14350 24452 14356
rect 21272 14340 21324 14346
rect 21272 14282 21324 14288
rect 22376 14340 22428 14346
rect 22376 14282 22428 14288
rect 23204 14340 23256 14346
rect 23204 14282 23256 14288
rect 21284 12986 21312 14282
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 21836 14006 21864 14214
rect 21824 14000 21876 14006
rect 21824 13942 21876 13948
rect 22192 14000 22244 14006
rect 22192 13942 22244 13948
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 22112 12918 22140 13126
rect 22100 12912 22152 12918
rect 22100 12854 22152 12860
rect 20916 11886 21036 11914
rect 19892 11688 19944 11694
rect 19892 11630 19944 11636
rect 19904 11150 19932 11630
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 20916 10742 20944 11886
rect 22204 11830 22232 13942
rect 22284 13252 22336 13258
rect 22284 13194 22336 13200
rect 22296 12442 22324 13194
rect 22284 12436 22336 12442
rect 22284 12378 22336 12384
rect 22388 11898 22416 14282
rect 23216 14074 23244 14282
rect 23204 14068 23256 14074
rect 23204 14010 23256 14016
rect 24412 13938 24440 14350
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 24412 13394 24440 13874
rect 24400 13388 24452 13394
rect 24400 13330 24452 13336
rect 24412 12850 24440 13330
rect 24504 12918 24532 14758
rect 26240 14340 26292 14346
rect 26240 14282 26292 14288
rect 24492 12912 24544 12918
rect 24492 12854 24544 12860
rect 24400 12844 24452 12850
rect 24400 12786 24452 12792
rect 24412 12306 24440 12786
rect 25136 12640 25188 12646
rect 25136 12582 25188 12588
rect 24124 12300 24176 12306
rect 24124 12242 24176 12248
rect 24400 12300 24452 12306
rect 24400 12242 24452 12248
rect 23480 12164 23532 12170
rect 23480 12106 23532 12112
rect 22376 11892 22428 11898
rect 22376 11834 22428 11840
rect 22192 11824 22244 11830
rect 22192 11766 22244 11772
rect 21272 11756 21324 11762
rect 21272 11698 21324 11704
rect 21284 11354 21312 11698
rect 22100 11552 22152 11558
rect 22100 11494 22152 11500
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 20996 11076 21048 11082
rect 20996 11018 21048 11024
rect 21008 10810 21036 11018
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 22112 10742 22140 11494
rect 23492 11354 23520 12106
rect 24136 11762 24164 12242
rect 25148 12238 25176 12582
rect 25136 12232 25188 12238
rect 25136 12174 25188 12180
rect 25780 12096 25832 12102
rect 25780 12038 25832 12044
rect 25792 11830 25820 12038
rect 25780 11824 25832 11830
rect 25780 11766 25832 11772
rect 24124 11756 24176 11762
rect 24124 11698 24176 11704
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 24136 11150 24164 11698
rect 25504 11552 25556 11558
rect 25504 11494 25556 11500
rect 25516 11150 25544 11494
rect 24124 11144 24176 11150
rect 24124 11086 24176 11092
rect 24400 11144 24452 11150
rect 24400 11086 24452 11092
rect 25504 11144 25556 11150
rect 25504 11086 25556 11092
rect 23204 11076 23256 11082
rect 23204 11018 23256 11024
rect 23216 10810 23244 11018
rect 23204 10804 23256 10810
rect 23204 10746 23256 10752
rect 20904 10736 20956 10742
rect 20904 10678 20956 10684
rect 22100 10736 22152 10742
rect 22100 10678 22152 10684
rect 24136 10674 24164 11086
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 24124 10668 24176 10674
rect 24124 10610 24176 10616
rect 20628 10600 20680 10606
rect 20628 10542 20680 10548
rect 20640 10266 20668 10542
rect 20628 10260 20680 10266
rect 20628 10202 20680 10208
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 20732 9722 20760 10610
rect 24412 10062 24440 11086
rect 25780 11008 25832 11014
rect 25780 10950 25832 10956
rect 25792 10742 25820 10950
rect 25780 10736 25832 10742
rect 25780 10678 25832 10684
rect 25412 10464 25464 10470
rect 25412 10406 25464 10412
rect 25424 10062 25452 10406
rect 26252 10266 26280 14282
rect 26424 13728 26476 13734
rect 26424 13670 26476 13676
rect 26436 13326 26464 13670
rect 26712 13530 26740 14758
rect 27528 14340 27580 14346
rect 27528 14282 27580 14288
rect 27540 13938 27568 14282
rect 28368 14006 28396 14758
rect 28356 14000 28408 14006
rect 28356 13942 28408 13948
rect 27068 13932 27120 13938
rect 27068 13874 27120 13880
rect 27528 13932 27580 13938
rect 27528 13874 27580 13880
rect 26700 13524 26752 13530
rect 26700 13466 26752 13472
rect 27080 13394 27108 13874
rect 28356 13728 28408 13734
rect 28356 13670 28408 13676
rect 27068 13388 27120 13394
rect 27068 13330 27120 13336
rect 28368 13326 28396 13670
rect 26424 13320 26476 13326
rect 26424 13262 26476 13268
rect 28356 13320 28408 13326
rect 28356 13262 28408 13268
rect 27344 12844 27396 12850
rect 27344 12786 27396 12792
rect 27356 12730 27384 12786
rect 27356 12702 27476 12730
rect 27448 12238 27476 12702
rect 27436 12232 27488 12238
rect 27436 12174 27488 12180
rect 27448 11762 27476 12174
rect 27436 11756 27488 11762
rect 27436 11698 27488 11704
rect 27528 10668 27580 10674
rect 27528 10610 27580 10616
rect 26240 10260 26292 10266
rect 26240 10202 26292 10208
rect 26252 10062 26280 10202
rect 24400 10056 24452 10062
rect 24400 9998 24452 10004
rect 25412 10056 25464 10062
rect 25412 9998 25464 10004
rect 26240 10056 26292 10062
rect 26240 9998 26292 10004
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 24412 9654 24440 9998
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 24400 9648 24452 9654
rect 24400 9590 24452 9596
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19352 9042 19380 9454
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19352 8634 19380 8978
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 20548 8634 20576 9522
rect 24412 8974 24440 9590
rect 24952 9580 25004 9586
rect 24952 9522 25004 9528
rect 24584 9376 24636 9382
rect 24584 9318 24636 9324
rect 23848 8968 23900 8974
rect 23848 8910 23900 8916
rect 24400 8968 24452 8974
rect 24400 8910 24452 8916
rect 22008 8900 22060 8906
rect 22008 8842 22060 8848
rect 23388 8900 23440 8906
rect 23388 8842 23440 8848
rect 21732 8832 21784 8838
rect 21732 8774 21784 8780
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 21744 8566 21772 8774
rect 21732 8560 21784 8566
rect 21732 8502 21784 8508
rect 21640 8424 21692 8430
rect 21640 8366 21692 8372
rect 21652 7886 21680 8366
rect 22020 8090 22048 8842
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 22008 8084 22060 8090
rect 22008 8026 22060 8032
rect 22204 7886 22232 8774
rect 23400 8634 23428 8842
rect 23388 8628 23440 8634
rect 23388 8570 23440 8576
rect 23860 8430 23888 8910
rect 24596 8566 24624 9318
rect 24964 8634 24992 9522
rect 25148 8974 25176 9862
rect 27540 9654 27568 10610
rect 26240 9648 26292 9654
rect 26240 9590 26292 9596
rect 27528 9648 27580 9654
rect 27528 9590 27580 9596
rect 25780 9580 25832 9586
rect 25780 9522 25832 9528
rect 25792 9178 25820 9522
rect 25780 9172 25832 9178
rect 25780 9114 25832 9120
rect 26252 9042 26280 9590
rect 27620 9580 27672 9586
rect 27620 9522 27672 9528
rect 26516 9376 26568 9382
rect 26516 9318 26568 9324
rect 26240 9036 26292 9042
rect 26240 8978 26292 8984
rect 25136 8968 25188 8974
rect 25136 8910 25188 8916
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 24584 8560 24636 8566
rect 24584 8502 24636 8508
rect 26252 8498 26280 8978
rect 26528 8974 26556 9318
rect 27632 9178 27660 9522
rect 28356 9376 28408 9382
rect 28356 9318 28408 9324
rect 27620 9172 27672 9178
rect 27620 9114 27672 9120
rect 26516 8968 26568 8974
rect 26516 8910 26568 8916
rect 25780 8492 25832 8498
rect 25780 8434 25832 8440
rect 26240 8492 26292 8498
rect 26240 8434 26292 8440
rect 27620 8492 27672 8498
rect 27620 8434 27672 8440
rect 23848 8424 23900 8430
rect 23848 8366 23900 8372
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 22008 7812 22060 7818
rect 22008 7754 22060 7760
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 20732 7478 20760 7686
rect 21100 7546 21128 7754
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 20720 7472 20772 7478
rect 20720 7414 20772 7420
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 19708 7336 19760 7342
rect 19708 7278 19760 7284
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 19260 6798 19288 7142
rect 19720 6798 19748 7278
rect 21192 7002 21220 7346
rect 21180 6996 21232 7002
rect 21180 6938 21232 6944
rect 22020 6798 22048 7754
rect 23860 7342 23888 8366
rect 25792 8090 25820 8434
rect 25780 8084 25832 8090
rect 25780 8026 25832 8032
rect 26252 7954 26280 8434
rect 27632 8090 27660 8434
rect 27620 8084 27672 8090
rect 27620 8026 27672 8032
rect 26240 7948 26292 7954
rect 26240 7890 26292 7896
rect 28368 7886 28396 9318
rect 24308 7880 24360 7886
rect 24308 7822 24360 7828
rect 28356 7880 28408 7886
rect 28356 7822 28408 7828
rect 23848 7336 23900 7342
rect 23848 7278 23900 7284
rect 24320 6798 24348 7822
rect 25228 7812 25280 7818
rect 25228 7754 25280 7760
rect 26976 7812 27028 7818
rect 26976 7754 27028 7760
rect 25240 7546 25268 7754
rect 25228 7540 25280 7546
rect 25228 7482 25280 7488
rect 24400 7472 24452 7478
rect 24400 7414 24452 7420
rect 24412 6866 24440 7414
rect 26988 7410 27016 7754
rect 25780 7404 25832 7410
rect 25780 7346 25832 7352
rect 26976 7404 27028 7410
rect 26976 7346 27028 7352
rect 25792 7002 25820 7346
rect 25780 6996 25832 7002
rect 25780 6938 25832 6944
rect 28460 6914 28488 26206
rect 28920 24818 28948 26318
rect 29092 25696 29144 25702
rect 29092 25638 29144 25644
rect 28908 24812 28960 24818
rect 28908 24754 28960 24760
rect 29104 23798 29132 25638
rect 29564 25362 29592 26318
rect 30116 25906 30144 26930
rect 30196 26784 30248 26790
rect 30196 26726 30248 26732
rect 30208 26382 30236 26726
rect 30196 26376 30248 26382
rect 30196 26318 30248 26324
rect 30104 25900 30156 25906
rect 30104 25842 30156 25848
rect 30840 25900 30892 25906
rect 30840 25842 30892 25848
rect 29552 25356 29604 25362
rect 29552 25298 29604 25304
rect 30116 25294 30144 25842
rect 30852 25498 30880 25842
rect 30840 25492 30892 25498
rect 30840 25434 30892 25440
rect 30104 25288 30156 25294
rect 30104 25230 30156 25236
rect 30196 25220 30248 25226
rect 30196 25162 30248 25168
rect 30208 24954 30236 25162
rect 30196 24948 30248 24954
rect 30196 24890 30248 24896
rect 30932 24812 30984 24818
rect 30932 24754 30984 24760
rect 30944 24410 30972 24754
rect 30932 24404 30984 24410
rect 30932 24346 30984 24352
rect 30288 24200 30340 24206
rect 30288 24142 30340 24148
rect 29092 23792 29144 23798
rect 29092 23734 29144 23740
rect 30196 23520 30248 23526
rect 30196 23462 30248 23468
rect 30208 22710 30236 23462
rect 30300 23202 30328 24142
rect 30932 24132 30984 24138
rect 30932 24074 30984 24080
rect 30300 23186 30420 23202
rect 30300 23180 30432 23186
rect 30300 23174 30380 23180
rect 30380 23122 30432 23128
rect 30840 23180 30892 23186
rect 30840 23122 30892 23128
rect 30196 22704 30248 22710
rect 30196 22646 30248 22652
rect 30852 22098 30880 23122
rect 30944 22778 30972 24074
rect 30932 22772 30984 22778
rect 30932 22714 30984 22720
rect 31128 22710 31156 31418
rect 31220 30326 31248 31894
rect 32140 31822 32168 32778
rect 33324 32768 33376 32774
rect 33324 32710 33376 32716
rect 33336 32502 33364 32710
rect 33324 32496 33376 32502
rect 33324 32438 33376 32444
rect 33508 32224 33560 32230
rect 33508 32166 33560 32172
rect 33520 31822 33548 32166
rect 33888 32026 33916 33458
rect 34716 33318 34744 33510
rect 37936 33454 37964 33934
rect 39672 33924 39724 33930
rect 39672 33866 39724 33872
rect 39304 33856 39356 33862
rect 39304 33798 39356 33804
rect 39316 33590 39344 33798
rect 39684 33658 39712 33866
rect 39672 33652 39724 33658
rect 39672 33594 39724 33600
rect 39304 33584 39356 33590
rect 39304 33526 39356 33532
rect 37924 33448 37976 33454
rect 37924 33390 37976 33396
rect 34704 33312 34756 33318
rect 34704 33254 34756 33260
rect 34612 32836 34664 32842
rect 34612 32778 34664 32784
rect 33876 32020 33928 32026
rect 33876 31962 33928 31968
rect 31484 31816 31536 31822
rect 31484 31758 31536 31764
rect 32128 31816 32180 31822
rect 32128 31758 32180 31764
rect 33508 31816 33560 31822
rect 33508 31758 33560 31764
rect 31208 30320 31260 30326
rect 31208 30262 31260 30268
rect 31392 30252 31444 30258
rect 31392 30194 31444 30200
rect 31404 29850 31432 30194
rect 31496 30122 31524 31758
rect 32140 30734 32168 31758
rect 34624 31482 34652 32778
rect 34716 32434 34744 33254
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 37004 33108 37056 33114
rect 37004 33050 37056 33056
rect 35900 32904 35952 32910
rect 35900 32846 35952 32852
rect 34704 32428 34756 32434
rect 34704 32370 34756 32376
rect 34612 31476 34664 31482
rect 34612 31418 34664 31424
rect 33600 31408 33652 31414
rect 33600 31350 33652 31356
rect 33232 31272 33284 31278
rect 33232 31214 33284 31220
rect 33244 30938 33272 31214
rect 33232 30932 33284 30938
rect 33232 30874 33284 30880
rect 32128 30728 32180 30734
rect 32128 30670 32180 30676
rect 31760 30592 31812 30598
rect 31760 30534 31812 30540
rect 31576 30252 31628 30258
rect 31576 30194 31628 30200
rect 31484 30116 31536 30122
rect 31484 30058 31536 30064
rect 31392 29844 31444 29850
rect 31392 29786 31444 29792
rect 31588 29306 31616 30194
rect 31772 29646 31800 30534
rect 32140 30190 32168 30670
rect 33508 30660 33560 30666
rect 33508 30602 33560 30608
rect 33520 30394 33548 30602
rect 33508 30388 33560 30394
rect 33508 30330 33560 30336
rect 32128 30184 32180 30190
rect 32128 30126 32180 30132
rect 31760 29640 31812 29646
rect 31760 29582 31812 29588
rect 31944 29640 31996 29646
rect 32140 29628 32168 30126
rect 31996 29600 32168 29628
rect 31944 29582 31996 29588
rect 31576 29300 31628 29306
rect 31576 29242 31628 29248
rect 32140 29170 32168 29600
rect 32128 29164 32180 29170
rect 32128 29106 32180 29112
rect 33140 28484 33192 28490
rect 33140 28426 33192 28432
rect 31484 28416 31536 28422
rect 31484 28358 31536 28364
rect 31496 27470 31524 28358
rect 32680 28076 32732 28082
rect 32680 28018 32732 28024
rect 31484 27464 31536 27470
rect 31484 27406 31536 27412
rect 32588 27396 32640 27402
rect 32588 27338 32640 27344
rect 32404 26784 32456 26790
rect 32404 26726 32456 26732
rect 31208 26512 31260 26518
rect 31208 26454 31260 26460
rect 31220 24138 31248 26454
rect 31300 26308 31352 26314
rect 31300 26250 31352 26256
rect 31312 26042 31340 26250
rect 31300 26036 31352 26042
rect 31300 25978 31352 25984
rect 31392 25288 31444 25294
rect 31392 25230 31444 25236
rect 31404 24818 31432 25230
rect 32416 24818 32444 26726
rect 31392 24812 31444 24818
rect 31392 24754 31444 24760
rect 32404 24812 32456 24818
rect 32404 24754 32456 24760
rect 31404 24274 31432 24754
rect 32404 24608 32456 24614
rect 32404 24550 32456 24556
rect 31392 24268 31444 24274
rect 31392 24210 31444 24216
rect 31208 24132 31260 24138
rect 31208 24074 31260 24080
rect 31404 23730 31432 24210
rect 32416 23798 32444 24550
rect 32600 24410 32628 27338
rect 32692 25498 32720 28018
rect 32772 27328 32824 27334
rect 32772 27270 32824 27276
rect 32784 26382 32812 27270
rect 33152 26994 33180 28426
rect 33508 27872 33560 27878
rect 33508 27814 33560 27820
rect 33520 27062 33548 27814
rect 33508 27056 33560 27062
rect 33508 26998 33560 27004
rect 33140 26988 33192 26994
rect 33140 26930 33192 26936
rect 32772 26376 32824 26382
rect 32772 26318 32824 26324
rect 32772 26240 32824 26246
rect 32772 26182 32824 26188
rect 32680 25492 32732 25498
rect 32680 25434 32732 25440
rect 32784 25294 32812 26182
rect 32956 25900 33008 25906
rect 32956 25842 33008 25848
rect 32772 25288 32824 25294
rect 32772 25230 32824 25236
rect 32588 24404 32640 24410
rect 32588 24346 32640 24352
rect 32404 23792 32456 23798
rect 32404 23734 32456 23740
rect 31392 23724 31444 23730
rect 31392 23666 31444 23672
rect 32772 23112 32824 23118
rect 32772 23054 32824 23060
rect 31852 23044 31904 23050
rect 31852 22986 31904 22992
rect 31116 22704 31168 22710
rect 31116 22646 31168 22652
rect 31864 22234 31892 22986
rect 32312 22976 32364 22982
rect 32312 22918 32364 22924
rect 31852 22228 31904 22234
rect 31852 22170 31904 22176
rect 30840 22092 30892 22098
rect 30840 22034 30892 22040
rect 28908 21956 28960 21962
rect 28908 21898 28960 21904
rect 28920 21690 28948 21898
rect 29000 21888 29052 21894
rect 29000 21830 29052 21836
rect 28908 21684 28960 21690
rect 28908 21626 28960 21632
rect 28816 21548 28868 21554
rect 28816 21490 28868 21496
rect 28828 21146 28856 21490
rect 28816 21140 28868 21146
rect 28816 21082 28868 21088
rect 28908 20868 28960 20874
rect 28908 20810 28960 20816
rect 28540 20460 28592 20466
rect 28540 20402 28592 20408
rect 28552 20058 28580 20402
rect 28724 20256 28776 20262
rect 28724 20198 28776 20204
rect 28540 20052 28592 20058
rect 28540 19994 28592 20000
rect 28736 18358 28764 20198
rect 28920 18426 28948 20810
rect 29012 20534 29040 21830
rect 30852 21554 30880 22034
rect 32324 21622 32352 22918
rect 32784 22642 32812 23054
rect 32772 22636 32824 22642
rect 32772 22578 32824 22584
rect 32312 21616 32364 21622
rect 32312 21558 32364 21564
rect 30012 21548 30064 21554
rect 30012 21490 30064 21496
rect 30840 21548 30892 21554
rect 30840 21490 30892 21496
rect 30024 21010 30052 21490
rect 31576 21344 31628 21350
rect 31576 21286 31628 21292
rect 30012 21004 30064 21010
rect 30012 20946 30064 20952
rect 29000 20528 29052 20534
rect 29000 20470 29052 20476
rect 30024 20466 30052 20946
rect 31588 20942 31616 21286
rect 32968 20942 32996 25842
rect 33612 23730 33640 31350
rect 34716 31346 34744 32370
rect 35912 32366 35940 32846
rect 36452 32768 36504 32774
rect 36452 32710 36504 32716
rect 36360 32428 36412 32434
rect 36360 32370 36412 32376
rect 35900 32360 35952 32366
rect 35900 32302 35952 32308
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 35912 31890 35940 32302
rect 35992 32224 36044 32230
rect 35992 32166 36044 32172
rect 35900 31884 35952 31890
rect 35900 31826 35952 31832
rect 34704 31340 34756 31346
rect 34704 31282 34756 31288
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 36004 30734 36032 32166
rect 36372 31482 36400 32370
rect 36464 31822 36492 32710
rect 36452 31816 36504 31822
rect 36452 31758 36504 31764
rect 36360 31476 36412 31482
rect 36360 31418 36412 31424
rect 34704 30728 34756 30734
rect 34704 30670 34756 30676
rect 35992 30728 36044 30734
rect 35992 30670 36044 30676
rect 34716 30054 34744 30670
rect 36084 30592 36136 30598
rect 36084 30534 36136 30540
rect 34704 30048 34756 30054
rect 34704 29990 34756 29996
rect 34716 29646 34744 29990
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 36096 29646 36124 30534
rect 34704 29640 34756 29646
rect 34704 29582 34756 29588
rect 36084 29640 36136 29646
rect 36084 29582 36136 29588
rect 33784 29572 33836 29578
rect 33784 29514 33836 29520
rect 33796 28762 33824 29514
rect 34716 29102 34744 29582
rect 36084 29504 36136 29510
rect 36084 29446 36136 29452
rect 36096 29238 36124 29446
rect 36084 29232 36136 29238
rect 36084 29174 36136 29180
rect 35992 29164 36044 29170
rect 35992 29106 36044 29112
rect 34704 29096 34756 29102
rect 34704 29038 34756 29044
rect 34244 28960 34296 28966
rect 34244 28902 34296 28908
rect 33784 28756 33836 28762
rect 33784 28698 33836 28704
rect 34256 28558 34284 28902
rect 34716 28558 34744 29038
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34244 28552 34296 28558
rect 34244 28494 34296 28500
rect 34704 28552 34756 28558
rect 34704 28494 34756 28500
rect 34716 28014 34744 28494
rect 34704 28008 34756 28014
rect 34704 27950 34756 27956
rect 34716 27470 34744 27950
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34704 27464 34756 27470
rect 34704 27406 34756 27412
rect 34716 26994 34744 27406
rect 34704 26988 34756 26994
rect 34704 26930 34756 26936
rect 35716 26988 35768 26994
rect 35716 26930 35768 26936
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 33968 26376 34020 26382
rect 33968 26318 34020 26324
rect 33980 25702 34008 26318
rect 34520 26308 34572 26314
rect 34520 26250 34572 26256
rect 33968 25696 34020 25702
rect 33968 25638 34020 25644
rect 33980 24750 34008 25638
rect 33968 24744 34020 24750
rect 33968 24686 34020 24692
rect 33980 24274 34008 24686
rect 33968 24268 34020 24274
rect 33968 24210 34020 24216
rect 33600 23724 33652 23730
rect 33600 23666 33652 23672
rect 33980 23662 34008 24210
rect 34532 23866 34560 26250
rect 35440 25696 35492 25702
rect 35440 25638 35492 25644
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 35452 25226 35480 25638
rect 35728 25362 35756 26930
rect 36004 26858 36032 29106
rect 36084 28960 36136 28966
rect 36084 28902 36136 28908
rect 36096 28558 36124 28902
rect 36084 28552 36136 28558
rect 36084 28494 36136 28500
rect 36176 28416 36228 28422
rect 36176 28358 36228 28364
rect 36188 28150 36216 28358
rect 36176 28144 36228 28150
rect 36176 28086 36228 28092
rect 36176 27872 36228 27878
rect 36176 27814 36228 27820
rect 36188 27470 36216 27814
rect 36176 27464 36228 27470
rect 36176 27406 36228 27412
rect 36084 27328 36136 27334
rect 36084 27270 36136 27276
rect 36096 27062 36124 27270
rect 36084 27056 36136 27062
rect 36084 26998 36136 27004
rect 35992 26852 36044 26858
rect 35992 26794 36044 26800
rect 36176 26308 36228 26314
rect 36176 26250 36228 26256
rect 36084 26240 36136 26246
rect 36084 26182 36136 26188
rect 36096 25974 36124 26182
rect 36084 25968 36136 25974
rect 36084 25910 36136 25916
rect 35716 25356 35768 25362
rect 35716 25298 35768 25304
rect 35440 25220 35492 25226
rect 35440 25162 35492 25168
rect 36084 25152 36136 25158
rect 36084 25094 36136 25100
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 36096 24206 36124 25094
rect 36084 24200 36136 24206
rect 36084 24142 36136 24148
rect 35348 24132 35400 24138
rect 35348 24074 35400 24080
rect 34520 23860 34572 23866
rect 34520 23802 34572 23808
rect 33968 23656 34020 23662
rect 33968 23598 34020 23604
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34796 23044 34848 23050
rect 34796 22986 34848 22992
rect 33508 22976 33560 22982
rect 33508 22918 33560 22924
rect 31576 20936 31628 20942
rect 31576 20878 31628 20884
rect 32956 20936 33008 20942
rect 32956 20878 33008 20884
rect 31392 20800 31444 20806
rect 31392 20742 31444 20748
rect 32496 20800 32548 20806
rect 32496 20742 32548 20748
rect 30012 20460 30064 20466
rect 30012 20402 30064 20408
rect 30024 19922 30052 20402
rect 30012 19916 30064 19922
rect 30012 19858 30064 19864
rect 30024 19378 30052 19858
rect 31404 19854 31432 20742
rect 32128 20460 32180 20466
rect 32128 20402 32180 20408
rect 32140 20058 32168 20402
rect 32508 20398 32536 20742
rect 33520 20534 33548 22918
rect 34152 22636 34204 22642
rect 34152 22578 34204 22584
rect 34164 22234 34192 22578
rect 34520 22432 34572 22438
rect 34520 22374 34572 22380
rect 34152 22228 34204 22234
rect 34152 22170 34204 22176
rect 33876 21888 33928 21894
rect 33876 21830 33928 21836
rect 33888 20602 33916 21830
rect 34532 21622 34560 22374
rect 34808 21690 34836 22986
rect 35360 22642 35388 24074
rect 36084 24064 36136 24070
rect 36084 24006 36136 24012
rect 36096 23798 36124 24006
rect 36188 23866 36216 26250
rect 36176 23860 36228 23866
rect 36176 23802 36228 23808
rect 36084 23792 36136 23798
rect 36084 23734 36136 23740
rect 36084 23112 36136 23118
rect 36084 23054 36136 23060
rect 35348 22636 35400 22642
rect 35348 22578 35400 22584
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 36096 22030 36124 23054
rect 36544 23044 36596 23050
rect 36544 22986 36596 22992
rect 36084 22024 36136 22030
rect 36084 21966 36136 21972
rect 34796 21684 34848 21690
rect 34796 21626 34848 21632
rect 36096 21622 36124 21966
rect 36268 21956 36320 21962
rect 36268 21898 36320 21904
rect 34520 21616 34572 21622
rect 34520 21558 34572 21564
rect 36084 21616 36136 21622
rect 36084 21558 36136 21564
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 36096 20942 36124 21558
rect 34980 20936 35032 20942
rect 34980 20878 35032 20884
rect 36084 20936 36136 20942
rect 36084 20878 36136 20884
rect 33876 20596 33928 20602
rect 33876 20538 33928 20544
rect 34992 20534 35020 20878
rect 33508 20528 33560 20534
rect 33508 20470 33560 20476
rect 34980 20528 35032 20534
rect 34980 20470 35032 20476
rect 32496 20392 32548 20398
rect 32496 20334 32548 20340
rect 36096 20262 36124 20878
rect 32680 20256 32732 20262
rect 32680 20198 32732 20204
rect 36084 20256 36136 20262
rect 36084 20198 36136 20204
rect 32128 20052 32180 20058
rect 32128 19994 32180 20000
rect 32128 19916 32180 19922
rect 32128 19858 32180 19864
rect 31392 19848 31444 19854
rect 31392 19790 31444 19796
rect 31760 19712 31812 19718
rect 31760 19654 31812 19660
rect 31208 19440 31260 19446
rect 31208 19382 31260 19388
rect 30012 19372 30064 19378
rect 30012 19314 30064 19320
rect 30024 18442 30052 19314
rect 28908 18420 28960 18426
rect 28908 18362 28960 18368
rect 29932 18414 30052 18442
rect 31220 18426 31248 19382
rect 31772 18766 31800 19654
rect 32140 19310 32168 19858
rect 32692 19854 32720 20198
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 36096 20058 36124 20198
rect 36280 20058 36308 21898
rect 36556 21690 36584 22986
rect 36636 22976 36688 22982
rect 36636 22918 36688 22924
rect 36544 21684 36596 21690
rect 36544 21626 36596 21632
rect 36084 20052 36136 20058
rect 36084 19994 36136 20000
rect 36268 20052 36320 20058
rect 36268 19994 36320 20000
rect 32680 19848 32732 19854
rect 32680 19790 32732 19796
rect 34520 19508 34572 19514
rect 34520 19450 34572 19456
rect 32220 19372 32272 19378
rect 32220 19314 32272 19320
rect 32128 19304 32180 19310
rect 32128 19246 32180 19252
rect 32232 18970 32260 19314
rect 33508 19168 33560 19174
rect 33508 19110 33560 19116
rect 32220 18964 32272 18970
rect 32220 18906 32272 18912
rect 31760 18760 31812 18766
rect 31760 18702 31812 18708
rect 32772 18692 32824 18698
rect 32772 18634 32824 18640
rect 31208 18420 31260 18426
rect 28724 18352 28776 18358
rect 28724 18294 28776 18300
rect 29932 18290 29960 18414
rect 31208 18362 31260 18368
rect 29920 18284 29972 18290
rect 29920 18226 29972 18232
rect 29932 17746 29960 18226
rect 32784 18222 32812 18634
rect 33520 18358 33548 19110
rect 34532 18358 34560 19450
rect 36096 19446 36124 19994
rect 36648 19854 36676 22918
rect 36728 22432 36780 22438
rect 36728 22374 36780 22380
rect 36740 20942 36768 22374
rect 36728 20936 36780 20942
rect 36728 20878 36780 20884
rect 36636 19848 36688 19854
rect 36636 19790 36688 19796
rect 36084 19440 36136 19446
rect 36084 19382 36136 19388
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 36096 18766 36124 19382
rect 36728 19372 36780 19378
rect 36728 19314 36780 19320
rect 36084 18760 36136 18766
rect 36084 18702 36136 18708
rect 36096 18358 36124 18702
rect 36740 18426 36768 19314
rect 36728 18420 36780 18426
rect 36728 18362 36780 18368
rect 33508 18352 33560 18358
rect 33508 18294 33560 18300
rect 34520 18352 34572 18358
rect 34520 18294 34572 18300
rect 36084 18352 36136 18358
rect 36084 18294 36136 18300
rect 32772 18216 32824 18222
rect 32772 18158 32824 18164
rect 32784 17746 32812 18158
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 29920 17740 29972 17746
rect 29920 17682 29972 17688
rect 32772 17740 32824 17746
rect 32772 17682 32824 17688
rect 29736 17604 29788 17610
rect 29736 17546 29788 17552
rect 29000 17536 29052 17542
rect 29000 17478 29052 17484
rect 29012 17338 29040 17478
rect 29000 17332 29052 17338
rect 29000 17274 29052 17280
rect 29748 17066 29776 17546
rect 29932 17134 29960 17682
rect 31576 17604 31628 17610
rect 31576 17546 31628 17552
rect 30472 17536 30524 17542
rect 30472 17478 30524 17484
rect 30484 17270 30512 17478
rect 30472 17264 30524 17270
rect 30472 17206 30524 17212
rect 29920 17128 29972 17134
rect 29920 17070 29972 17076
rect 29736 17060 29788 17066
rect 29736 17002 29788 17008
rect 31588 16250 31616 17546
rect 32784 17270 32812 17682
rect 35348 17604 35400 17610
rect 35348 17546 35400 17552
rect 34796 17536 34848 17542
rect 34796 17478 34848 17484
rect 32772 17264 32824 17270
rect 32772 17206 32824 17212
rect 33508 17196 33560 17202
rect 33508 17138 33560 17144
rect 32312 16992 32364 16998
rect 32312 16934 32364 16940
rect 33232 16992 33284 16998
rect 33232 16934 33284 16940
rect 31760 16584 31812 16590
rect 31760 16526 31812 16532
rect 31576 16244 31628 16250
rect 31576 16186 31628 16192
rect 31772 16114 31800 16526
rect 31852 16516 31904 16522
rect 31852 16458 31904 16464
rect 31760 16108 31812 16114
rect 31760 16050 31812 16056
rect 28816 14952 28868 14958
rect 28816 14894 28868 14900
rect 28828 14414 28856 14894
rect 30196 14816 30248 14822
rect 30196 14758 30248 14764
rect 28816 14408 28868 14414
rect 28816 14350 28868 14356
rect 30208 14074 30236 14758
rect 31864 14618 31892 16458
rect 32220 16448 32272 16454
rect 32220 16390 32272 16396
rect 32232 16182 32260 16390
rect 32324 16250 32352 16934
rect 32312 16244 32364 16250
rect 32312 16186 32364 16192
rect 32220 16176 32272 16182
rect 32220 16118 32272 16124
rect 32864 16108 32916 16114
rect 32864 16050 32916 16056
rect 32876 15502 32904 16050
rect 32864 15496 32916 15502
rect 32864 15438 32916 15444
rect 32128 15360 32180 15366
rect 32128 15302 32180 15308
rect 31852 14612 31904 14618
rect 31852 14554 31904 14560
rect 32140 14414 32168 15302
rect 32876 14958 32904 15438
rect 33244 15094 33272 16934
rect 33520 16250 33548 17138
rect 33508 16244 33560 16250
rect 33508 16186 33560 16192
rect 34808 16182 34836 17478
rect 35360 17338 35388 17546
rect 35348 17332 35400 17338
rect 35348 17274 35400 17280
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 36096 16658 36124 18294
rect 36360 18080 36412 18086
rect 36360 18022 36412 18028
rect 36084 16652 36136 16658
rect 36084 16594 36136 16600
rect 36372 16590 36400 18022
rect 37016 17338 37044 33050
rect 37936 32502 37964 33390
rect 39868 33318 39896 34002
rect 40144 33590 40172 34954
rect 40132 33584 40184 33590
rect 40132 33526 40184 33532
rect 39856 33312 39908 33318
rect 39856 33254 39908 33260
rect 39868 32978 39896 33254
rect 39856 32972 39908 32978
rect 39856 32914 39908 32920
rect 38660 32836 38712 32842
rect 38660 32778 38712 32784
rect 38672 32570 38700 32778
rect 38660 32564 38712 32570
rect 38660 32506 38712 32512
rect 37924 32496 37976 32502
rect 37924 32438 37976 32444
rect 37280 32360 37332 32366
rect 37280 32302 37332 32308
rect 37292 31890 37320 32302
rect 37936 31890 37964 32438
rect 39304 32428 39356 32434
rect 39304 32370 39356 32376
rect 40408 32428 40460 32434
rect 40408 32370 40460 32376
rect 39316 32026 39344 32370
rect 39304 32020 39356 32026
rect 39304 31962 39356 31968
rect 40420 31890 40448 32370
rect 37280 31884 37332 31890
rect 37280 31826 37332 31832
rect 37924 31884 37976 31890
rect 37924 31826 37976 31832
rect 40408 31884 40460 31890
rect 40408 31826 40460 31832
rect 37280 31680 37332 31686
rect 37280 31622 37332 31628
rect 37292 31414 37320 31622
rect 37280 31408 37332 31414
rect 37280 31350 37332 31356
rect 37936 31346 37964 31826
rect 39304 31816 39356 31822
rect 39304 31758 39356 31764
rect 37924 31340 37976 31346
rect 37924 31282 37976 31288
rect 39316 30938 39344 31758
rect 40512 31414 40540 35866
rect 41432 35766 41460 35974
rect 42444 35894 42472 36110
rect 42444 35866 42564 35894
rect 41420 35760 41472 35766
rect 41420 35702 41472 35708
rect 42536 35698 42564 35866
rect 42524 35692 42576 35698
rect 42576 35652 42656 35680
rect 42524 35634 42576 35640
rect 40684 35488 40736 35494
rect 40684 35430 40736 35436
rect 40696 35086 40724 35430
rect 40684 35080 40736 35086
rect 40684 35022 40736 35028
rect 41788 34944 41840 34950
rect 41788 34886 41840 34892
rect 41800 34678 41828 34886
rect 41788 34672 41840 34678
rect 41788 34614 41840 34620
rect 42628 33998 42656 35652
rect 42616 33992 42668 33998
rect 42616 33934 42668 33940
rect 40592 33856 40644 33862
rect 40592 33798 40644 33804
rect 40604 32910 40632 33798
rect 42156 33448 42208 33454
rect 42156 33390 42208 33396
rect 42168 32978 42196 33390
rect 42156 32972 42208 32978
rect 42156 32914 42208 32920
rect 40592 32904 40644 32910
rect 40592 32846 40644 32852
rect 41788 32836 41840 32842
rect 41788 32778 41840 32784
rect 41696 32768 41748 32774
rect 41696 32710 41748 32716
rect 41708 32502 41736 32710
rect 41696 32496 41748 32502
rect 41696 32438 41748 32444
rect 41236 32224 41288 32230
rect 41236 32166 41288 32172
rect 41248 31822 41276 32166
rect 41800 32026 41828 32778
rect 42168 32434 42196 32914
rect 42156 32428 42208 32434
rect 42156 32370 42208 32376
rect 41788 32020 41840 32026
rect 41788 31962 41840 31968
rect 42168 31890 42196 32370
rect 42156 31884 42208 31890
rect 42156 31826 42208 31832
rect 41236 31816 41288 31822
rect 41236 31758 41288 31764
rect 40500 31408 40552 31414
rect 40500 31350 40552 31356
rect 39580 31272 39632 31278
rect 39580 31214 39632 31220
rect 39304 30932 39356 30938
rect 39304 30874 39356 30880
rect 39592 30666 39620 31214
rect 39672 31136 39724 31142
rect 39672 31078 39724 31084
rect 39684 30734 39712 31078
rect 39672 30728 39724 30734
rect 39672 30670 39724 30676
rect 37740 30660 37792 30666
rect 37740 30602 37792 30608
rect 39580 30660 39632 30666
rect 39580 30602 39632 30608
rect 37752 30258 37780 30602
rect 37740 30252 37792 30258
rect 37740 30194 37792 30200
rect 38844 30252 38896 30258
rect 38844 30194 38896 30200
rect 37752 29850 37780 30194
rect 38660 30048 38712 30054
rect 38660 29990 38712 29996
rect 37740 29844 37792 29850
rect 37740 29786 37792 29792
rect 37372 28960 37424 28966
rect 37372 28902 37424 28908
rect 37384 28626 37412 28902
rect 37372 28620 37424 28626
rect 37372 28562 37424 28568
rect 38672 28150 38700 29990
rect 38856 29850 38884 30194
rect 39592 30190 39620 30602
rect 39580 30184 39632 30190
rect 39580 30126 39632 30132
rect 38844 29844 38896 29850
rect 38844 29786 38896 29792
rect 38752 29572 38804 29578
rect 38752 29514 38804 29520
rect 38764 28762 38792 29514
rect 39592 29170 39620 30126
rect 39580 29164 39632 29170
rect 39580 29106 39632 29112
rect 38936 28960 38988 28966
rect 38936 28902 38988 28908
rect 38752 28756 38804 28762
rect 38752 28698 38804 28704
rect 38948 28558 38976 28902
rect 39592 28626 39620 29106
rect 39580 28620 39632 28626
rect 39580 28562 39632 28568
rect 39948 28620 40000 28626
rect 39948 28562 40000 28568
rect 38936 28552 38988 28558
rect 38936 28494 38988 28500
rect 39960 28218 39988 28562
rect 39948 28212 40000 28218
rect 39948 28154 40000 28160
rect 38660 28144 38712 28150
rect 38660 28086 38712 28092
rect 39960 27538 39988 28154
rect 39948 27532 40000 27538
rect 39948 27474 40000 27480
rect 37280 27464 37332 27470
rect 37280 27406 37332 27412
rect 37292 27062 37320 27406
rect 39304 27328 39356 27334
rect 39304 27270 39356 27276
rect 37280 27056 37332 27062
rect 37280 26998 37332 27004
rect 37292 26382 37320 26998
rect 38660 26988 38712 26994
rect 38660 26930 38712 26936
rect 37280 26376 37332 26382
rect 37280 26318 37332 26324
rect 37292 25838 37320 26318
rect 37924 26240 37976 26246
rect 37924 26182 37976 26188
rect 37280 25832 37332 25838
rect 37280 25774 37332 25780
rect 37292 25226 37320 25774
rect 37936 25294 37964 26182
rect 38672 26042 38700 26930
rect 39028 26784 39080 26790
rect 39028 26726 39080 26732
rect 38660 26036 38712 26042
rect 38660 25978 38712 25984
rect 38660 25900 38712 25906
rect 38660 25842 38712 25848
rect 37924 25288 37976 25294
rect 37924 25230 37976 25236
rect 37280 25220 37332 25226
rect 37280 25162 37332 25168
rect 37292 24818 37320 25162
rect 37924 25152 37976 25158
rect 37924 25094 37976 25100
rect 37936 24886 37964 25094
rect 38672 24954 38700 25842
rect 38660 24948 38712 24954
rect 38660 24890 38712 24896
rect 37924 24880 37976 24886
rect 37924 24822 37976 24828
rect 37280 24812 37332 24818
rect 37280 24754 37332 24760
rect 37832 24812 37884 24818
rect 37832 24754 37884 24760
rect 38016 24812 38068 24818
rect 38016 24754 38068 24760
rect 37844 24698 37872 24754
rect 37844 24670 37964 24698
rect 37648 23656 37700 23662
rect 37648 23598 37700 23604
rect 37660 23118 37688 23598
rect 37648 23112 37700 23118
rect 37648 23054 37700 23060
rect 37372 22976 37424 22982
rect 37372 22918 37424 22924
rect 37384 22030 37412 22918
rect 37464 22636 37516 22642
rect 37464 22578 37516 22584
rect 37476 22234 37504 22578
rect 37660 22574 37688 23054
rect 37648 22568 37700 22574
rect 37648 22510 37700 22516
rect 37464 22228 37516 22234
rect 37464 22170 37516 22176
rect 37660 22098 37688 22510
rect 37648 22092 37700 22098
rect 37648 22034 37700 22040
rect 37372 22024 37424 22030
rect 37372 21966 37424 21972
rect 37556 21548 37608 21554
rect 37556 21490 37608 21496
rect 37568 21146 37596 21490
rect 37556 21140 37608 21146
rect 37556 21082 37608 21088
rect 37832 19712 37884 19718
rect 37832 19654 37884 19660
rect 37844 18766 37872 19654
rect 37832 18760 37884 18766
rect 37832 18702 37884 18708
rect 37464 18624 37516 18630
rect 37464 18566 37516 18572
rect 37096 18284 37148 18290
rect 37096 18226 37148 18232
rect 37108 17882 37136 18226
rect 37096 17876 37148 17882
rect 37096 17818 37148 17824
rect 37372 17740 37424 17746
rect 37372 17682 37424 17688
rect 37004 17332 37056 17338
rect 37004 17274 37056 17280
rect 37384 17202 37412 17682
rect 37476 17270 37504 18566
rect 37464 17264 37516 17270
rect 37464 17206 37516 17212
rect 37936 17202 37964 24670
rect 38028 24410 38056 24754
rect 38016 24404 38068 24410
rect 38016 24346 38068 24352
rect 39040 24206 39068 26726
rect 39316 26042 39344 27270
rect 39960 27062 39988 27474
rect 40408 27396 40460 27402
rect 40408 27338 40460 27344
rect 39948 27056 40000 27062
rect 39948 26998 40000 27004
rect 39856 26376 39908 26382
rect 39856 26318 39908 26324
rect 39304 26036 39356 26042
rect 39304 25978 39356 25984
rect 39868 25906 39896 26318
rect 39856 25900 39908 25906
rect 39856 25842 39908 25848
rect 39868 25294 39896 25842
rect 39856 25288 39908 25294
rect 39856 25230 39908 25236
rect 39868 24614 39896 25230
rect 40420 24682 40448 27338
rect 40512 26234 40540 31350
rect 42628 31346 42656 33934
rect 43812 33924 43864 33930
rect 43812 33866 43864 33872
rect 43824 33658 43852 33866
rect 43904 33856 43956 33862
rect 43904 33798 43956 33804
rect 43812 33652 43864 33658
rect 43812 33594 43864 33600
rect 43916 33590 43944 33798
rect 43904 33584 43956 33590
rect 43904 33526 43956 33532
rect 43812 33516 43864 33522
rect 43812 33458 43864 33464
rect 43536 32768 43588 32774
rect 43536 32710 43588 32716
rect 43548 31822 43576 32710
rect 43824 32570 43852 33458
rect 43812 32564 43864 32570
rect 43812 32506 43864 32512
rect 43628 32428 43680 32434
rect 43628 32370 43680 32376
rect 43640 32026 43668 32370
rect 43628 32020 43680 32026
rect 43628 31962 43680 31968
rect 43536 31816 43588 31822
rect 43536 31758 43588 31764
rect 44008 31482 44036 38898
rect 45204 38350 45232 38898
rect 46756 38752 46808 38758
rect 46756 38694 46808 38700
rect 46768 38350 46796 38694
rect 46860 38554 46888 41074
rect 47964 40118 47992 43658
rect 48332 43654 48360 44338
rect 48320 43648 48372 43654
rect 48320 43590 48372 43596
rect 48332 43314 48360 43590
rect 48320 43308 48372 43314
rect 48320 43250 48372 43256
rect 48332 42906 48360 43250
rect 48320 42900 48372 42906
rect 48320 42842 48372 42848
rect 48332 42226 48360 42842
rect 48884 42566 48912 44746
rect 48964 44736 49016 44742
rect 48964 44678 49016 44684
rect 48976 44470 49004 44678
rect 48964 44464 49016 44470
rect 48964 44406 49016 44412
rect 49436 44334 49464 45358
rect 51552 45082 51580 45426
rect 52736 45416 52788 45422
rect 52736 45358 52788 45364
rect 52092 45280 52144 45286
rect 52092 45222 52144 45228
rect 51540 45076 51592 45082
rect 51540 45018 51592 45024
rect 51356 44804 51408 44810
rect 51356 44746 51408 44752
rect 50294 44636 50602 44656
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44560 50602 44580
rect 49424 44328 49476 44334
rect 49424 44270 49476 44276
rect 49436 43654 49464 44270
rect 49700 44192 49752 44198
rect 49700 44134 49752 44140
rect 49608 43716 49660 43722
rect 49608 43658 49660 43664
rect 49424 43648 49476 43654
rect 49424 43590 49476 43596
rect 49436 43314 49464 43590
rect 49620 43450 49648 43658
rect 49608 43444 49660 43450
rect 49608 43386 49660 43392
rect 49712 43382 49740 44134
rect 50294 43548 50602 43568
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43472 50602 43492
rect 49700 43376 49752 43382
rect 49700 43318 49752 43324
rect 49424 43308 49476 43314
rect 49424 43250 49476 43256
rect 49436 42770 49464 43250
rect 49424 42764 49476 42770
rect 49424 42706 49476 42712
rect 51368 42566 51396 44746
rect 52104 43790 52132 45222
rect 52748 44878 52776 45358
rect 53392 45082 53420 45834
rect 53748 45824 53800 45830
rect 53748 45766 53800 45772
rect 53380 45076 53432 45082
rect 53380 45018 53432 45024
rect 52736 44872 52788 44878
rect 52736 44814 52788 44820
rect 52748 44402 52776 44814
rect 53380 44804 53432 44810
rect 53380 44746 53432 44752
rect 52736 44396 52788 44402
rect 52736 44338 52788 44344
rect 53288 44396 53340 44402
rect 53288 44338 53340 44344
rect 52092 43784 52144 43790
rect 52092 43726 52144 43732
rect 53300 43722 53328 44338
rect 53392 43994 53420 44746
rect 53760 44470 53788 45766
rect 54024 45484 54076 45490
rect 54024 45426 54076 45432
rect 54036 44538 54064 45426
rect 54576 44872 54628 44878
rect 54576 44814 54628 44820
rect 54024 44532 54076 44538
rect 54024 44474 54076 44480
rect 53748 44464 53800 44470
rect 53748 44406 53800 44412
rect 54588 44402 54616 44814
rect 55048 44470 55076 46310
rect 55324 46034 55352 46446
rect 55312 46028 55364 46034
rect 55312 45970 55364 45976
rect 55508 45626 55536 46514
rect 56704 46170 56732 46514
rect 57244 46368 57296 46374
rect 57244 46310 57296 46316
rect 56692 46164 56744 46170
rect 56692 46106 56744 46112
rect 56692 45892 56744 45898
rect 56692 45834 56744 45840
rect 55496 45620 55548 45626
rect 55496 45562 55548 45568
rect 56508 45280 56560 45286
rect 56508 45222 56560 45228
rect 56520 44946 56548 45222
rect 56704 45082 56732 45834
rect 56692 45076 56744 45082
rect 56692 45018 56744 45024
rect 56508 44940 56560 44946
rect 56508 44882 56560 44888
rect 55956 44804 56008 44810
rect 55956 44746 56008 44752
rect 55968 44538 55996 44746
rect 55956 44532 56008 44538
rect 55956 44474 56008 44480
rect 55036 44464 55088 44470
rect 55036 44406 55088 44412
rect 54576 44396 54628 44402
rect 54576 44338 54628 44344
rect 53380 43988 53432 43994
rect 53380 43930 53432 43936
rect 51632 43716 51684 43722
rect 51632 43658 51684 43664
rect 53288 43716 53340 43722
rect 53288 43658 53340 43664
rect 51540 43648 51592 43654
rect 51540 43590 51592 43596
rect 51552 43382 51580 43590
rect 51540 43376 51592 43382
rect 51540 43318 51592 43324
rect 51448 43104 51500 43110
rect 51448 43046 51500 43052
rect 51460 42702 51488 43046
rect 51448 42696 51500 42702
rect 51448 42638 51500 42644
rect 48872 42560 48924 42566
rect 48872 42502 48924 42508
rect 51356 42560 51408 42566
rect 51356 42502 51408 42508
rect 50294 42460 50602 42480
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42384 50602 42404
rect 51644 42294 51672 43658
rect 53104 43308 53156 43314
rect 53104 43250 53156 43256
rect 51632 42288 51684 42294
rect 51632 42230 51684 42236
rect 48320 42220 48372 42226
rect 48320 42162 48372 42168
rect 50160 42220 50212 42226
rect 50160 42162 50212 42168
rect 48332 41614 48360 42162
rect 49700 42016 49752 42022
rect 49700 41958 49752 41964
rect 48320 41608 48372 41614
rect 48320 41550 48372 41556
rect 48332 41138 48360 41550
rect 49332 41540 49384 41546
rect 49332 41482 49384 41488
rect 49056 41472 49108 41478
rect 49056 41414 49108 41420
rect 48320 41132 48372 41138
rect 48320 41074 48372 41080
rect 48332 40526 48360 41074
rect 48320 40520 48372 40526
rect 48320 40462 48372 40468
rect 47952 40112 48004 40118
rect 47952 40054 48004 40060
rect 47768 40044 47820 40050
rect 47768 39986 47820 39992
rect 47032 39840 47084 39846
rect 47032 39782 47084 39788
rect 47044 39030 47072 39782
rect 47780 39642 47808 39986
rect 48228 39840 48280 39846
rect 48228 39782 48280 39788
rect 47768 39636 47820 39642
rect 47768 39578 47820 39584
rect 48240 39506 48268 39782
rect 47952 39500 48004 39506
rect 47952 39442 48004 39448
rect 48228 39500 48280 39506
rect 48228 39442 48280 39448
rect 47032 39024 47084 39030
rect 47032 38966 47084 38972
rect 47964 38894 47992 39442
rect 49068 39370 49096 41414
rect 49056 39364 49108 39370
rect 49056 39306 49108 39312
rect 49344 39098 49372 41482
rect 49712 40526 49740 41958
rect 50172 41274 50200 42162
rect 51644 41614 51672 42230
rect 52184 42016 52236 42022
rect 52184 41958 52236 41964
rect 51080 41608 51132 41614
rect 51080 41550 51132 41556
rect 51632 41608 51684 41614
rect 51632 41550 51684 41556
rect 50294 41372 50602 41392
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41296 50602 41316
rect 50160 41268 50212 41274
rect 50160 41210 50212 41216
rect 51092 40934 51120 41550
rect 51540 41132 51592 41138
rect 51540 41074 51592 41080
rect 51080 40928 51132 40934
rect 51080 40870 51132 40876
rect 51092 40730 51120 40870
rect 51080 40724 51132 40730
rect 51080 40666 51132 40672
rect 49700 40520 49752 40526
rect 49700 40462 49752 40468
rect 49608 40384 49660 40390
rect 49608 40326 49660 40332
rect 49620 39438 49648 40326
rect 50294 40284 50602 40304
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40208 50602 40228
rect 51092 40118 51120 40666
rect 51552 40186 51580 41074
rect 51644 40594 51672 41550
rect 52196 41206 52224 41958
rect 52736 41608 52788 41614
rect 52736 41550 52788 41556
rect 52184 41200 52236 41206
rect 52184 41142 52236 41148
rect 52748 41070 52776 41550
rect 52920 41472 52972 41478
rect 52920 41414 52972 41420
rect 52736 41064 52788 41070
rect 52736 41006 52788 41012
rect 52184 40928 52236 40934
rect 52184 40870 52236 40876
rect 51632 40588 51684 40594
rect 51632 40530 51684 40536
rect 52196 40526 52224 40870
rect 52184 40520 52236 40526
rect 52184 40462 52236 40468
rect 51816 40384 51868 40390
rect 51816 40326 51868 40332
rect 51540 40180 51592 40186
rect 51540 40122 51592 40128
rect 49792 40112 49844 40118
rect 49792 40054 49844 40060
rect 51080 40112 51132 40118
rect 51080 40054 51132 40060
rect 49804 39846 49832 40054
rect 51828 40050 51856 40326
rect 51816 40044 51868 40050
rect 51816 39986 51868 39992
rect 49792 39840 49844 39846
rect 49792 39782 49844 39788
rect 49608 39432 49660 39438
rect 49608 39374 49660 39380
rect 49608 39296 49660 39302
rect 49608 39238 49660 39244
rect 49332 39092 49384 39098
rect 49332 39034 49384 39040
rect 49620 39030 49648 39238
rect 49608 39024 49660 39030
rect 49608 38966 49660 38972
rect 47492 38888 47544 38894
rect 47492 38830 47544 38836
rect 47952 38888 48004 38894
rect 47952 38830 48004 38836
rect 46848 38548 46900 38554
rect 46848 38490 46900 38496
rect 47504 38418 47532 38830
rect 49804 38758 49832 39782
rect 52748 39438 52776 41006
rect 52932 40526 52960 41414
rect 52920 40520 52972 40526
rect 52920 40462 52972 40468
rect 53116 39846 53144 43250
rect 53300 42770 53328 43658
rect 54588 43450 54616 44338
rect 56520 43858 56548 44882
rect 57256 44878 57284 46310
rect 57244 44872 57296 44878
rect 57244 44814 57296 44820
rect 56508 43852 56560 43858
rect 56508 43794 56560 43800
rect 54576 43444 54628 43450
rect 54576 43386 54628 43392
rect 56520 43382 56548 43794
rect 56508 43376 56560 43382
rect 56508 43318 56560 43324
rect 55588 43308 55640 43314
rect 55588 43250 55640 43256
rect 53288 42764 53340 42770
rect 53288 42706 53340 42712
rect 55128 42628 55180 42634
rect 55128 42570 55180 42576
rect 54760 42560 54812 42566
rect 54760 42502 54812 42508
rect 53656 42220 53708 42226
rect 53656 42162 53708 42168
rect 53380 42152 53432 42158
rect 53380 42094 53432 42100
rect 53392 41614 53420 42094
rect 53380 41608 53432 41614
rect 53380 41550 53432 41556
rect 53392 40594 53420 41550
rect 53668 40730 53696 42162
rect 54772 41614 54800 42502
rect 55140 42362 55168 42570
rect 55128 42356 55180 42362
rect 55128 42298 55180 42304
rect 55600 42294 55628 43250
rect 56520 42770 56548 43318
rect 57336 43104 57388 43110
rect 57336 43046 57388 43052
rect 56508 42764 56560 42770
rect 56508 42706 56560 42712
rect 56520 42362 56548 42706
rect 56508 42356 56560 42362
rect 56508 42298 56560 42304
rect 55588 42288 55640 42294
rect 55588 42230 55640 42236
rect 56232 42220 56284 42226
rect 56232 42162 56284 42168
rect 54760 41608 54812 41614
rect 54760 41550 54812 41556
rect 53748 41540 53800 41546
rect 53748 41482 53800 41488
rect 55680 41540 55732 41546
rect 55680 41482 55732 41488
rect 53760 41274 53788 41482
rect 54760 41472 54812 41478
rect 54760 41414 54812 41420
rect 53748 41268 53800 41274
rect 53748 41210 53800 41216
rect 54772 41206 54800 41414
rect 54760 41200 54812 41206
rect 54760 41142 54812 41148
rect 55692 41138 55720 41482
rect 55680 41132 55732 41138
rect 55680 41074 55732 41080
rect 55692 40730 55720 41074
rect 56244 40730 56272 42162
rect 56520 41546 56548 42298
rect 57348 41614 57376 43046
rect 57336 41608 57388 41614
rect 57336 41550 57388 41556
rect 56508 41540 56560 41546
rect 56508 41482 56560 41488
rect 57336 41472 57388 41478
rect 57336 41414 57388 41420
rect 57348 41206 57376 41414
rect 57336 41200 57388 41206
rect 57336 41142 57388 41148
rect 57060 40928 57112 40934
rect 57060 40870 57112 40876
rect 53656 40724 53708 40730
rect 53656 40666 53708 40672
rect 55680 40724 55732 40730
rect 55680 40666 55732 40672
rect 56232 40724 56284 40730
rect 56232 40666 56284 40672
rect 53380 40588 53432 40594
rect 53380 40530 53432 40536
rect 57072 40526 57100 40870
rect 57060 40520 57112 40526
rect 57060 40462 57112 40468
rect 53104 39840 53156 39846
rect 53104 39782 53156 39788
rect 54668 39840 54720 39846
rect 54668 39782 54720 39788
rect 52736 39432 52788 39438
rect 52736 39374 52788 39380
rect 53472 39432 53524 39438
rect 53472 39374 53524 39380
rect 52828 39364 52880 39370
rect 52828 39306 52880 39312
rect 53012 39364 53064 39370
rect 53012 39306 53064 39312
rect 52276 39296 52328 39302
rect 52276 39238 52328 39244
rect 50294 39196 50602 39216
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39120 50602 39140
rect 51540 39024 51592 39030
rect 51540 38966 51592 38972
rect 49792 38752 49844 38758
rect 49792 38694 49844 38700
rect 49884 38752 49936 38758
rect 49884 38694 49936 38700
rect 47492 38412 47544 38418
rect 47492 38354 47544 38360
rect 45192 38344 45244 38350
rect 45192 38286 45244 38292
rect 46756 38344 46808 38350
rect 46756 38286 46808 38292
rect 47504 38282 47532 38354
rect 44456 38276 44508 38282
rect 44456 38218 44508 38224
rect 47492 38276 47544 38282
rect 47492 38218 47544 38224
rect 44272 38208 44324 38214
rect 44272 38150 44324 38156
rect 44180 35080 44232 35086
rect 44180 35022 44232 35028
rect 44192 34678 44220 35022
rect 44180 34672 44232 34678
rect 44180 34614 44232 34620
rect 44180 33448 44232 33454
rect 44180 33390 44232 33396
rect 44192 32502 44220 33390
rect 44180 32496 44232 32502
rect 44180 32438 44232 32444
rect 43996 31476 44048 31482
rect 43996 31418 44048 31424
rect 44284 31414 44312 38150
rect 44468 38010 44496 38218
rect 47032 38208 47084 38214
rect 47032 38150 47084 38156
rect 44456 38004 44508 38010
rect 44456 37946 44508 37952
rect 44456 37868 44508 37874
rect 44456 37810 44508 37816
rect 44468 35290 44496 37810
rect 45560 37800 45612 37806
rect 45560 37742 45612 37748
rect 45572 37262 45600 37742
rect 46940 37664 46992 37670
rect 46940 37606 46992 37612
rect 45560 37256 45612 37262
rect 45560 37198 45612 37204
rect 45572 36718 45600 37198
rect 46952 36786 46980 37606
rect 47044 37262 47072 38150
rect 47504 37874 47532 38218
rect 47124 37868 47176 37874
rect 47124 37810 47176 37816
rect 47492 37868 47544 37874
rect 47492 37810 47544 37816
rect 48228 37868 48280 37874
rect 48228 37810 48280 37816
rect 47032 37256 47084 37262
rect 47032 37198 47084 37204
rect 46940 36780 46992 36786
rect 46940 36722 46992 36728
rect 45560 36712 45612 36718
rect 45560 36654 45612 36660
rect 45572 35630 45600 36654
rect 45652 36576 45704 36582
rect 45652 36518 45704 36524
rect 47032 36576 47084 36582
rect 47032 36518 47084 36524
rect 45560 35624 45612 35630
rect 45560 35566 45612 35572
rect 45572 35290 45600 35566
rect 44456 35284 44508 35290
rect 44456 35226 44508 35232
rect 45560 35284 45612 35290
rect 45560 35226 45612 35232
rect 45572 35034 45600 35226
rect 45480 35006 45600 35034
rect 45480 34542 45508 35006
rect 45664 34746 45692 36518
rect 46848 36236 46900 36242
rect 46848 36178 46900 36184
rect 46860 35222 46888 36178
rect 47044 35766 47072 36518
rect 47032 35760 47084 35766
rect 47032 35702 47084 35708
rect 47032 35488 47084 35494
rect 47032 35430 47084 35436
rect 46848 35216 46900 35222
rect 46848 35158 46900 35164
rect 47044 35086 47072 35430
rect 47136 35290 47164 37810
rect 48240 37330 48268 37810
rect 48228 37324 48280 37330
rect 48228 37266 48280 37272
rect 47768 37120 47820 37126
rect 47768 37062 47820 37068
rect 47780 36854 47808 37062
rect 47768 36848 47820 36854
rect 47768 36790 47820 36796
rect 48228 36712 48280 36718
rect 48228 36654 48280 36660
rect 48240 36242 48268 36654
rect 48228 36236 48280 36242
rect 48228 36178 48280 36184
rect 49804 36106 49832 38694
rect 49896 37942 49924 38694
rect 51552 38350 51580 38966
rect 52092 38956 52144 38962
rect 52092 38898 52144 38904
rect 51540 38344 51592 38350
rect 51540 38286 51592 38292
rect 51448 38276 51500 38282
rect 51448 38218 51500 38224
rect 50294 38108 50602 38128
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38032 50602 38052
rect 49884 37936 49936 37942
rect 49884 37878 49936 37884
rect 50804 37800 50856 37806
rect 50804 37742 50856 37748
rect 49884 37664 49936 37670
rect 49884 37606 49936 37612
rect 49896 36854 49924 37606
rect 50160 37188 50212 37194
rect 50160 37130 50212 37136
rect 50068 37120 50120 37126
rect 50068 37062 50120 37068
rect 49884 36848 49936 36854
rect 49884 36790 49936 36796
rect 50080 36106 50108 37062
rect 50172 36922 50200 37130
rect 50294 37020 50602 37040
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36944 50602 36964
rect 50160 36916 50212 36922
rect 50160 36858 50212 36864
rect 50816 36786 50844 37742
rect 50160 36780 50212 36786
rect 50160 36722 50212 36728
rect 50804 36780 50856 36786
rect 50804 36722 50856 36728
rect 50172 36174 50200 36722
rect 51460 36378 51488 38218
rect 52104 36650 52132 38898
rect 52288 37942 52316 39238
rect 52276 37936 52328 37942
rect 52276 37878 52328 37884
rect 52184 37664 52236 37670
rect 52184 37606 52236 37612
rect 52196 36854 52224 37606
rect 52840 37126 52868 39306
rect 53024 38554 53052 39306
rect 53484 38962 53512 39374
rect 53932 39296 53984 39302
rect 53932 39238 53984 39244
rect 53472 38956 53524 38962
rect 53472 38898 53524 38904
rect 53748 38752 53800 38758
rect 53748 38694 53800 38700
rect 53760 38554 53788 38694
rect 53012 38548 53064 38554
rect 53012 38490 53064 38496
rect 53748 38548 53800 38554
rect 53748 38490 53800 38496
rect 53748 38276 53800 38282
rect 53748 38218 53800 38224
rect 53760 37126 53788 38218
rect 53840 38208 53892 38214
rect 53840 38150 53892 38156
rect 53852 37194 53880 38150
rect 53840 37188 53892 37194
rect 53840 37130 53892 37136
rect 52828 37120 52880 37126
rect 52828 37062 52880 37068
rect 53564 37120 53616 37126
rect 53564 37062 53616 37068
rect 53748 37120 53800 37126
rect 53748 37062 53800 37068
rect 53576 36938 53604 37062
rect 53944 36938 53972 39238
rect 54680 37942 54708 39782
rect 56692 38956 56744 38962
rect 56692 38898 56744 38904
rect 55312 38888 55364 38894
rect 55312 38830 55364 38836
rect 54852 38752 54904 38758
rect 54852 38694 54904 38700
rect 54864 38350 54892 38694
rect 55324 38350 55352 38830
rect 56704 38554 56732 38898
rect 56692 38548 56744 38554
rect 56692 38490 56744 38496
rect 54852 38344 54904 38350
rect 54852 38286 54904 38292
rect 55312 38344 55364 38350
rect 55312 38286 55364 38292
rect 54668 37936 54720 37942
rect 54668 37878 54720 37884
rect 53576 36910 53972 36938
rect 52184 36848 52236 36854
rect 52184 36790 52236 36796
rect 52092 36644 52144 36650
rect 52092 36586 52144 36592
rect 51448 36372 51500 36378
rect 51448 36314 51500 36320
rect 50160 36168 50212 36174
rect 50160 36110 50212 36116
rect 52736 36168 52788 36174
rect 52736 36110 52788 36116
rect 49792 36100 49844 36106
rect 49792 36042 49844 36048
rect 50068 36100 50120 36106
rect 50068 36042 50120 36048
rect 47124 35284 47176 35290
rect 47124 35226 47176 35232
rect 47032 35080 47084 35086
rect 47032 35022 47084 35028
rect 46848 35012 46900 35018
rect 46848 34954 46900 34960
rect 48964 35012 49016 35018
rect 48964 34954 49016 34960
rect 46860 34746 46888 34954
rect 48976 34746 49004 34954
rect 49700 34944 49752 34950
rect 49700 34886 49752 34892
rect 45652 34740 45704 34746
rect 45652 34682 45704 34688
rect 46848 34740 46900 34746
rect 46848 34682 46900 34688
rect 48964 34740 49016 34746
rect 48964 34682 49016 34688
rect 46296 34604 46348 34610
rect 46296 34546 46348 34552
rect 48964 34604 49016 34610
rect 48964 34546 49016 34552
rect 44916 34536 44968 34542
rect 44916 34478 44968 34484
rect 45468 34536 45520 34542
rect 45468 34478 45520 34484
rect 44928 33998 44956 34478
rect 45008 34400 45060 34406
rect 45008 34342 45060 34348
rect 44916 33992 44968 33998
rect 44916 33934 44968 33940
rect 44928 31890 44956 33934
rect 45020 32502 45048 34342
rect 45560 33924 45612 33930
rect 45560 33866 45612 33872
rect 45572 32570 45600 33866
rect 45652 33312 45704 33318
rect 45652 33254 45704 33260
rect 45664 32910 45692 33254
rect 46308 33114 46336 34546
rect 47584 34536 47636 34542
rect 47584 34478 47636 34484
rect 47596 33998 47624 34478
rect 47584 33992 47636 33998
rect 47584 33934 47636 33940
rect 46388 33856 46440 33862
rect 46388 33798 46440 33804
rect 46296 33108 46348 33114
rect 46296 33050 46348 33056
rect 45652 32904 45704 32910
rect 45652 32846 45704 32852
rect 45652 32768 45704 32774
rect 45652 32710 45704 32716
rect 45560 32564 45612 32570
rect 45560 32506 45612 32512
rect 45008 32496 45060 32502
rect 45008 32438 45060 32444
rect 44916 31884 44968 31890
rect 44916 31826 44968 31832
rect 44272 31408 44324 31414
rect 44272 31350 44324 31356
rect 45664 31346 45692 32710
rect 46400 31822 46428 33798
rect 47596 33454 47624 33934
rect 48872 33924 48924 33930
rect 48872 33866 48924 33872
rect 48228 33856 48280 33862
rect 48228 33798 48280 33804
rect 48240 33590 48268 33798
rect 48228 33584 48280 33590
rect 48228 33526 48280 33532
rect 47584 33448 47636 33454
rect 47584 33390 47636 33396
rect 47596 32910 47624 33390
rect 47584 32904 47636 32910
rect 47584 32846 47636 32852
rect 46480 32836 46532 32842
rect 46480 32778 46532 32784
rect 46492 32026 46520 32778
rect 47596 32434 47624 32846
rect 48228 32768 48280 32774
rect 48228 32710 48280 32716
rect 48240 32502 48268 32710
rect 48884 32570 48912 33866
rect 48976 33658 49004 34546
rect 48964 33652 49016 33658
rect 48964 33594 49016 33600
rect 49712 33590 49740 34886
rect 49804 34678 49832 36042
rect 50172 35494 50200 36110
rect 51264 36100 51316 36106
rect 51264 36042 51316 36048
rect 50294 35932 50602 35952
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35856 50602 35876
rect 50804 35692 50856 35698
rect 50804 35634 50856 35640
rect 50160 35488 50212 35494
rect 50160 35430 50212 35436
rect 50172 35086 50200 35430
rect 50160 35080 50212 35086
rect 50160 35022 50212 35028
rect 49792 34672 49844 34678
rect 49792 34614 49844 34620
rect 50172 34406 50200 35022
rect 50294 34844 50602 34864
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34768 50602 34788
rect 50160 34400 50212 34406
rect 50160 34342 50212 34348
rect 50172 33998 50200 34342
rect 50816 34202 50844 35634
rect 51172 35488 51224 35494
rect 51172 35430 51224 35436
rect 50804 34196 50856 34202
rect 50804 34138 50856 34144
rect 50160 33992 50212 33998
rect 50160 33934 50212 33940
rect 50804 33924 50856 33930
rect 50804 33866 50856 33872
rect 51080 33924 51132 33930
rect 51080 33866 51132 33872
rect 50294 33756 50602 33776
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33680 50602 33700
rect 50816 33658 50844 33866
rect 50804 33652 50856 33658
rect 50804 33594 50856 33600
rect 49700 33584 49752 33590
rect 49700 33526 49752 33532
rect 51092 33454 51120 33866
rect 51080 33448 51132 33454
rect 51080 33390 51132 33396
rect 51092 33130 51120 33390
rect 51000 33102 51120 33130
rect 51000 32910 51028 33102
rect 51184 32910 51212 35430
rect 50804 32904 50856 32910
rect 50804 32846 50856 32852
rect 50988 32904 51040 32910
rect 50988 32846 51040 32852
rect 51172 32904 51224 32910
rect 51172 32846 51224 32852
rect 50294 32668 50602 32688
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32592 50602 32612
rect 48872 32564 48924 32570
rect 48872 32506 48924 32512
rect 48228 32496 48280 32502
rect 48228 32438 48280 32444
rect 47584 32428 47636 32434
rect 47584 32370 47636 32376
rect 46480 32020 46532 32026
rect 46480 31962 46532 31968
rect 46388 31816 46440 31822
rect 46388 31758 46440 31764
rect 47596 31346 47624 32370
rect 50816 32366 50844 32846
rect 50804 32360 50856 32366
rect 50804 32302 50856 32308
rect 50816 32026 50844 32302
rect 51080 32224 51132 32230
rect 51080 32166 51132 32172
rect 50804 32020 50856 32026
rect 50804 31962 50856 31968
rect 50816 31890 50844 31962
rect 50804 31884 50856 31890
rect 50804 31826 50856 31832
rect 50160 31816 50212 31822
rect 50160 31758 50212 31764
rect 49608 31680 49660 31686
rect 49608 31622 49660 31628
rect 40592 31340 40644 31346
rect 40592 31282 40644 31288
rect 42432 31340 42484 31346
rect 42432 31282 42484 31288
rect 42616 31340 42668 31346
rect 42616 31282 42668 31288
rect 45652 31340 45704 31346
rect 45652 31282 45704 31288
rect 46940 31340 46992 31346
rect 46940 31282 46992 31288
rect 47584 31340 47636 31346
rect 47584 31282 47636 31288
rect 40604 30394 40632 31282
rect 41696 31136 41748 31142
rect 41696 31078 41748 31084
rect 41236 30864 41288 30870
rect 41236 30806 41288 30812
rect 40592 30388 40644 30394
rect 40592 30330 40644 30336
rect 41248 30326 41276 30806
rect 41236 30320 41288 30326
rect 41236 30262 41288 30268
rect 41248 29714 41276 30262
rect 41236 29708 41288 29714
rect 41236 29650 41288 29656
rect 41512 29164 41564 29170
rect 41512 29106 41564 29112
rect 41052 29028 41104 29034
rect 41052 28970 41104 28976
rect 40684 28484 40736 28490
rect 40684 28426 40736 28432
rect 40512 26206 40632 26234
rect 40500 25696 40552 25702
rect 40500 25638 40552 25644
rect 40512 25294 40540 25638
rect 40500 25288 40552 25294
rect 40500 25230 40552 25236
rect 40408 24676 40460 24682
rect 40408 24618 40460 24624
rect 39856 24608 39908 24614
rect 39856 24550 39908 24556
rect 39868 24206 39896 24550
rect 39028 24200 39080 24206
rect 39028 24142 39080 24148
rect 39856 24200 39908 24206
rect 39856 24142 39908 24148
rect 40040 23724 40092 23730
rect 40040 23666 40092 23672
rect 38200 23520 38252 23526
rect 38200 23462 38252 23468
rect 38212 22030 38240 23462
rect 39304 23044 39356 23050
rect 39304 22986 39356 22992
rect 39316 22234 39344 22986
rect 39856 22432 39908 22438
rect 39856 22374 39908 22380
rect 39304 22228 39356 22234
rect 39304 22170 39356 22176
rect 38200 22024 38252 22030
rect 38200 21966 38252 21972
rect 39868 21622 39896 22374
rect 40052 21690 40080 23666
rect 40604 23322 40632 26206
rect 40592 23316 40644 23322
rect 40592 23258 40644 23264
rect 40604 23118 40632 23258
rect 40408 23112 40460 23118
rect 40408 23054 40460 23060
rect 40592 23112 40644 23118
rect 40592 23054 40644 23060
rect 40316 23044 40368 23050
rect 40316 22986 40368 22992
rect 40132 22976 40184 22982
rect 40132 22918 40184 22924
rect 40040 21684 40092 21690
rect 40040 21626 40092 21632
rect 39856 21616 39908 21622
rect 39856 21558 39908 21564
rect 40144 20602 40172 22918
rect 40328 22642 40356 22986
rect 40224 22636 40276 22642
rect 40224 22578 40276 22584
rect 40316 22636 40368 22642
rect 40316 22578 40368 22584
rect 40236 21146 40264 22578
rect 40328 22030 40356 22578
rect 40316 22024 40368 22030
rect 40316 21966 40368 21972
rect 40328 21554 40356 21966
rect 40316 21548 40368 21554
rect 40316 21490 40368 21496
rect 40224 21140 40276 21146
rect 40224 21082 40276 21088
rect 40328 20874 40356 21490
rect 40316 20868 40368 20874
rect 40316 20810 40368 20816
rect 40132 20596 40184 20602
rect 40132 20538 40184 20544
rect 38660 20528 38712 20534
rect 38660 20470 38712 20476
rect 38672 19854 38700 20470
rect 38752 20460 38804 20466
rect 38752 20402 38804 20408
rect 38660 19848 38712 19854
rect 38660 19790 38712 19796
rect 38672 19310 38700 19790
rect 38292 19304 38344 19310
rect 38292 19246 38344 19252
rect 38660 19304 38712 19310
rect 38660 19246 38712 19252
rect 38304 18630 38332 19246
rect 38660 19168 38712 19174
rect 38660 19110 38712 19116
rect 38292 18624 38344 18630
rect 38292 18566 38344 18572
rect 38304 18290 38332 18566
rect 38672 18358 38700 19110
rect 38660 18352 38712 18358
rect 38660 18294 38712 18300
rect 38292 18284 38344 18290
rect 38292 18226 38344 18232
rect 38304 17882 38332 18226
rect 38292 17876 38344 17882
rect 38292 17818 38344 17824
rect 38764 17338 38792 20402
rect 38844 20256 38896 20262
rect 38844 20198 38896 20204
rect 38856 17610 38884 20198
rect 39120 19780 39172 19786
rect 39120 19722 39172 19728
rect 39132 17882 39160 19722
rect 39856 19440 39908 19446
rect 39856 19382 39908 19388
rect 39868 19242 39896 19382
rect 39856 19236 39908 19242
rect 39856 19178 39908 19184
rect 39868 18834 39896 19178
rect 39856 18828 39908 18834
rect 39856 18770 39908 18776
rect 39672 18692 39724 18698
rect 39672 18634 39724 18640
rect 39304 18624 39356 18630
rect 39304 18566 39356 18572
rect 39120 17876 39172 17882
rect 39120 17818 39172 17824
rect 39316 17678 39344 18566
rect 39684 18426 39712 18634
rect 39672 18420 39724 18426
rect 39672 18362 39724 18368
rect 39868 18034 39896 18770
rect 40144 18358 40172 20538
rect 40328 20466 40356 20810
rect 40316 20460 40368 20466
rect 40316 20402 40368 20408
rect 40328 19922 40356 20402
rect 40316 19916 40368 19922
rect 40316 19858 40368 19864
rect 40132 18352 40184 18358
rect 40132 18294 40184 18300
rect 39868 18006 40080 18034
rect 39304 17672 39356 17678
rect 39304 17614 39356 17620
rect 38844 17604 38896 17610
rect 38844 17546 38896 17552
rect 38752 17332 38804 17338
rect 38752 17274 38804 17280
rect 37280 17196 37332 17202
rect 37280 17138 37332 17144
rect 37372 17196 37424 17202
rect 37372 17138 37424 17144
rect 37924 17196 37976 17202
rect 37924 17138 37976 17144
rect 37292 16794 37320 17138
rect 37280 16788 37332 16794
rect 37280 16730 37332 16736
rect 37832 16652 37884 16658
rect 37832 16594 37884 16600
rect 39764 16652 39816 16658
rect 39764 16594 39816 16600
rect 36360 16584 36412 16590
rect 36360 16526 36412 16532
rect 34796 16176 34848 16182
rect 34796 16118 34848 16124
rect 37844 16046 37872 16594
rect 39776 16182 39804 16594
rect 39856 16516 39908 16522
rect 39856 16458 39908 16464
rect 39764 16176 39816 16182
rect 39764 16118 39816 16124
rect 39028 16108 39080 16114
rect 39028 16050 39080 16056
rect 34704 16040 34756 16046
rect 34704 15982 34756 15988
rect 37832 16040 37884 16046
rect 37832 15982 37884 15988
rect 34612 15496 34664 15502
rect 34612 15438 34664 15444
rect 33968 15428 34020 15434
rect 33968 15370 34020 15376
rect 33692 15360 33744 15366
rect 33692 15302 33744 15308
rect 33232 15088 33284 15094
rect 33232 15030 33284 15036
rect 32864 14952 32916 14958
rect 32864 14894 32916 14900
rect 32876 14482 32904 14894
rect 32864 14476 32916 14482
rect 32864 14418 32916 14424
rect 32128 14408 32180 14414
rect 32128 14350 32180 14356
rect 32312 14340 32364 14346
rect 32312 14282 32364 14288
rect 30196 14068 30248 14074
rect 30196 14010 30248 14016
rect 29092 13932 29144 13938
rect 29092 13874 29144 13880
rect 28540 13184 28592 13190
rect 28540 13126 28592 13132
rect 28552 12918 28580 13126
rect 28540 12912 28592 12918
rect 28540 12854 28592 12860
rect 29000 12844 29052 12850
rect 29000 12786 29052 12792
rect 28632 12640 28684 12646
rect 28632 12582 28684 12588
rect 28644 12238 28672 12582
rect 29012 12442 29040 12786
rect 29000 12436 29052 12442
rect 29000 12378 29052 12384
rect 28632 12232 28684 12238
rect 28632 12174 28684 12180
rect 29104 11898 29132 13874
rect 30196 13728 30248 13734
rect 30196 13670 30248 13676
rect 29276 12640 29328 12646
rect 29276 12582 29328 12588
rect 29368 12640 29420 12646
rect 29368 12582 29420 12588
rect 29288 12238 29316 12582
rect 29276 12232 29328 12238
rect 29276 12174 29328 12180
rect 29092 11892 29144 11898
rect 29092 11834 29144 11840
rect 29380 11830 29408 12582
rect 30208 12238 30236 13670
rect 31944 13252 31996 13258
rect 31944 13194 31996 13200
rect 30196 12232 30248 12238
rect 30196 12174 30248 12180
rect 31116 12164 31168 12170
rect 31116 12106 31168 12112
rect 30932 12096 30984 12102
rect 30932 12038 30984 12044
rect 30944 11830 30972 12038
rect 31128 11898 31156 12106
rect 31208 12096 31260 12102
rect 31208 12038 31260 12044
rect 31116 11892 31168 11898
rect 31116 11834 31168 11840
rect 29368 11824 29420 11830
rect 29368 11766 29420 11772
rect 30932 11824 30984 11830
rect 30932 11766 30984 11772
rect 29552 11688 29604 11694
rect 29552 11630 29604 11636
rect 29564 10742 29592 11630
rect 31220 11150 31248 12038
rect 31956 11354 31984 13194
rect 32128 12844 32180 12850
rect 32128 12786 32180 12792
rect 32140 12238 32168 12786
rect 32128 12232 32180 12238
rect 32128 12174 32180 12180
rect 32140 11762 32168 12174
rect 32128 11756 32180 11762
rect 32128 11698 32180 11704
rect 31944 11348 31996 11354
rect 31944 11290 31996 11296
rect 31208 11144 31260 11150
rect 31208 11086 31260 11092
rect 32140 11082 32168 11698
rect 32128 11076 32180 11082
rect 32128 11018 32180 11024
rect 29552 10736 29604 10742
rect 29552 10678 29604 10684
rect 29564 10130 29592 10678
rect 32140 10674 32168 11018
rect 30196 10668 30248 10674
rect 30196 10610 30248 10616
rect 32128 10668 32180 10674
rect 32128 10610 32180 10616
rect 29828 10464 29880 10470
rect 29828 10406 29880 10412
rect 29552 10124 29604 10130
rect 29552 10066 29604 10072
rect 29092 9580 29144 9586
rect 29092 9522 29144 9528
rect 29000 9376 29052 9382
rect 29000 9318 29052 9324
rect 28540 8628 28592 8634
rect 28540 8570 28592 8576
rect 28552 7478 28580 8570
rect 28724 8424 28776 8430
rect 28724 8366 28776 8372
rect 28540 7472 28592 7478
rect 28540 7414 28592 7420
rect 28460 6886 28580 6914
rect 24400 6860 24452 6866
rect 24400 6802 24452 6808
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19708 6792 19760 6798
rect 19708 6734 19760 6740
rect 22008 6792 22060 6798
rect 22008 6734 22060 6740
rect 24308 6792 24360 6798
rect 24308 6734 24360 6740
rect 20904 6724 20956 6730
rect 20904 6666 20956 6672
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18708 6390 18736 6598
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 20916 6458 20944 6666
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 18696 6384 18748 6390
rect 18696 6326 18748 6332
rect 22020 6322 22048 6734
rect 23480 6724 23532 6730
rect 23480 6666 23532 6672
rect 23492 6458 23520 6666
rect 23848 6656 23900 6662
rect 23848 6598 23900 6604
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23860 6390 23888 6598
rect 23848 6384 23900 6390
rect 23848 6326 23900 6332
rect 20628 6316 20680 6322
rect 20628 6258 20680 6264
rect 22008 6316 22060 6322
rect 22008 6258 22060 6264
rect 23204 6316 23256 6322
rect 23204 6258 23256 6264
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 17132 4548 17184 4554
rect 17132 4490 17184 4496
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16316 3738 16344 4082
rect 17144 3738 17172 4490
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 17132 3732 17184 3738
rect 17132 3674 17184 3680
rect 14740 3460 14792 3466
rect 14740 3402 14792 3408
rect 14752 3194 14780 3402
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 13820 3120 13872 3126
rect 13820 3062 13872 3068
rect 16316 3058 16344 3674
rect 17328 3126 17356 4422
rect 18616 4214 18644 5170
rect 19444 4622 19472 6190
rect 20640 5914 20668 6258
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 21916 5704 21968 5710
rect 22020 5658 22048 6258
rect 23216 5914 23244 6258
rect 24320 6254 24348 6734
rect 25780 6724 25832 6730
rect 25780 6666 25832 6672
rect 25792 6458 25820 6666
rect 25780 6452 25832 6458
rect 25780 6394 25832 6400
rect 24308 6248 24360 6254
rect 24308 6190 24360 6196
rect 26976 6248 27028 6254
rect 26976 6190 27028 6196
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 26056 6112 26108 6118
rect 26056 6054 26108 6060
rect 23204 5908 23256 5914
rect 23204 5850 23256 5856
rect 24688 5710 24716 6054
rect 26068 5710 26096 6054
rect 26988 5914 27016 6190
rect 26976 5908 27028 5914
rect 26976 5850 27028 5856
rect 21968 5652 22048 5658
rect 21916 5646 22048 5652
rect 24676 5704 24728 5710
rect 24676 5646 24728 5652
rect 26056 5704 26108 5710
rect 26056 5646 26108 5652
rect 21928 5630 22048 5646
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 22020 5098 22048 5630
rect 23296 5636 23348 5642
rect 23296 5578 23348 5584
rect 22008 5092 22060 5098
rect 22008 5034 22060 5040
rect 22020 4622 22048 5034
rect 22744 5024 22796 5030
rect 22744 4966 22796 4972
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 20628 4616 20680 4622
rect 20628 4558 20680 4564
rect 22008 4616 22060 4622
rect 22008 4558 22060 4564
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 18604 4208 18656 4214
rect 18604 4150 18656 4156
rect 20640 4078 20668 4558
rect 21824 4548 21876 4554
rect 21824 4490 21876 4496
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18064 3534 18092 3878
rect 20640 3534 20668 4014
rect 21836 3738 21864 4490
rect 22020 4214 22048 4558
rect 22008 4208 22060 4214
rect 22008 4150 22060 4156
rect 22112 4146 22140 4762
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 21824 3732 21876 3738
rect 21824 3674 21876 3680
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 18144 3460 18196 3466
rect 18144 3402 18196 3408
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 17316 3120 17368 3126
rect 17316 3062 17368 3068
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 13084 2576 13136 2582
rect 13084 2518 13136 2524
rect 17236 2514 17264 2994
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 18064 2446 18092 3334
rect 18156 3194 18184 3402
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 19352 3126 19380 3470
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19340 3120 19392 3126
rect 19340 3062 19392 3068
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18616 2650 18644 2994
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 19996 2446 20024 2790
rect 20640 2446 20668 3470
rect 22756 3126 22784 4966
rect 23308 4826 23336 5578
rect 24688 5030 24716 5646
rect 25780 5296 25832 5302
rect 25780 5238 25832 5244
rect 24032 5024 24084 5030
rect 24032 4966 24084 4972
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 23296 4820 23348 4826
rect 23296 4762 23348 4768
rect 23204 4548 23256 4554
rect 23204 4490 23256 4496
rect 23216 4282 23244 4490
rect 23204 4276 23256 4282
rect 23204 4218 23256 4224
rect 24044 4078 24072 4966
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 24032 4072 24084 4078
rect 24032 4014 24084 4020
rect 23204 3460 23256 3466
rect 23204 3402 23256 3408
rect 22744 3120 22796 3126
rect 22744 3062 22796 3068
rect 23216 2650 23244 3402
rect 24044 2990 24072 4014
rect 25412 3936 25464 3942
rect 25412 3878 25464 3884
rect 24032 2984 24084 2990
rect 24032 2926 24084 2932
rect 24308 2848 24360 2854
rect 24308 2790 24360 2796
rect 23204 2644 23256 2650
rect 23204 2586 23256 2592
rect 24320 2514 24348 2790
rect 24308 2508 24360 2514
rect 24308 2450 24360 2456
rect 25424 2446 25452 3878
rect 25700 3194 25728 4082
rect 25688 3188 25740 3194
rect 25688 3130 25740 3136
rect 25792 2650 25820 5238
rect 26988 4690 27016 5850
rect 27252 5568 27304 5574
rect 27252 5510 27304 5516
rect 26976 4684 27028 4690
rect 26976 4626 27028 4632
rect 26516 4480 26568 4486
rect 26516 4422 26568 4428
rect 26528 4214 26556 4422
rect 26516 4208 26568 4214
rect 26516 4150 26568 4156
rect 26988 4146 27016 4626
rect 27264 4622 27292 5510
rect 27252 4616 27304 4622
rect 27252 4558 27304 4564
rect 26976 4140 27028 4146
rect 26976 4082 27028 4088
rect 26988 3738 27016 4082
rect 28356 3936 28408 3942
rect 28356 3878 28408 3884
rect 26976 3732 27028 3738
rect 26976 3674 27028 3680
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 26252 3126 26280 3334
rect 26240 3120 26292 3126
rect 26240 3062 26292 3068
rect 26988 2990 27016 3674
rect 28368 3534 28396 3878
rect 28356 3528 28408 3534
rect 28356 3470 28408 3476
rect 27344 3460 27396 3466
rect 27344 3402 27396 3408
rect 26976 2984 27028 2990
rect 26976 2926 27028 2932
rect 25780 2644 25832 2650
rect 25780 2586 25832 2592
rect 26988 2514 27016 2926
rect 27356 2650 27384 3402
rect 28080 3392 28132 3398
rect 28080 3334 28132 3340
rect 28092 3126 28120 3334
rect 28080 3120 28132 3126
rect 28080 3062 28132 3068
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 27344 2644 27396 2650
rect 27344 2586 27396 2592
rect 26976 2508 27028 2514
rect 26976 2450 27028 2456
rect 28368 2446 28396 2790
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 25412 2440 25464 2446
rect 25412 2382 25464 2388
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 28552 2378 28580 6886
rect 28736 6866 28764 8366
rect 29012 6914 29040 9318
rect 29104 7546 29132 9522
rect 29644 8968 29696 8974
rect 29644 8910 29696 8916
rect 29092 7540 29144 7546
rect 29092 7482 29144 7488
rect 29184 7336 29236 7342
rect 29184 7278 29236 7284
rect 28828 6886 29040 6914
rect 28724 6860 28776 6866
rect 28724 6802 28776 6808
rect 28828 6798 28856 6886
rect 29196 6798 29224 7278
rect 29656 6866 29684 8910
rect 29840 7886 29868 10406
rect 30208 9722 30236 10610
rect 30840 9988 30892 9994
rect 30840 9930 30892 9936
rect 30196 9716 30248 9722
rect 30196 9658 30248 9664
rect 30472 8900 30524 8906
rect 30472 8842 30524 8848
rect 30484 8090 30512 8842
rect 30472 8084 30524 8090
rect 30472 8026 30524 8032
rect 29828 7880 29880 7886
rect 29828 7822 29880 7828
rect 30852 7274 30880 9930
rect 32220 9920 32272 9926
rect 32220 9862 32272 9868
rect 30932 8832 30984 8838
rect 30932 8774 30984 8780
rect 30944 7478 30972 8774
rect 32232 7886 32260 9862
rect 32324 8974 32352 14282
rect 32876 14278 32904 14418
rect 32864 14272 32916 14278
rect 32864 14214 32916 14220
rect 32876 13938 32904 14214
rect 32864 13932 32916 13938
rect 32864 13874 32916 13880
rect 32876 13326 32904 13874
rect 32864 13320 32916 13326
rect 32864 13262 32916 13268
rect 32404 13184 32456 13190
rect 32404 13126 32456 13132
rect 32416 11762 32444 13126
rect 32876 12918 32904 13262
rect 32864 12912 32916 12918
rect 32864 12854 32916 12860
rect 33416 12844 33468 12850
rect 33416 12786 33468 12792
rect 33428 11898 33456 12786
rect 33508 12640 33560 12646
rect 33508 12582 33560 12588
rect 33416 11892 33468 11898
rect 33416 11834 33468 11840
rect 32404 11756 32456 11762
rect 32404 11698 32456 11704
rect 33520 11150 33548 12582
rect 33508 11144 33560 11150
rect 33508 11086 33560 11092
rect 33416 11076 33468 11082
rect 33416 11018 33468 11024
rect 33428 10606 33456 11018
rect 33704 10810 33732 15302
rect 33980 14074 34008 15370
rect 34152 15360 34204 15366
rect 34152 15302 34204 15308
rect 33968 14068 34020 14074
rect 33968 14010 34020 14016
rect 33784 13252 33836 13258
rect 33784 13194 33836 13200
rect 33796 11354 33824 13194
rect 33968 11688 34020 11694
rect 33968 11630 34020 11636
rect 33784 11348 33836 11354
rect 33784 11290 33836 11296
rect 33980 11082 34008 11630
rect 33968 11076 34020 11082
rect 33968 11018 34020 11024
rect 33692 10804 33744 10810
rect 33692 10746 33744 10752
rect 34164 10742 34192 15302
rect 34624 15026 34652 15438
rect 34520 15020 34572 15026
rect 34520 14962 34572 14968
rect 34612 15020 34664 15026
rect 34612 14962 34664 14968
rect 34532 13530 34560 14962
rect 34624 14482 34652 14962
rect 34716 14906 34744 15982
rect 36084 15904 36136 15910
rect 36084 15846 36136 15852
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 36096 15502 36124 15846
rect 37844 15586 37872 15982
rect 39040 15706 39068 16050
rect 39212 15904 39264 15910
rect 39212 15846 39264 15852
rect 39028 15700 39080 15706
rect 39028 15642 39080 15648
rect 37752 15558 37872 15586
rect 37752 15502 37780 15558
rect 36084 15496 36136 15502
rect 36084 15438 36136 15444
rect 37740 15496 37792 15502
rect 37740 15438 37792 15444
rect 36084 15360 36136 15366
rect 36084 15302 36136 15308
rect 36096 15094 36124 15302
rect 37752 15094 37780 15438
rect 38936 15428 38988 15434
rect 38936 15370 38988 15376
rect 38948 15162 38976 15370
rect 38936 15156 38988 15162
rect 38936 15098 38988 15104
rect 39224 15094 39252 15846
rect 39776 15570 39804 16118
rect 39764 15564 39816 15570
rect 39764 15506 39816 15512
rect 36084 15088 36136 15094
rect 36084 15030 36136 15036
rect 37740 15088 37792 15094
rect 37740 15030 37792 15036
rect 39212 15088 39264 15094
rect 39212 15030 39264 15036
rect 37556 15020 37608 15026
rect 37556 14962 37608 14968
rect 38936 15020 38988 15026
rect 38936 14962 38988 14968
rect 34716 14878 34836 14906
rect 34704 14816 34756 14822
rect 34704 14758 34756 14764
rect 34612 14476 34664 14482
rect 34612 14418 34664 14424
rect 34520 13524 34572 13530
rect 34520 13466 34572 13472
rect 34244 13184 34296 13190
rect 34244 13126 34296 13132
rect 34256 11762 34284 13126
rect 34716 12918 34744 14758
rect 34808 14482 34836 14878
rect 36084 14816 36136 14822
rect 36084 14758 36136 14764
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34796 14476 34848 14482
rect 34796 14418 34848 14424
rect 34808 13938 34836 14418
rect 36096 14414 36124 14758
rect 36084 14408 36136 14414
rect 36084 14350 36136 14356
rect 36268 14272 36320 14278
rect 36268 14214 36320 14220
rect 36280 14006 36308 14214
rect 36268 14000 36320 14006
rect 36268 13942 36320 13948
rect 37568 13938 37596 14962
rect 38948 14074 38976 14962
rect 39776 14482 39804 15506
rect 39868 15162 39896 16458
rect 39948 16448 40000 16454
rect 39948 16390 40000 16396
rect 39960 15502 39988 16390
rect 40052 16046 40080 18006
rect 40040 16040 40092 16046
rect 40040 15982 40092 15988
rect 39948 15496 40000 15502
rect 39948 15438 40000 15444
rect 39856 15156 39908 15162
rect 39856 15098 39908 15104
rect 40052 15026 40080 15982
rect 40040 15020 40092 15026
rect 40040 14962 40092 14968
rect 39764 14476 39816 14482
rect 39764 14418 39816 14424
rect 39856 14340 39908 14346
rect 39856 14282 39908 14288
rect 38936 14068 38988 14074
rect 38936 14010 38988 14016
rect 34796 13932 34848 13938
rect 34796 13874 34848 13880
rect 36084 13932 36136 13938
rect 36084 13874 36136 13880
rect 37556 13932 37608 13938
rect 37556 13874 37608 13880
rect 38936 13932 38988 13938
rect 38936 13874 38988 13880
rect 34808 13394 34836 13874
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34796 13388 34848 13394
rect 34796 13330 34848 13336
rect 34704 12912 34756 12918
rect 34704 12854 34756 12860
rect 34808 12850 34836 13330
rect 36096 12986 36124 13874
rect 36360 13728 36412 13734
rect 36360 13670 36412 13676
rect 36372 13326 36400 13670
rect 37568 13394 37596 13874
rect 38948 13530 38976 13874
rect 38936 13524 38988 13530
rect 38936 13466 38988 13472
rect 37556 13388 37608 13394
rect 37556 13330 37608 13336
rect 36360 13320 36412 13326
rect 36360 13262 36412 13268
rect 37568 13258 37596 13330
rect 37556 13252 37608 13258
rect 37556 13194 37608 13200
rect 38844 13252 38896 13258
rect 38844 13194 38896 13200
rect 36084 12980 36136 12986
rect 36084 12922 36136 12928
rect 37568 12850 37596 13194
rect 38856 12986 38884 13194
rect 38844 12980 38896 12986
rect 38844 12922 38896 12928
rect 34796 12844 34848 12850
rect 34796 12786 34848 12792
rect 37556 12844 37608 12850
rect 37556 12786 37608 12792
rect 38936 12844 38988 12850
rect 38936 12786 38988 12792
rect 34808 12238 34836 12786
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 37568 12306 37596 12786
rect 38948 12442 38976 12786
rect 39868 12442 39896 14282
rect 38936 12436 38988 12442
rect 38936 12378 38988 12384
rect 39856 12436 39908 12442
rect 39856 12378 39908 12384
rect 37556 12300 37608 12306
rect 37556 12242 37608 12248
rect 34796 12232 34848 12238
rect 34796 12174 34848 12180
rect 35992 12164 36044 12170
rect 35992 12106 36044 12112
rect 34244 11756 34296 11762
rect 34244 11698 34296 11704
rect 35348 11552 35400 11558
rect 35348 11494 35400 11500
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 35360 11150 35388 11494
rect 36004 11354 36032 12106
rect 36084 12096 36136 12102
rect 36084 12038 36136 12044
rect 35992 11348 36044 11354
rect 35992 11290 36044 11296
rect 35348 11144 35400 11150
rect 35348 11086 35400 11092
rect 36096 10742 36124 12038
rect 37568 11762 37596 12242
rect 38844 12164 38896 12170
rect 38844 12106 38896 12112
rect 38856 11898 38884 12106
rect 38844 11892 38896 11898
rect 38844 11834 38896 11840
rect 37556 11756 37608 11762
rect 37556 11698 37608 11704
rect 38752 11756 38804 11762
rect 38752 11698 38804 11704
rect 37568 11234 37596 11698
rect 38764 11354 38792 11698
rect 39868 11354 39896 12378
rect 40420 11558 40448 23054
rect 40696 17338 40724 28426
rect 41064 27470 41092 28970
rect 41524 28762 41552 29106
rect 41512 28756 41564 28762
rect 41512 28698 41564 28704
rect 41052 27464 41104 27470
rect 41052 27406 41104 27412
rect 41236 26988 41288 26994
rect 41236 26930 41288 26936
rect 41248 26586 41276 26930
rect 41236 26580 41288 26586
rect 41236 26522 41288 26528
rect 41144 26308 41196 26314
rect 41144 26250 41196 26256
rect 41156 24410 41184 26250
rect 41236 25152 41288 25158
rect 41236 25094 41288 25100
rect 41144 24404 41196 24410
rect 41144 24346 41196 24352
rect 41248 24206 41276 25094
rect 41420 24268 41472 24274
rect 41420 24210 41472 24216
rect 41236 24200 41288 24206
rect 41236 24142 41288 24148
rect 41432 24138 41460 24210
rect 41420 24132 41472 24138
rect 41420 24074 41472 24080
rect 41432 23526 41460 24074
rect 41708 23730 41736 31078
rect 42444 29850 42472 31282
rect 42800 30796 42852 30802
rect 42800 30738 42852 30744
rect 42616 30592 42668 30598
rect 42616 30534 42668 30540
rect 42524 30320 42576 30326
rect 42524 30262 42576 30268
rect 42432 29844 42484 29850
rect 42432 29786 42484 29792
rect 41880 29232 41932 29238
rect 41880 29174 41932 29180
rect 41892 27606 41920 29174
rect 42064 28144 42116 28150
rect 42064 28086 42116 28092
rect 41880 27600 41932 27606
rect 41880 27542 41932 27548
rect 41788 26784 41840 26790
rect 41788 26726 41840 26732
rect 41800 25294 41828 26726
rect 42076 26382 42104 28086
rect 42536 26994 42564 30262
rect 42628 29646 42656 30534
rect 42812 30326 42840 30738
rect 42984 30728 43036 30734
rect 42984 30670 43036 30676
rect 44272 30728 44324 30734
rect 44272 30670 44324 30676
rect 45652 30728 45704 30734
rect 45652 30670 45704 30676
rect 42800 30320 42852 30326
rect 42800 30262 42852 30268
rect 42996 30190 43024 30670
rect 44180 30592 44232 30598
rect 44180 30534 44232 30540
rect 42984 30184 43036 30190
rect 42984 30126 43036 30132
rect 42996 29714 43024 30126
rect 42984 29708 43036 29714
rect 42984 29650 43036 29656
rect 42616 29640 42668 29646
rect 42616 29582 42668 29588
rect 42996 29170 43024 29650
rect 42984 29164 43036 29170
rect 42984 29106 43036 29112
rect 42996 28626 43024 29106
rect 42984 28620 43036 28626
rect 42984 28562 43036 28568
rect 42996 28218 43024 28562
rect 42984 28212 43036 28218
rect 42984 28154 43036 28160
rect 42996 27538 43024 28154
rect 42984 27532 43036 27538
rect 42984 27474 43036 27480
rect 44192 27470 44220 30534
rect 44284 27606 44312 30670
rect 44364 30660 44416 30666
rect 44364 30602 44416 30608
rect 44376 28762 44404 30602
rect 45664 30190 45692 30670
rect 45652 30184 45704 30190
rect 45652 30126 45704 30132
rect 46848 30184 46900 30190
rect 46848 30126 46900 30132
rect 45100 29572 45152 29578
rect 45100 29514 45152 29520
rect 44456 29504 44508 29510
rect 44456 29446 44508 29452
rect 44364 28756 44416 28762
rect 44364 28698 44416 28704
rect 44468 28558 44496 29446
rect 44456 28552 44508 28558
rect 44456 28494 44508 28500
rect 44364 28076 44416 28082
rect 44364 28018 44416 28024
rect 44272 27600 44324 27606
rect 44272 27542 44324 27548
rect 44376 27470 44404 28018
rect 45112 27946 45140 29514
rect 45664 29306 45692 30126
rect 45836 30048 45888 30054
rect 45836 29990 45888 29996
rect 45652 29300 45704 29306
rect 45652 29242 45704 29248
rect 45664 29102 45692 29242
rect 45652 29096 45704 29102
rect 45652 29038 45704 29044
rect 45192 28960 45244 28966
rect 45192 28902 45244 28908
rect 45204 28150 45232 28902
rect 45848 28558 45876 29990
rect 46860 29850 46888 30126
rect 46848 29844 46900 29850
rect 46848 29786 46900 29792
rect 46952 29034 46980 31282
rect 47032 31136 47084 31142
rect 47032 31078 47084 31084
rect 47044 30258 47072 31078
rect 47596 30802 47624 31282
rect 47584 30796 47636 30802
rect 47584 30738 47636 30744
rect 49620 30734 49648 31622
rect 49608 30728 49660 30734
rect 49608 30670 49660 30676
rect 47124 30660 47176 30666
rect 47124 30602 47176 30608
rect 47032 30252 47084 30258
rect 47032 30194 47084 30200
rect 47032 30048 47084 30054
rect 47032 29990 47084 29996
rect 47044 29238 47072 29990
rect 47136 29850 47164 30602
rect 47768 30592 47820 30598
rect 47768 30534 47820 30540
rect 49608 30592 49660 30598
rect 49608 30534 49660 30540
rect 47780 30326 47808 30534
rect 47768 30320 47820 30326
rect 47768 30262 47820 30268
rect 47124 29844 47176 29850
rect 47124 29786 47176 29792
rect 49620 29646 49648 30534
rect 50172 30122 50200 31758
rect 50294 31580 50602 31600
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31504 50602 31524
rect 50816 31346 50844 31826
rect 50804 31340 50856 31346
rect 50804 31282 50856 31288
rect 50804 30728 50856 30734
rect 50804 30670 50856 30676
rect 50294 30492 50602 30512
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30416 50602 30436
rect 50816 30190 50844 30670
rect 51092 30326 51120 32166
rect 51276 31482 51304 36042
rect 52552 36032 52604 36038
rect 52552 35974 52604 35980
rect 51908 35012 51960 35018
rect 51908 34954 51960 34960
rect 51920 33114 51948 34954
rect 52092 34944 52144 34950
rect 52092 34886 52144 34892
rect 52104 33998 52132 34886
rect 52092 33992 52144 33998
rect 52092 33934 52144 33940
rect 51908 33108 51960 33114
rect 51908 33050 51960 33056
rect 52368 32768 52420 32774
rect 52368 32710 52420 32716
rect 52276 32428 52328 32434
rect 52276 32370 52328 32376
rect 51264 31476 51316 31482
rect 51264 31418 51316 31424
rect 52184 31340 52236 31346
rect 52184 31282 52236 31288
rect 52196 30394 52224 31282
rect 52288 30938 52316 32370
rect 52380 31822 52408 32710
rect 52368 31816 52420 31822
rect 52368 31758 52420 31764
rect 52460 31680 52512 31686
rect 52460 31622 52512 31628
rect 52276 30932 52328 30938
rect 52276 30874 52328 30880
rect 52472 30734 52500 31622
rect 52460 30728 52512 30734
rect 52460 30670 52512 30676
rect 52184 30388 52236 30394
rect 52184 30330 52236 30336
rect 51080 30320 51132 30326
rect 51080 30262 51132 30268
rect 52564 30258 52592 35974
rect 52748 35630 52776 36110
rect 53932 35692 53984 35698
rect 53932 35634 53984 35640
rect 52736 35624 52788 35630
rect 52736 35566 52788 35572
rect 52748 34542 52776 35566
rect 53012 34944 53064 34950
rect 53012 34886 53064 34892
rect 52736 34536 52788 34542
rect 52736 34478 52788 34484
rect 52748 33930 52776 34478
rect 52736 33924 52788 33930
rect 52736 33866 52788 33872
rect 52748 33454 52776 33866
rect 53024 33590 53052 34886
rect 53380 34604 53432 34610
rect 53380 34546 53432 34552
rect 53392 34202 53420 34546
rect 53380 34196 53432 34202
rect 53380 34138 53432 34144
rect 53944 33658 53972 35634
rect 54116 35488 54168 35494
rect 54116 35430 54168 35436
rect 54024 35012 54076 35018
rect 54024 34954 54076 34960
rect 54036 34542 54064 34954
rect 54128 34678 54156 35430
rect 54116 34672 54168 34678
rect 54116 34614 54168 34620
rect 54024 34536 54076 34542
rect 54024 34478 54076 34484
rect 53932 33652 53984 33658
rect 53932 33594 53984 33600
rect 54680 33590 54708 37878
rect 55324 37670 55352 38286
rect 56692 38276 56744 38282
rect 56692 38218 56744 38224
rect 55312 37664 55364 37670
rect 55312 37606 55364 37612
rect 55324 37466 55352 37606
rect 56704 37466 56732 38218
rect 55312 37460 55364 37466
rect 55312 37402 55364 37408
rect 56692 37460 56744 37466
rect 56692 37402 56744 37408
rect 55324 37262 55352 37402
rect 55312 37256 55364 37262
rect 55312 37198 55364 37204
rect 55220 36848 55272 36854
rect 55324 36802 55352 37198
rect 56416 37188 56468 37194
rect 56416 37130 56468 37136
rect 56428 36922 56456 37130
rect 56416 36916 56468 36922
rect 56416 36858 56468 36864
rect 55272 36796 55352 36802
rect 55220 36790 55352 36796
rect 55232 36774 55352 36790
rect 55324 36174 55352 36774
rect 56692 36780 56744 36786
rect 56692 36722 56744 36728
rect 56704 36378 56732 36722
rect 56692 36372 56744 36378
rect 56692 36314 56744 36320
rect 55312 36168 55364 36174
rect 55312 36110 55364 36116
rect 55324 35766 55352 36110
rect 56600 36100 56652 36106
rect 56600 36042 56652 36048
rect 55312 35760 55364 35766
rect 55312 35702 55364 35708
rect 55324 35154 55352 35702
rect 55956 35488 56008 35494
rect 55956 35430 56008 35436
rect 55312 35148 55364 35154
rect 55312 35090 55364 35096
rect 55968 35086 55996 35430
rect 55956 35080 56008 35086
rect 55956 35022 56008 35028
rect 55956 34400 56008 34406
rect 55956 34342 56008 34348
rect 53012 33584 53064 33590
rect 53012 33526 53064 33532
rect 54668 33584 54720 33590
rect 54668 33526 54720 33532
rect 52736 33448 52788 33454
rect 52736 33390 52788 33396
rect 52748 32978 52776 33390
rect 52736 32972 52788 32978
rect 52736 32914 52788 32920
rect 52748 32434 52776 32914
rect 55968 32910 55996 34342
rect 56612 34202 56640 36042
rect 56784 35692 56836 35698
rect 56784 35634 56836 35640
rect 56692 34944 56744 34950
rect 56692 34886 56744 34892
rect 56600 34196 56652 34202
rect 56600 34138 56652 34144
rect 56704 33998 56732 34886
rect 56692 33992 56744 33998
rect 56692 33934 56744 33940
rect 56796 33114 56824 35634
rect 57152 35080 57204 35086
rect 57152 35022 57204 35028
rect 56876 35012 56928 35018
rect 56876 34954 56928 34960
rect 56784 33108 56836 33114
rect 56784 33050 56836 33056
rect 55956 32904 56008 32910
rect 55956 32846 56008 32852
rect 52736 32428 52788 32434
rect 52736 32370 52788 32376
rect 52748 31890 52776 32370
rect 55496 32224 55548 32230
rect 55496 32166 55548 32172
rect 52736 31884 52788 31890
rect 52736 31826 52788 31832
rect 55508 31822 55536 32166
rect 56888 32026 56916 34954
rect 57164 34066 57192 35022
rect 57152 34060 57204 34066
rect 57152 34002 57204 34008
rect 57164 33930 57192 34002
rect 57152 33924 57204 33930
rect 57152 33866 57204 33872
rect 57164 33590 57192 33866
rect 57152 33584 57204 33590
rect 57152 33526 57204 33532
rect 57164 32978 57192 33526
rect 57152 32972 57204 32978
rect 57152 32914 57204 32920
rect 57428 32836 57480 32842
rect 57428 32778 57480 32784
rect 57440 32570 57468 32778
rect 57428 32564 57480 32570
rect 57428 32506 57480 32512
rect 56876 32020 56928 32026
rect 56876 31962 56928 31968
rect 55496 31816 55548 31822
rect 55496 31758 55548 31764
rect 57060 31748 57112 31754
rect 57060 31690 57112 31696
rect 56692 31340 56744 31346
rect 56692 31282 56744 31288
rect 52736 31272 52788 31278
rect 52736 31214 52788 31220
rect 52748 30734 52776 31214
rect 55588 31136 55640 31142
rect 55588 31078 55640 31084
rect 55600 30734 55628 31078
rect 52736 30728 52788 30734
rect 52736 30670 52788 30676
rect 55588 30728 55640 30734
rect 55588 30670 55640 30676
rect 52552 30252 52604 30258
rect 52552 30194 52604 30200
rect 52748 30190 52776 30670
rect 56600 30660 56652 30666
rect 56600 30602 56652 30608
rect 55404 30592 55456 30598
rect 55404 30534 55456 30540
rect 53012 30252 53064 30258
rect 53012 30194 53064 30200
rect 50804 30184 50856 30190
rect 50804 30126 50856 30132
rect 52736 30184 52788 30190
rect 52736 30126 52788 30132
rect 50160 30116 50212 30122
rect 50160 30058 50212 30064
rect 50816 29714 50844 30126
rect 52748 29714 52776 30126
rect 53024 29850 53052 30194
rect 54116 30048 54168 30054
rect 54116 29990 54168 29996
rect 53012 29844 53064 29850
rect 53012 29786 53064 29792
rect 50804 29708 50856 29714
rect 50804 29650 50856 29656
rect 52736 29708 52788 29714
rect 52736 29650 52788 29656
rect 49608 29640 49660 29646
rect 49608 29582 49660 29588
rect 47952 29572 48004 29578
rect 47952 29514 48004 29520
rect 47032 29232 47084 29238
rect 47032 29174 47084 29180
rect 47124 29164 47176 29170
rect 47124 29106 47176 29112
rect 46940 29028 46992 29034
rect 46940 28970 46992 28976
rect 45836 28552 45888 28558
rect 47136 28506 47164 29106
rect 45836 28494 45888 28500
rect 45652 28484 45704 28490
rect 45652 28426 45704 28432
rect 47044 28478 47164 28506
rect 45664 28218 45692 28426
rect 47044 28218 47072 28478
rect 47124 28416 47176 28422
rect 47124 28358 47176 28364
rect 45652 28212 45704 28218
rect 45652 28154 45704 28160
rect 47032 28212 47084 28218
rect 47032 28154 47084 28160
rect 45192 28144 45244 28150
rect 45192 28086 45244 28092
rect 45664 28082 45692 28154
rect 47136 28150 47164 28358
rect 47124 28144 47176 28150
rect 47124 28086 47176 28092
rect 45652 28076 45704 28082
rect 45652 28018 45704 28024
rect 45100 27940 45152 27946
rect 45100 27882 45152 27888
rect 44180 27464 44232 27470
rect 44180 27406 44232 27412
rect 44364 27464 44416 27470
rect 44364 27406 44416 27412
rect 44376 26994 44404 27406
rect 45652 27396 45704 27402
rect 45652 27338 45704 27344
rect 45664 27130 45692 27338
rect 46940 27328 46992 27334
rect 46940 27270 46992 27276
rect 45652 27124 45704 27130
rect 45652 27066 45704 27072
rect 46296 27056 46348 27062
rect 46296 26998 46348 27004
rect 42524 26988 42576 26994
rect 42524 26930 42576 26936
rect 44364 26988 44416 26994
rect 44364 26930 44416 26936
rect 42536 26586 42564 26930
rect 42524 26580 42576 26586
rect 42524 26522 42576 26528
rect 42064 26376 42116 26382
rect 42064 26318 42116 26324
rect 41788 25288 41840 25294
rect 41788 25230 41840 25236
rect 41696 23724 41748 23730
rect 41696 23666 41748 23672
rect 41420 23520 41472 23526
rect 41420 23462 41472 23468
rect 42076 22982 42104 26318
rect 42536 26234 42564 26522
rect 42444 26206 42564 26234
rect 42444 25838 42472 26206
rect 44376 25906 44404 26930
rect 44456 26784 44508 26790
rect 44456 26726 44508 26732
rect 44468 26042 44496 26726
rect 45008 26376 45060 26382
rect 45008 26318 45060 26324
rect 44456 26036 44508 26042
rect 44456 25978 44508 25984
rect 43076 25900 43128 25906
rect 43076 25842 43128 25848
rect 44364 25900 44416 25906
rect 44364 25842 44416 25848
rect 42432 25832 42484 25838
rect 42432 25774 42484 25780
rect 42444 25226 42472 25774
rect 43088 25498 43116 25842
rect 43812 25696 43864 25702
rect 43812 25638 43864 25644
rect 43076 25492 43128 25498
rect 43076 25434 43128 25440
rect 42432 25220 42484 25226
rect 42432 25162 42484 25168
rect 42444 24750 42472 25162
rect 43076 24812 43128 24818
rect 43076 24754 43128 24760
rect 42432 24744 42484 24750
rect 42432 24686 42484 24692
rect 42444 24410 42472 24686
rect 43088 24410 43116 24754
rect 42432 24404 42484 24410
rect 42432 24346 42484 24352
rect 43076 24404 43128 24410
rect 43076 24346 43128 24352
rect 43824 24206 43852 25638
rect 44376 25226 44404 25842
rect 45020 25362 45048 26318
rect 45928 26308 45980 26314
rect 45928 26250 45980 26256
rect 45652 25696 45704 25702
rect 45652 25638 45704 25644
rect 45008 25356 45060 25362
rect 45008 25298 45060 25304
rect 44364 25220 44416 25226
rect 44364 25162 44416 25168
rect 44916 25220 44968 25226
rect 44916 25162 44968 25168
rect 44928 24274 44956 25162
rect 45020 24750 45048 25298
rect 45664 25294 45692 25638
rect 45940 25498 45968 26250
rect 45928 25492 45980 25498
rect 45928 25434 45980 25440
rect 45652 25288 45704 25294
rect 45652 25230 45704 25236
rect 45008 24744 45060 24750
rect 45008 24686 45060 24692
rect 46308 24682 46336 26998
rect 46388 26988 46440 26994
rect 46388 26930 46440 26936
rect 46400 26586 46428 26930
rect 46848 26920 46900 26926
rect 46848 26862 46900 26868
rect 46388 26580 46440 26586
rect 46388 26522 46440 26528
rect 46860 26450 46888 26862
rect 46848 26444 46900 26450
rect 46848 26386 46900 26392
rect 46860 25294 46888 26386
rect 46952 25294 46980 27270
rect 47964 25906 47992 29514
rect 48320 29504 48372 29510
rect 48320 29446 48372 29452
rect 48332 29238 48360 29446
rect 50294 29404 50602 29424
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29328 50602 29348
rect 49792 29300 49844 29306
rect 49792 29242 49844 29248
rect 48320 29232 48372 29238
rect 48320 29174 48372 29180
rect 48964 29164 49016 29170
rect 48964 29106 49016 29112
rect 48976 28762 49004 29106
rect 49424 29096 49476 29102
rect 49424 29038 49476 29044
rect 48964 28756 49016 28762
rect 48964 28698 49016 28704
rect 48320 28552 48372 28558
rect 48320 28494 48372 28500
rect 48332 28150 48360 28494
rect 49056 28484 49108 28490
rect 49056 28426 49108 28432
rect 49068 28218 49096 28426
rect 49056 28212 49108 28218
rect 49056 28154 49108 28160
rect 49436 28150 49464 29038
rect 49804 28150 49832 29242
rect 50712 29028 50764 29034
rect 50712 28970 50764 28976
rect 50160 28552 50212 28558
rect 50160 28494 50212 28500
rect 48320 28144 48372 28150
rect 48320 28086 48372 28092
rect 49424 28144 49476 28150
rect 49424 28086 49476 28092
rect 49792 28144 49844 28150
rect 49792 28086 49844 28092
rect 48964 28076 49016 28082
rect 48964 28018 49016 28024
rect 48136 27396 48188 27402
rect 48136 27338 48188 27344
rect 48148 26586 48176 27338
rect 48228 27328 48280 27334
rect 48228 27270 48280 27276
rect 48240 27062 48268 27270
rect 48976 27130 49004 28018
rect 49436 28014 49464 28086
rect 49424 28008 49476 28014
rect 49424 27950 49476 27956
rect 48964 27124 49016 27130
rect 48964 27066 49016 27072
rect 48228 27056 48280 27062
rect 48228 26998 48280 27004
rect 49436 26994 49464 27950
rect 50172 27538 50200 28494
rect 50620 28416 50672 28422
rect 50620 28358 50672 28364
rect 50294 28316 50602 28336
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28240 50602 28260
rect 50160 27532 50212 27538
rect 50160 27474 50212 27480
rect 49424 26988 49476 26994
rect 49424 26930 49476 26936
rect 48136 26580 48188 26586
rect 48136 26522 48188 26528
rect 50172 26450 50200 27474
rect 50294 27228 50602 27248
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27152 50602 27172
rect 50160 26444 50212 26450
rect 50160 26386 50212 26392
rect 48136 26308 48188 26314
rect 48136 26250 48188 26256
rect 47952 25900 48004 25906
rect 47952 25842 48004 25848
rect 48148 25498 48176 26250
rect 50172 25906 50200 26386
rect 50294 26140 50602 26160
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26064 50602 26084
rect 50632 25974 50660 28358
rect 50724 27062 50752 28970
rect 50816 28558 50844 29650
rect 51816 29572 51868 29578
rect 51816 29514 51868 29520
rect 51828 29238 51856 29514
rect 51816 29232 51868 29238
rect 51816 29174 51868 29180
rect 50896 29164 50948 29170
rect 50896 29106 50948 29112
rect 50804 28552 50856 28558
rect 50804 28494 50856 28500
rect 50908 28218 50936 29106
rect 52748 28626 52776 29650
rect 54128 29238 54156 29990
rect 55416 29646 55444 30534
rect 55404 29640 55456 29646
rect 55404 29582 55456 29588
rect 54576 29572 54628 29578
rect 54576 29514 54628 29520
rect 54116 29232 54168 29238
rect 54116 29174 54168 29180
rect 53196 29028 53248 29034
rect 53196 28970 53248 28976
rect 53208 28626 53236 28970
rect 54588 28762 54616 29514
rect 56508 29504 56560 29510
rect 56508 29446 56560 29452
rect 54576 28756 54628 28762
rect 54576 28698 54628 28704
rect 52736 28620 52788 28626
rect 52736 28562 52788 28568
rect 53196 28620 53248 28626
rect 53196 28562 53248 28568
rect 51448 28484 51500 28490
rect 51448 28426 51500 28432
rect 50896 28212 50948 28218
rect 50896 28154 50948 28160
rect 50804 27396 50856 27402
rect 50804 27338 50856 27344
rect 50816 27130 50844 27338
rect 50804 27124 50856 27130
rect 50804 27066 50856 27072
rect 50712 27056 50764 27062
rect 50712 26998 50764 27004
rect 51460 26586 51488 28426
rect 53208 28082 53236 28562
rect 54760 28484 54812 28490
rect 54760 28426 54812 28432
rect 54772 28218 54800 28426
rect 54760 28212 54812 28218
rect 54760 28154 54812 28160
rect 53196 28076 53248 28082
rect 53196 28018 53248 28024
rect 54760 28076 54812 28082
rect 54760 28018 54812 28024
rect 51540 27328 51592 27334
rect 51540 27270 51592 27276
rect 51448 26580 51500 26586
rect 51448 26522 51500 26528
rect 51552 26382 51580 27270
rect 53208 26994 53236 28018
rect 54772 27606 54800 28018
rect 54760 27600 54812 27606
rect 54760 27542 54812 27548
rect 54116 27464 54168 27470
rect 54116 27406 54168 27412
rect 53196 26988 53248 26994
rect 53196 26930 53248 26936
rect 54128 26382 54156 27406
rect 54668 27396 54720 27402
rect 54668 27338 54720 27344
rect 54680 27130 54708 27338
rect 54668 27124 54720 27130
rect 54668 27066 54720 27072
rect 54760 26988 54812 26994
rect 54760 26930 54812 26936
rect 54772 26586 54800 26930
rect 54760 26580 54812 26586
rect 54760 26522 54812 26528
rect 56520 26382 56548 29446
rect 56612 29306 56640 30602
rect 56704 30394 56732 31282
rect 57072 30734 57100 31690
rect 57060 30728 57112 30734
rect 57060 30670 57112 30676
rect 56784 30660 56836 30666
rect 56784 30602 56836 30608
rect 56692 30388 56744 30394
rect 56692 30330 56744 30336
rect 56692 30252 56744 30258
rect 56692 30194 56744 30200
rect 56704 29850 56732 30194
rect 56692 29844 56744 29850
rect 56692 29786 56744 29792
rect 56600 29300 56652 29306
rect 56600 29242 56652 29248
rect 56692 28484 56744 28490
rect 56692 28426 56744 28432
rect 56600 27872 56652 27878
rect 56600 27814 56652 27820
rect 51540 26376 51592 26382
rect 51540 26318 51592 26324
rect 54116 26376 54168 26382
rect 54116 26318 54168 26324
rect 56508 26376 56560 26382
rect 56508 26318 56560 26324
rect 50620 25968 50672 25974
rect 50620 25910 50672 25916
rect 49424 25900 49476 25906
rect 49424 25842 49476 25848
rect 50160 25900 50212 25906
rect 50160 25842 50212 25848
rect 48136 25492 48188 25498
rect 48136 25434 48188 25440
rect 46848 25288 46900 25294
rect 46848 25230 46900 25236
rect 46940 25288 46992 25294
rect 46940 25230 46992 25236
rect 46860 24818 46888 25230
rect 46848 24812 46900 24818
rect 46848 24754 46900 24760
rect 48964 24812 49016 24818
rect 48964 24754 49016 24760
rect 46296 24676 46348 24682
rect 46296 24618 46348 24624
rect 45928 24608 45980 24614
rect 45928 24550 45980 24556
rect 44916 24268 44968 24274
rect 44916 24210 44968 24216
rect 43812 24200 43864 24206
rect 43812 24142 43864 24148
rect 45940 23798 45968 24550
rect 48976 24410 49004 24754
rect 48964 24404 49016 24410
rect 48964 24346 49016 24352
rect 47584 24200 47636 24206
rect 47584 24142 47636 24148
rect 48320 24200 48372 24206
rect 48320 24142 48372 24148
rect 46848 24132 46900 24138
rect 46848 24074 46900 24080
rect 46388 24064 46440 24070
rect 46388 24006 46440 24012
rect 45928 23792 45980 23798
rect 45928 23734 45980 23740
rect 44824 23724 44876 23730
rect 44824 23666 44876 23672
rect 43076 23656 43128 23662
rect 43076 23598 43128 23604
rect 43088 23118 43116 23598
rect 43076 23112 43128 23118
rect 43076 23054 43128 23060
rect 42432 23044 42484 23050
rect 42432 22986 42484 22992
rect 42064 22976 42116 22982
rect 42064 22918 42116 22924
rect 41880 22636 41932 22642
rect 41880 22578 41932 22584
rect 41696 22432 41748 22438
rect 41696 22374 41748 22380
rect 41708 20942 41736 22374
rect 41892 21690 41920 22578
rect 42076 22438 42104 22918
rect 42064 22432 42116 22438
rect 42064 22374 42116 22380
rect 42444 22234 42472 22986
rect 42616 22976 42668 22982
rect 42616 22918 42668 22924
rect 42432 22228 42484 22234
rect 42432 22170 42484 22176
rect 41880 21684 41932 21690
rect 41880 21626 41932 21632
rect 42628 21622 42656 22918
rect 43088 22642 43116 23054
rect 44180 23044 44232 23050
rect 44180 22986 44232 22992
rect 43076 22636 43128 22642
rect 43076 22578 43128 22584
rect 42800 22432 42852 22438
rect 42800 22374 42852 22380
rect 42812 21622 42840 22374
rect 44192 22234 44220 22986
rect 44456 22976 44508 22982
rect 44456 22918 44508 22924
rect 44364 22432 44416 22438
rect 44364 22374 44416 22380
rect 44180 22228 44232 22234
rect 44180 22170 44232 22176
rect 44376 22030 44404 22374
rect 44364 22024 44416 22030
rect 44364 21966 44416 21972
rect 44088 21956 44140 21962
rect 44088 21898 44140 21904
rect 42616 21616 42668 21622
rect 42616 21558 42668 21564
rect 42800 21616 42852 21622
rect 42800 21558 42852 21564
rect 42432 21344 42484 21350
rect 42432 21286 42484 21292
rect 42444 20942 42472 21286
rect 44100 21146 44128 21898
rect 44180 21548 44232 21554
rect 44180 21490 44232 21496
rect 44088 21140 44140 21146
rect 44088 21082 44140 21088
rect 41696 20936 41748 20942
rect 41696 20878 41748 20884
rect 42432 20936 42484 20942
rect 42432 20878 42484 20884
rect 41788 20460 41840 20466
rect 41788 20402 41840 20408
rect 41420 20256 41472 20262
rect 41420 20198 41472 20204
rect 41236 19372 41288 19378
rect 41236 19314 41288 19320
rect 41248 18970 41276 19314
rect 41236 18964 41288 18970
rect 41236 18906 41288 18912
rect 41432 18766 41460 20198
rect 41800 19378 41828 20402
rect 42444 20398 42472 20878
rect 44192 20602 44220 21490
rect 44468 20942 44496 22918
rect 44836 22778 44864 23666
rect 45560 23656 45612 23662
rect 45560 23598 45612 23604
rect 45192 23520 45244 23526
rect 45192 23462 45244 23468
rect 44824 22772 44876 22778
rect 44824 22714 44876 22720
rect 45204 22710 45232 23462
rect 45572 23118 45600 23598
rect 45560 23112 45612 23118
rect 45560 23054 45612 23060
rect 45192 22704 45244 22710
rect 45192 22646 45244 22652
rect 45572 22438 45600 23054
rect 46400 22642 46428 24006
rect 46860 23322 46888 24074
rect 47596 23730 47624 24142
rect 47584 23724 47636 23730
rect 47584 23666 47636 23672
rect 47032 23520 47084 23526
rect 47032 23462 47084 23468
rect 46848 23316 46900 23322
rect 46848 23258 46900 23264
rect 47044 23118 47072 23462
rect 47596 23186 47624 23666
rect 48332 23322 48360 24142
rect 48872 24132 48924 24138
rect 48872 24074 48924 24080
rect 48884 23866 48912 24074
rect 49436 24070 49464 25842
rect 54128 25838 54156 26318
rect 54760 26308 54812 26314
rect 54760 26250 54812 26256
rect 54116 25832 54168 25838
rect 54116 25774 54168 25780
rect 49516 25696 49568 25702
rect 49516 25638 49568 25644
rect 51540 25696 51592 25702
rect 51540 25638 51592 25644
rect 49528 25294 49556 25638
rect 51552 25294 51580 25638
rect 54128 25294 54156 25774
rect 54772 25498 54800 26250
rect 56520 26234 56548 26318
rect 56428 26206 56548 26234
rect 55496 25696 55548 25702
rect 55496 25638 55548 25644
rect 54760 25492 54812 25498
rect 54760 25434 54812 25440
rect 49516 25288 49568 25294
rect 49516 25230 49568 25236
rect 51540 25288 51592 25294
rect 51540 25230 51592 25236
rect 54116 25288 54168 25294
rect 54116 25230 54168 25236
rect 49528 24818 49556 25230
rect 51540 25152 51592 25158
rect 51540 25094 51592 25100
rect 50294 25052 50602 25072
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24976 50602 24996
rect 51552 24818 51580 25094
rect 49516 24812 49568 24818
rect 49516 24754 49568 24760
rect 51540 24812 51592 24818
rect 51540 24754 51592 24760
rect 49424 24064 49476 24070
rect 49424 24006 49476 24012
rect 48872 23860 48924 23866
rect 48872 23802 48924 23808
rect 49528 23730 49556 24754
rect 54128 24750 54156 25230
rect 54760 25220 54812 25226
rect 54760 25162 54812 25168
rect 54116 24744 54168 24750
rect 54116 24686 54168 24692
rect 49700 24608 49752 24614
rect 49700 24550 49752 24556
rect 49712 23798 49740 24550
rect 54128 24410 54156 24686
rect 54116 24404 54168 24410
rect 54116 24346 54168 24352
rect 50160 24200 50212 24206
rect 50160 24142 50212 24148
rect 49976 24064 50028 24070
rect 49976 24006 50028 24012
rect 49700 23792 49752 23798
rect 49700 23734 49752 23740
rect 49332 23724 49384 23730
rect 49332 23666 49384 23672
rect 49516 23724 49568 23730
rect 49516 23666 49568 23672
rect 49344 23322 49372 23666
rect 48320 23316 48372 23322
rect 48320 23258 48372 23264
rect 49332 23316 49384 23322
rect 49332 23258 49384 23264
rect 47584 23180 47636 23186
rect 47584 23122 47636 23128
rect 47032 23112 47084 23118
rect 47032 23054 47084 23060
rect 49608 23044 49660 23050
rect 49608 22986 49660 22992
rect 49620 22778 49648 22986
rect 49608 22772 49660 22778
rect 49608 22714 49660 22720
rect 46388 22636 46440 22642
rect 46388 22578 46440 22584
rect 49700 22636 49752 22642
rect 49700 22578 49752 22584
rect 45560 22432 45612 22438
rect 45560 22374 45612 22380
rect 45572 20942 45600 22374
rect 47584 21888 47636 21894
rect 47584 21830 47636 21836
rect 46388 21344 46440 21350
rect 46388 21286 46440 21292
rect 44456 20936 44508 20942
rect 44456 20878 44508 20884
rect 45560 20936 45612 20942
rect 45560 20878 45612 20884
rect 45572 20618 45600 20878
rect 44180 20596 44232 20602
rect 44180 20538 44232 20544
rect 45480 20590 45600 20618
rect 45480 20466 45508 20590
rect 43720 20460 43772 20466
rect 43720 20402 43772 20408
rect 45468 20460 45520 20466
rect 45468 20402 45520 20408
rect 42432 20392 42484 20398
rect 42432 20334 42484 20340
rect 42444 19854 42472 20334
rect 43732 20058 43760 20402
rect 45100 20392 45152 20398
rect 45100 20334 45152 20340
rect 43720 20052 43772 20058
rect 43720 19994 43772 20000
rect 45112 19854 45140 20334
rect 42432 19848 42484 19854
rect 42432 19790 42484 19796
rect 45100 19848 45152 19854
rect 45100 19790 45152 19796
rect 41880 19712 41932 19718
rect 41880 19654 41932 19660
rect 41892 19446 41920 19654
rect 41880 19440 41932 19446
rect 41880 19382 41932 19388
rect 42444 19378 42472 19790
rect 43812 19780 43864 19786
rect 43812 19722 43864 19728
rect 43824 19514 43852 19722
rect 43812 19508 43864 19514
rect 43812 19450 43864 19456
rect 41788 19372 41840 19378
rect 41788 19314 41840 19320
rect 42432 19372 42484 19378
rect 42432 19314 42484 19320
rect 43720 19372 43772 19378
rect 43720 19314 43772 19320
rect 41512 19168 41564 19174
rect 41512 19110 41564 19116
rect 41420 18760 41472 18766
rect 41420 18702 41472 18708
rect 41524 18290 41552 19110
rect 42444 18766 42472 19314
rect 43732 18970 43760 19314
rect 45112 19310 45140 19790
rect 46400 19718 46428 21286
rect 47596 20942 47624 21830
rect 49712 21690 49740 22578
rect 49988 22030 50016 24006
rect 50172 23730 50200 24142
rect 50804 24132 50856 24138
rect 50804 24074 50856 24080
rect 50294 23964 50602 23984
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23888 50602 23908
rect 50816 23866 50844 24074
rect 51540 24064 51592 24070
rect 51540 24006 51592 24012
rect 54484 24064 54536 24070
rect 54484 24006 54536 24012
rect 50804 23860 50856 23866
rect 50804 23802 50856 23808
rect 50160 23724 50212 23730
rect 50160 23666 50212 23672
rect 50172 22642 50200 23666
rect 51552 23118 51580 24006
rect 54496 23798 54524 24006
rect 54772 23866 54800 25162
rect 55508 24818 55536 25638
rect 55496 24812 55548 24818
rect 55496 24754 55548 24760
rect 54760 23860 54812 23866
rect 54760 23802 54812 23808
rect 54484 23792 54536 23798
rect 54484 23734 54536 23740
rect 53380 23724 53432 23730
rect 53380 23666 53432 23672
rect 53392 23118 53420 23666
rect 51540 23112 51592 23118
rect 51540 23054 51592 23060
rect 53380 23112 53432 23118
rect 53380 23054 53432 23060
rect 50620 23044 50672 23050
rect 50620 22986 50672 22992
rect 52092 23044 52144 23050
rect 52092 22986 52144 22992
rect 50294 22876 50602 22896
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22800 50602 22820
rect 50632 22778 50660 22986
rect 51540 22976 51592 22982
rect 51540 22918 51592 22924
rect 50620 22772 50672 22778
rect 50620 22714 50672 22720
rect 50160 22636 50212 22642
rect 50160 22578 50212 22584
rect 50632 22030 50660 22714
rect 51552 22710 51580 22918
rect 51540 22704 51592 22710
rect 51540 22646 51592 22652
rect 52000 22568 52052 22574
rect 52000 22510 52052 22516
rect 51172 22432 51224 22438
rect 51172 22374 51224 22380
rect 51184 22030 51212 22374
rect 49976 22024 50028 22030
rect 49976 21966 50028 21972
rect 50620 22024 50672 22030
rect 50620 21966 50672 21972
rect 51172 22024 51224 22030
rect 51172 21966 51224 21972
rect 49700 21684 49752 21690
rect 49700 21626 49752 21632
rect 47584 20936 47636 20942
rect 47584 20878 47636 20884
rect 46756 20868 46808 20874
rect 46756 20810 46808 20816
rect 46768 20602 46796 20810
rect 47308 20800 47360 20806
rect 47308 20742 47360 20748
rect 46756 20596 46808 20602
rect 46756 20538 46808 20544
rect 46572 20460 46624 20466
rect 46572 20402 46624 20408
rect 46584 20058 46612 20402
rect 46572 20052 46624 20058
rect 46572 19994 46624 20000
rect 47320 19854 47348 20742
rect 47596 20466 47624 20878
rect 48596 20868 48648 20874
rect 48596 20810 48648 20816
rect 47584 20460 47636 20466
rect 47584 20402 47636 20408
rect 48608 20058 48636 20810
rect 48872 20800 48924 20806
rect 48872 20742 48924 20748
rect 48596 20052 48648 20058
rect 48596 19994 48648 20000
rect 47216 19848 47268 19854
rect 47216 19790 47268 19796
rect 47308 19848 47360 19854
rect 47308 19790 47360 19796
rect 46572 19780 46624 19786
rect 46572 19722 46624 19728
rect 46388 19712 46440 19718
rect 46388 19654 46440 19660
rect 46584 19514 46612 19722
rect 46572 19508 46624 19514
rect 46572 19450 46624 19456
rect 47228 19378 47256 19790
rect 48884 19446 48912 20742
rect 49988 20534 50016 21966
rect 50988 21956 51040 21962
rect 50988 21898 51040 21904
rect 50294 21788 50602 21808
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21712 50602 21732
rect 50068 21548 50120 21554
rect 50068 21490 50120 21496
rect 50080 20924 50108 21490
rect 51000 20942 51028 21898
rect 51540 21548 51592 21554
rect 51540 21490 51592 21496
rect 51552 21146 51580 21490
rect 52012 21350 52040 22510
rect 52104 22234 52132 22986
rect 52736 22976 52788 22982
rect 52736 22918 52788 22924
rect 52092 22228 52144 22234
rect 52092 22170 52144 22176
rect 52748 22030 52776 22918
rect 55956 22636 56008 22642
rect 55956 22578 56008 22584
rect 55128 22500 55180 22506
rect 55128 22442 55180 22448
rect 52736 22024 52788 22030
rect 52736 21966 52788 21972
rect 53840 21888 53892 21894
rect 53840 21830 53892 21836
rect 53852 21622 53880 21830
rect 53840 21616 53892 21622
rect 53840 21558 53892 21564
rect 55140 21554 55168 22442
rect 55404 22432 55456 22438
rect 55404 22374 55456 22380
rect 55128 21548 55180 21554
rect 55128 21490 55180 21496
rect 52000 21344 52052 21350
rect 52000 21286 52052 21292
rect 54576 21344 54628 21350
rect 54576 21286 54628 21292
rect 51540 21140 51592 21146
rect 51540 21082 51592 21088
rect 52012 21010 52040 21286
rect 52000 21004 52052 21010
rect 52000 20946 52052 20952
rect 50160 20936 50212 20942
rect 50080 20896 50160 20924
rect 50160 20878 50212 20884
rect 50988 20936 51040 20942
rect 50988 20878 51040 20884
rect 49976 20528 50028 20534
rect 49976 20470 50028 20476
rect 48964 20460 49016 20466
rect 48964 20402 49016 20408
rect 48976 19514 49004 20402
rect 50172 19922 50200 20878
rect 50804 20868 50856 20874
rect 50804 20810 50856 20816
rect 50294 20700 50602 20720
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20624 50602 20644
rect 50252 20256 50304 20262
rect 50252 20198 50304 20204
rect 50160 19916 50212 19922
rect 50160 19858 50212 19864
rect 48964 19508 49016 19514
rect 48964 19450 49016 19456
rect 48872 19440 48924 19446
rect 48872 19382 48924 19388
rect 50172 19378 50200 19858
rect 50264 19854 50292 20198
rect 50252 19848 50304 19854
rect 50252 19790 50304 19796
rect 50294 19612 50602 19632
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19536 50602 19556
rect 50816 19514 50844 20810
rect 51000 20602 51028 20878
rect 50988 20596 51040 20602
rect 50988 20538 51040 20544
rect 52012 20398 52040 20946
rect 54588 20942 54616 21286
rect 54576 20936 54628 20942
rect 54576 20878 54628 20884
rect 55312 20936 55364 20942
rect 55312 20878 55364 20884
rect 52552 20800 52604 20806
rect 52552 20742 52604 20748
rect 52000 20392 52052 20398
rect 52000 20334 52052 20340
rect 52012 19922 52040 20334
rect 52000 19916 52052 19922
rect 52000 19858 52052 19864
rect 51540 19712 51592 19718
rect 51540 19654 51592 19660
rect 50804 19508 50856 19514
rect 50804 19450 50856 19456
rect 51552 19446 51580 19654
rect 51540 19440 51592 19446
rect 51540 19382 51592 19388
rect 46480 19372 46532 19378
rect 46480 19314 46532 19320
rect 47216 19372 47268 19378
rect 47216 19314 47268 19320
rect 50160 19372 50212 19378
rect 50160 19314 50212 19320
rect 45100 19304 45152 19310
rect 45100 19246 45152 19252
rect 43720 18964 43772 18970
rect 43720 18906 43772 18912
rect 42432 18760 42484 18766
rect 42432 18702 42484 18708
rect 45008 18760 45060 18766
rect 45008 18702 45060 18708
rect 41512 18284 41564 18290
rect 41512 18226 41564 18232
rect 42444 17882 42472 18702
rect 43812 18692 43864 18698
rect 43812 18634 43864 18640
rect 43824 18426 43852 18634
rect 43812 18420 43864 18426
rect 43812 18362 43864 18368
rect 43536 18284 43588 18290
rect 43536 18226 43588 18232
rect 43548 17882 43576 18226
rect 42432 17876 42484 17882
rect 42432 17818 42484 17824
rect 43536 17876 43588 17882
rect 43536 17818 43588 17824
rect 45020 17746 45048 18702
rect 45112 18290 45140 19246
rect 46492 18970 46520 19314
rect 46480 18964 46532 18970
rect 46480 18906 46532 18912
rect 46388 18692 46440 18698
rect 46388 18634 46440 18640
rect 46400 18426 46428 18634
rect 46388 18420 46440 18426
rect 46388 18362 46440 18368
rect 45100 18284 45152 18290
rect 45100 18226 45152 18232
rect 46388 18284 46440 18290
rect 46388 18226 46440 18232
rect 46400 17882 46428 18226
rect 46388 17876 46440 17882
rect 46388 17818 46440 17824
rect 47228 17746 47256 19314
rect 52012 18766 52040 19858
rect 52564 19854 52592 20742
rect 53380 20460 53432 20466
rect 53380 20402 53432 20408
rect 54576 20460 54628 20466
rect 54576 20402 54628 20408
rect 53392 20058 53420 20402
rect 53380 20052 53432 20058
rect 53380 19994 53432 20000
rect 54588 19854 54616 20402
rect 55324 19854 55352 20878
rect 55416 19854 55444 22374
rect 55680 22024 55732 22030
rect 55680 21966 55732 21972
rect 52552 19848 52604 19854
rect 52552 19790 52604 19796
rect 54576 19848 54628 19854
rect 54576 19790 54628 19796
rect 55312 19848 55364 19854
rect 55312 19790 55364 19796
rect 55404 19848 55456 19854
rect 55404 19790 55456 19796
rect 55692 19446 55720 21966
rect 55968 20602 55996 22578
rect 56428 22030 56456 26206
rect 56612 25974 56640 27814
rect 56600 25968 56652 25974
rect 56600 25910 56652 25916
rect 56600 25356 56652 25362
rect 56600 25298 56652 25304
rect 56612 24426 56640 25298
rect 56704 24614 56732 28426
rect 56692 24608 56744 24614
rect 56692 24550 56744 24556
rect 56520 24410 56640 24426
rect 56796 24410 56824 30602
rect 57072 30054 57100 30670
rect 57244 30592 57296 30598
rect 57244 30534 57296 30540
rect 57060 30048 57112 30054
rect 57060 29990 57112 29996
rect 57072 29646 57100 29990
rect 57256 29646 57284 30534
rect 57060 29640 57112 29646
rect 57060 29582 57112 29588
rect 57244 29640 57296 29646
rect 57244 29582 57296 29588
rect 57072 29170 57100 29582
rect 57060 29164 57112 29170
rect 57060 29106 57112 29112
rect 57072 28558 57100 29106
rect 57060 28552 57112 28558
rect 57060 28494 57112 28500
rect 57072 28150 57100 28494
rect 57060 28144 57112 28150
rect 57060 28086 57112 28092
rect 57072 27470 57100 28086
rect 57244 28076 57296 28082
rect 57244 28018 57296 28024
rect 57060 27464 57112 27470
rect 57060 27406 57112 27412
rect 57072 26994 57100 27406
rect 57256 27130 57284 28018
rect 57336 27396 57388 27402
rect 57336 27338 57388 27344
rect 57244 27124 57296 27130
rect 57244 27066 57296 27072
rect 57060 26988 57112 26994
rect 57060 26930 57112 26936
rect 57072 26518 57100 26930
rect 57060 26512 57112 26518
rect 57060 26454 57112 26460
rect 56876 25696 56928 25702
rect 56876 25638 56928 25644
rect 56888 24886 56916 25638
rect 57072 25498 57100 26454
rect 57348 26042 57376 27338
rect 57336 26036 57388 26042
rect 57336 25978 57388 25984
rect 57060 25492 57112 25498
rect 57060 25434 57112 25440
rect 57336 25220 57388 25226
rect 57336 25162 57388 25168
rect 57348 24954 57376 25162
rect 57336 24948 57388 24954
rect 57336 24890 57388 24896
rect 56876 24880 56928 24886
rect 56876 24822 56928 24828
rect 56508 24404 56640 24410
rect 56560 24398 56640 24404
rect 56784 24404 56836 24410
rect 56508 24346 56560 24352
rect 56784 24346 56836 24352
rect 56888 24290 56916 24822
rect 57336 24812 57388 24818
rect 57336 24754 57388 24760
rect 56796 24262 56916 24290
rect 56796 24138 56824 24262
rect 56784 24132 56836 24138
rect 56784 24074 56836 24080
rect 57244 24132 57296 24138
rect 57244 24074 57296 24080
rect 56796 23730 56824 24074
rect 56784 23724 56836 23730
rect 56784 23666 56836 23672
rect 56796 23118 56824 23666
rect 56784 23112 56836 23118
rect 56784 23054 56836 23060
rect 56796 22438 56824 23054
rect 57256 22778 57284 24074
rect 57348 23866 57376 24754
rect 57336 23860 57388 23866
rect 57336 23802 57388 23808
rect 57244 22772 57296 22778
rect 57244 22714 57296 22720
rect 56784 22432 56836 22438
rect 56784 22374 56836 22380
rect 56416 22024 56468 22030
rect 56416 21966 56468 21972
rect 56796 21894 56824 22374
rect 56784 21888 56836 21894
rect 56784 21830 56836 21836
rect 56692 21548 56744 21554
rect 56692 21490 56744 21496
rect 56704 21146 56732 21490
rect 56692 21140 56744 21146
rect 56692 21082 56744 21088
rect 56796 20942 56824 21830
rect 57244 21344 57296 21350
rect 57244 21286 57296 21292
rect 56784 20936 56836 20942
rect 56784 20878 56836 20884
rect 56692 20868 56744 20874
rect 56692 20810 56744 20816
rect 55956 20596 56008 20602
rect 55956 20538 56008 20544
rect 56704 20058 56732 20810
rect 56692 20052 56744 20058
rect 56692 19994 56744 20000
rect 56796 19938 56824 20878
rect 56704 19910 56824 19938
rect 55864 19848 55916 19854
rect 55864 19790 55916 19796
rect 55876 19446 55904 19790
rect 55680 19440 55732 19446
rect 55680 19382 55732 19388
rect 55864 19440 55916 19446
rect 55864 19382 55916 19388
rect 56704 18766 56732 19910
rect 57256 19854 57284 21286
rect 57244 19848 57296 19854
rect 57244 19790 57296 19796
rect 52000 18760 52052 18766
rect 52000 18702 52052 18708
rect 56692 18760 56744 18766
rect 56692 18702 56744 18708
rect 51816 18624 51868 18630
rect 51816 18566 51868 18572
rect 50294 18524 50602 18544
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18448 50602 18468
rect 51264 18352 51316 18358
rect 51264 18294 51316 18300
rect 50620 18080 50672 18086
rect 50620 18022 50672 18028
rect 45008 17740 45060 17746
rect 45008 17682 45060 17688
rect 47216 17740 47268 17746
rect 47216 17682 47268 17688
rect 43812 17604 43864 17610
rect 43812 17546 43864 17552
rect 43824 17338 43852 17546
rect 40684 17332 40736 17338
rect 40684 17274 40736 17280
rect 43812 17332 43864 17338
rect 43812 17274 43864 17280
rect 45020 17202 45048 17682
rect 46296 17604 46348 17610
rect 46296 17546 46348 17552
rect 46308 17338 46336 17546
rect 46296 17332 46348 17338
rect 46296 17274 46348 17280
rect 47228 17202 47256 17682
rect 48780 17604 48832 17610
rect 48780 17546 48832 17552
rect 43904 17196 43956 17202
rect 43904 17138 43956 17144
rect 45008 17196 45060 17202
rect 45008 17138 45060 17144
rect 46388 17196 46440 17202
rect 46388 17138 46440 17144
rect 47216 17196 47268 17202
rect 47216 17138 47268 17144
rect 42432 17128 42484 17134
rect 42432 17070 42484 17076
rect 42444 16658 42472 17070
rect 43916 16794 43944 17138
rect 43904 16788 43956 16794
rect 43904 16730 43956 16736
rect 42432 16652 42484 16658
rect 42432 16594 42484 16600
rect 42064 16448 42116 16454
rect 42064 16390 42116 16396
rect 42076 16182 42104 16390
rect 42064 16176 42116 16182
rect 42064 16118 42116 16124
rect 42444 16114 42472 16594
rect 45020 16590 45048 17138
rect 46400 16794 46428 17138
rect 48792 16794 48820 17546
rect 49056 17536 49108 17542
rect 49056 17478 49108 17484
rect 46388 16788 46440 16794
rect 46388 16730 46440 16736
rect 48780 16788 48832 16794
rect 48780 16730 48832 16736
rect 47400 16652 47452 16658
rect 47400 16594 47452 16600
rect 45008 16584 45060 16590
rect 45008 16526 45060 16532
rect 47412 16538 47440 16594
rect 42616 16516 42668 16522
rect 42616 16458 42668 16464
rect 43812 16516 43864 16522
rect 43812 16458 43864 16464
rect 41236 16108 41288 16114
rect 41236 16050 41288 16056
rect 42432 16108 42484 16114
rect 42432 16050 42484 16056
rect 41248 15706 41276 16050
rect 41512 15904 41564 15910
rect 41512 15846 41564 15852
rect 41236 15700 41288 15706
rect 41236 15642 41288 15648
rect 41524 14414 41552 15846
rect 42628 15706 42656 16458
rect 43824 16250 43852 16458
rect 43812 16244 43864 16250
rect 43812 16186 43864 16192
rect 45020 16114 45048 16526
rect 46388 16516 46440 16522
rect 47412 16510 47624 16538
rect 46388 16458 46440 16464
rect 46400 16250 46428 16458
rect 46388 16244 46440 16250
rect 46388 16186 46440 16192
rect 45008 16108 45060 16114
rect 45008 16050 45060 16056
rect 46388 16108 46440 16114
rect 46388 16050 46440 16056
rect 46400 15706 46428 16050
rect 47596 16046 47624 16510
rect 49068 16182 49096 17478
rect 50294 17436 50602 17456
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17360 50602 17380
rect 49332 16992 49384 16998
rect 49332 16934 49384 16940
rect 49344 16590 49372 16934
rect 49332 16584 49384 16590
rect 49332 16526 49384 16532
rect 50294 16348 50602 16368
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16272 50602 16292
rect 50632 16182 50660 18022
rect 51276 17746 51304 18294
rect 51264 17740 51316 17746
rect 51264 17682 51316 17688
rect 50804 17264 50856 17270
rect 50804 17206 50856 17212
rect 50816 17134 50844 17206
rect 50896 17196 50948 17202
rect 50896 17138 50948 17144
rect 50804 17128 50856 17134
rect 50804 17070 50856 17076
rect 50908 16250 50936 17138
rect 51828 16590 51856 18566
rect 52012 18358 52040 18702
rect 52644 18692 52696 18698
rect 52644 18634 52696 18640
rect 52000 18352 52052 18358
rect 52000 18294 52052 18300
rect 52184 18284 52236 18290
rect 52184 18226 52236 18232
rect 52196 17338 52224 18226
rect 52656 17882 52684 18634
rect 56704 18290 56732 18702
rect 57244 18692 57296 18698
rect 57244 18634 57296 18640
rect 54760 18284 54812 18290
rect 54760 18226 54812 18232
rect 56692 18284 56744 18290
rect 56692 18226 56744 18232
rect 53840 18216 53892 18222
rect 53840 18158 53892 18164
rect 53852 17882 53880 18158
rect 54300 18080 54352 18086
rect 54300 18022 54352 18028
rect 52644 17876 52696 17882
rect 52644 17818 52696 17824
rect 53840 17876 53892 17882
rect 53840 17818 53892 17824
rect 52184 17332 52236 17338
rect 52184 17274 52236 17280
rect 53852 17202 53880 17818
rect 54312 17678 54340 18022
rect 54300 17672 54352 17678
rect 54300 17614 54352 17620
rect 52920 17196 52972 17202
rect 52920 17138 52972 17144
rect 53840 17196 53892 17202
rect 53840 17138 53892 17144
rect 52932 16794 52960 17138
rect 52920 16788 52972 16794
rect 52920 16730 52972 16736
rect 51540 16584 51592 16590
rect 51540 16526 51592 16532
rect 51816 16584 51868 16590
rect 51816 16526 51868 16532
rect 50896 16244 50948 16250
rect 50896 16186 50948 16192
rect 49056 16176 49108 16182
rect 49056 16118 49108 16124
rect 50620 16176 50672 16182
rect 50620 16118 50672 16124
rect 51552 16114 51580 16526
rect 54772 16454 54800 18226
rect 55864 18080 55916 18086
rect 55864 18022 55916 18028
rect 55876 17270 55904 18022
rect 55956 17672 56008 17678
rect 55956 17614 56008 17620
rect 55864 17264 55916 17270
rect 55864 17206 55916 17212
rect 55968 17202 55996 17614
rect 57256 17338 57284 18634
rect 57336 17604 57388 17610
rect 57336 17546 57388 17552
rect 57244 17332 57296 17338
rect 57244 17274 57296 17280
rect 55956 17196 56008 17202
rect 55956 17138 56008 17144
rect 55496 16992 55548 16998
rect 55496 16934 55548 16940
rect 55404 16516 55456 16522
rect 55404 16458 55456 16464
rect 54760 16448 54812 16454
rect 54760 16390 54812 16396
rect 51540 16108 51592 16114
rect 51540 16050 51592 16056
rect 52000 16108 52052 16114
rect 52000 16050 52052 16056
rect 47584 16040 47636 16046
rect 47584 15982 47636 15988
rect 42616 15700 42668 15706
rect 42616 15642 42668 15648
rect 46388 15700 46440 15706
rect 46388 15642 46440 15648
rect 45008 15496 45060 15502
rect 45008 15438 45060 15444
rect 41604 15428 41656 15434
rect 41604 15370 41656 15376
rect 41616 14618 41644 15370
rect 41604 14612 41656 14618
rect 41604 14554 41656 14560
rect 45020 14482 45048 15438
rect 46388 15428 46440 15434
rect 46388 15370 46440 15376
rect 46400 15162 46428 15370
rect 47596 15366 47624 15982
rect 49056 15904 49108 15910
rect 49056 15846 49108 15852
rect 48136 15564 48188 15570
rect 48136 15506 48188 15512
rect 47584 15360 47636 15366
rect 47584 15302 47636 15308
rect 46388 15156 46440 15162
rect 46388 15098 46440 15104
rect 45560 15088 45612 15094
rect 45560 15030 45612 15036
rect 45008 14476 45060 14482
rect 45008 14418 45060 14424
rect 41512 14408 41564 14414
rect 41512 14350 41564 14356
rect 45020 14090 45048 14418
rect 44548 14068 44600 14074
rect 44548 14010 44600 14016
rect 44928 14062 45048 14090
rect 42984 13932 43036 13938
rect 42984 13874 43036 13880
rect 42996 13530 43024 13874
rect 44272 13728 44324 13734
rect 44272 13670 44324 13676
rect 42984 13524 43036 13530
rect 42984 13466 43036 13472
rect 42524 13320 42576 13326
rect 42524 13262 42576 13268
rect 41696 12436 41748 12442
rect 41696 12378 41748 12384
rect 40500 12232 40552 12238
rect 40500 12174 40552 12180
rect 40512 11762 40540 12174
rect 40500 11756 40552 11762
rect 40500 11698 40552 11704
rect 40408 11552 40460 11558
rect 40408 11494 40460 11500
rect 38752 11348 38804 11354
rect 38752 11290 38804 11296
rect 39856 11348 39908 11354
rect 39856 11290 39908 11296
rect 37476 11206 37596 11234
rect 37476 11150 37504 11206
rect 37464 11144 37516 11150
rect 37464 11086 37516 11092
rect 34152 10736 34204 10742
rect 34152 10678 34204 10684
rect 36084 10736 36136 10742
rect 36084 10678 36136 10684
rect 33416 10600 33468 10606
rect 33416 10542 33468 10548
rect 37280 10600 37332 10606
rect 37280 10542 37332 10548
rect 33428 10062 33456 10542
rect 35624 10464 35676 10470
rect 35624 10406 35676 10412
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 33416 10056 33468 10062
rect 33416 9998 33468 10004
rect 33428 9518 33456 9998
rect 34060 9988 34112 9994
rect 34060 9930 34112 9936
rect 33416 9512 33468 9518
rect 33416 9454 33468 9460
rect 32312 8968 32364 8974
rect 32312 8910 32364 8916
rect 33428 8838 33456 9454
rect 34072 9382 34100 9930
rect 34152 9920 34204 9926
rect 34152 9862 34204 9868
rect 34060 9376 34112 9382
rect 34060 9318 34112 9324
rect 33416 8832 33468 8838
rect 33416 8774 33468 8780
rect 33428 8430 33456 8774
rect 34164 8566 34192 9862
rect 35636 9654 35664 10406
rect 35624 9648 35676 9654
rect 35624 9590 35676 9596
rect 37292 9586 37320 10542
rect 37476 10266 37504 11086
rect 38660 11076 38712 11082
rect 38660 11018 38712 11024
rect 38672 10810 38700 11018
rect 38660 10804 38712 10810
rect 38660 10746 38712 10752
rect 38568 10668 38620 10674
rect 38568 10610 38620 10616
rect 38580 10266 38608 10610
rect 37464 10260 37516 10266
rect 37464 10202 37516 10208
rect 38568 10260 38620 10266
rect 38568 10202 38620 10208
rect 38660 9988 38712 9994
rect 38660 9930 38712 9936
rect 38672 9722 38700 9930
rect 38660 9716 38712 9722
rect 38660 9658 38712 9664
rect 37280 9580 37332 9586
rect 37280 9522 37332 9528
rect 37372 9580 37424 9586
rect 37372 9522 37424 9528
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34428 8968 34480 8974
rect 34428 8910 34480 8916
rect 35808 8968 35860 8974
rect 35808 8910 35860 8916
rect 34152 8560 34204 8566
rect 34152 8502 34204 8508
rect 34440 8498 34468 8910
rect 34796 8900 34848 8906
rect 34796 8842 34848 8848
rect 34808 8634 34836 8842
rect 34796 8628 34848 8634
rect 34796 8570 34848 8576
rect 34428 8492 34480 8498
rect 34428 8434 34480 8440
rect 33416 8424 33468 8430
rect 33416 8366 33468 8372
rect 32128 7880 32180 7886
rect 32128 7822 32180 7828
rect 32220 7880 32272 7886
rect 32220 7822 32272 7828
rect 30932 7472 30984 7478
rect 30932 7414 30984 7420
rect 32140 7342 32168 7822
rect 33428 7818 33456 8366
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 35820 7818 35848 8910
rect 36636 8900 36688 8906
rect 36636 8842 36688 8848
rect 36084 8832 36136 8838
rect 36084 8774 36136 8780
rect 35992 8492 36044 8498
rect 35992 8434 36044 8440
rect 36004 8090 36032 8434
rect 35992 8084 36044 8090
rect 35992 8026 36044 8032
rect 36096 7886 36124 8774
rect 36648 8634 36676 8842
rect 36636 8628 36688 8634
rect 36636 8570 36688 8576
rect 37292 8498 37320 9522
rect 37280 8492 37332 8498
rect 37280 8434 37332 8440
rect 36084 7880 36136 7886
rect 36084 7822 36136 7828
rect 33416 7812 33468 7818
rect 33416 7754 33468 7760
rect 35808 7812 35860 7818
rect 35808 7754 35860 7760
rect 33508 7744 33560 7750
rect 33508 7686 33560 7692
rect 33520 7478 33548 7686
rect 35820 7478 35848 7754
rect 37384 7546 37412 9522
rect 37924 8832 37976 8838
rect 37924 8774 37976 8780
rect 37936 8566 37964 8774
rect 37924 8560 37976 8566
rect 37924 8502 37976 8508
rect 38844 8492 38896 8498
rect 38844 8434 38896 8440
rect 38660 8288 38712 8294
rect 38660 8230 38712 8236
rect 38672 7886 38700 8230
rect 38856 8090 38884 8434
rect 38844 8084 38896 8090
rect 38844 8026 38896 8032
rect 38660 7880 38712 7886
rect 38660 7822 38712 7828
rect 37372 7540 37424 7546
rect 37372 7482 37424 7488
rect 33508 7472 33560 7478
rect 33508 7414 33560 7420
rect 35808 7472 35860 7478
rect 35808 7414 35860 7420
rect 35348 7404 35400 7410
rect 35348 7346 35400 7352
rect 39212 7404 39264 7410
rect 39212 7346 39264 7352
rect 32128 7336 32180 7342
rect 32128 7278 32180 7284
rect 30840 7268 30892 7274
rect 30840 7210 30892 7216
rect 32140 6866 32168 7278
rect 32312 7200 32364 7206
rect 32312 7142 32364 7148
rect 29644 6860 29696 6866
rect 29644 6802 29696 6808
rect 32128 6860 32180 6866
rect 32128 6802 32180 6808
rect 28816 6792 28868 6798
rect 28816 6734 28868 6740
rect 29184 6792 29236 6798
rect 29184 6734 29236 6740
rect 29000 6656 29052 6662
rect 29000 6598 29052 6604
rect 28908 6316 28960 6322
rect 28908 6258 28960 6264
rect 28920 5914 28948 6258
rect 28908 5908 28960 5914
rect 28908 5850 28960 5856
rect 29012 5710 29040 6598
rect 29196 5778 29224 6734
rect 29656 6322 29684 6802
rect 30288 6792 30340 6798
rect 30288 6734 30340 6740
rect 30300 6390 30328 6734
rect 31024 6724 31076 6730
rect 31024 6666 31076 6672
rect 30288 6384 30340 6390
rect 30288 6326 30340 6332
rect 29644 6316 29696 6322
rect 29644 6258 29696 6264
rect 30932 6316 30984 6322
rect 30932 6258 30984 6264
rect 29656 5794 29684 6258
rect 30944 5914 30972 6258
rect 29736 5908 29788 5914
rect 29736 5850 29788 5856
rect 30932 5908 30984 5914
rect 30932 5850 30984 5856
rect 29748 5794 29776 5850
rect 29184 5772 29236 5778
rect 29656 5766 29776 5794
rect 29184 5714 29236 5720
rect 29000 5704 29052 5710
rect 29000 5646 29052 5652
rect 29196 4690 29224 5714
rect 29644 5636 29696 5642
rect 29644 5578 29696 5584
rect 29184 4684 29236 4690
rect 29184 4626 29236 4632
rect 29656 3194 29684 5578
rect 29748 5302 29776 5766
rect 29736 5296 29788 5302
rect 29736 5238 29788 5244
rect 29748 3534 29776 5238
rect 31036 3738 31064 6666
rect 32140 6254 32168 6802
rect 32324 6798 32352 7142
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 32312 6792 32364 6798
rect 32312 6734 32364 6740
rect 34060 6656 34112 6662
rect 34060 6598 34112 6604
rect 34072 6390 34100 6598
rect 34060 6384 34112 6390
rect 34060 6326 34112 6332
rect 35360 6254 35388 7346
rect 38660 7336 38712 7342
rect 38660 7278 38712 7284
rect 38672 6798 38700 7278
rect 39224 7002 39252 7346
rect 39212 6996 39264 7002
rect 39212 6938 39264 6944
rect 35808 6792 35860 6798
rect 35808 6734 35860 6740
rect 37740 6792 37792 6798
rect 37740 6734 37792 6740
rect 38660 6792 38712 6798
rect 38660 6734 38712 6740
rect 32128 6248 32180 6254
rect 32128 6190 32180 6196
rect 35348 6248 35400 6254
rect 35348 6190 35400 6196
rect 31116 6112 31168 6118
rect 31116 6054 31168 6060
rect 31128 4622 31156 6054
rect 32140 5778 32168 6190
rect 33508 6112 33560 6118
rect 33508 6054 33560 6060
rect 32128 5772 32180 5778
rect 32128 5714 32180 5720
rect 33520 5710 33548 6054
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 35360 5914 35388 6190
rect 35820 5914 35848 6734
rect 36728 6724 36780 6730
rect 36728 6666 36780 6672
rect 36740 6458 36768 6666
rect 36728 6452 36780 6458
rect 36728 6394 36780 6400
rect 36728 6316 36780 6322
rect 36728 6258 36780 6264
rect 35348 5908 35400 5914
rect 35348 5850 35400 5856
rect 35808 5908 35860 5914
rect 35808 5850 35860 5856
rect 33508 5704 33560 5710
rect 33508 5646 33560 5652
rect 34060 5568 34112 5574
rect 34060 5510 34112 5516
rect 34072 5302 34100 5510
rect 34060 5296 34112 5302
rect 34060 5238 34112 5244
rect 32588 5228 32640 5234
rect 32588 5170 32640 5176
rect 32600 4622 32628 5170
rect 34612 5160 34664 5166
rect 34612 5102 34664 5108
rect 33876 5024 33928 5030
rect 33876 4966 33928 4972
rect 33888 4622 33916 4966
rect 34624 4622 34652 5102
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 31116 4616 31168 4622
rect 31116 4558 31168 4564
rect 32588 4616 32640 4622
rect 32588 4558 32640 4564
rect 33876 4616 33928 4622
rect 33876 4558 33928 4564
rect 34612 4616 34664 4622
rect 34612 4558 34664 4564
rect 31392 4480 31444 4486
rect 31392 4422 31444 4428
rect 31404 4146 31432 4422
rect 31392 4140 31444 4146
rect 31392 4082 31444 4088
rect 32600 4078 32628 4558
rect 34152 4480 34204 4486
rect 34152 4422 34204 4428
rect 34164 4146 34192 4422
rect 34152 4140 34204 4146
rect 34152 4082 34204 4088
rect 34624 4078 34652 4558
rect 35820 4554 35848 5850
rect 35992 5568 36044 5574
rect 35992 5510 36044 5516
rect 35808 4548 35860 4554
rect 35808 4490 35860 4496
rect 32588 4072 32640 4078
rect 32588 4014 32640 4020
rect 34612 4072 34664 4078
rect 34612 4014 34664 4020
rect 31116 3936 31168 3942
rect 31116 3878 31168 3884
rect 31024 3732 31076 3738
rect 31024 3674 31076 3680
rect 31128 3534 31156 3878
rect 32600 3602 32628 4014
rect 34624 3602 34652 4014
rect 36004 4010 36032 5510
rect 36544 5024 36596 5030
rect 36544 4966 36596 4972
rect 36556 4622 36584 4966
rect 36740 4826 36768 6258
rect 37752 6254 37780 6734
rect 37740 6248 37792 6254
rect 37740 6190 37792 6196
rect 37752 5710 37780 6190
rect 39396 6112 39448 6118
rect 39396 6054 39448 6060
rect 39408 5914 39436 6054
rect 39396 5908 39448 5914
rect 39396 5850 39448 5856
rect 37740 5704 37792 5710
rect 37740 5646 37792 5652
rect 37752 5166 37780 5646
rect 39212 5568 39264 5574
rect 39212 5510 39264 5516
rect 39224 5302 39252 5510
rect 39868 5302 39896 11290
rect 40420 11150 40448 11494
rect 40512 11218 40540 11698
rect 40500 11212 40552 11218
rect 40500 11154 40552 11160
rect 40408 11144 40460 11150
rect 40408 11086 40460 11092
rect 40512 10674 40540 11154
rect 40500 10668 40552 10674
rect 40500 10610 40552 10616
rect 40500 9580 40552 9586
rect 40500 9522 40552 9528
rect 40512 9042 40540 9522
rect 40500 9036 40552 9042
rect 40500 8978 40552 8984
rect 40512 8430 40540 8978
rect 41420 8492 41472 8498
rect 41420 8434 41472 8440
rect 40500 8424 40552 8430
rect 40420 8372 40500 8378
rect 40420 8366 40552 8372
rect 40420 8350 40540 8366
rect 40420 7342 40448 8350
rect 40500 8288 40552 8294
rect 40500 8230 40552 8236
rect 40512 7478 40540 8230
rect 41432 7546 41460 8434
rect 41708 7886 41736 12378
rect 42536 12238 42564 13262
rect 43904 13252 43956 13258
rect 43904 13194 43956 13200
rect 43168 12844 43220 12850
rect 43168 12786 43220 12792
rect 43180 12442 43208 12786
rect 43916 12442 43944 13194
rect 43168 12436 43220 12442
rect 43168 12378 43220 12384
rect 43904 12436 43956 12442
rect 43904 12378 43956 12384
rect 42524 12232 42576 12238
rect 42524 12174 42576 12180
rect 41880 12164 41932 12170
rect 41880 12106 41932 12112
rect 41892 11898 41920 12106
rect 41880 11892 41932 11898
rect 41880 11834 41932 11840
rect 42536 11762 42564 12174
rect 44284 11830 44312 13670
rect 44560 11830 44588 14010
rect 44928 14006 44956 14062
rect 44916 14000 44968 14006
rect 44916 13942 44968 13948
rect 44928 12918 44956 13942
rect 45572 13326 45600 15030
rect 46664 15020 46716 15026
rect 46664 14962 46716 14968
rect 46676 14618 46704 14962
rect 47596 14958 47624 15302
rect 47584 14952 47636 14958
rect 47584 14894 47636 14900
rect 46664 14612 46716 14618
rect 46664 14554 46716 14560
rect 47596 14414 47624 14894
rect 47584 14408 47636 14414
rect 47584 14350 47636 14356
rect 46388 14340 46440 14346
rect 46388 14282 46440 14288
rect 46400 13530 46428 14282
rect 46756 13932 46808 13938
rect 46756 13874 46808 13880
rect 46388 13524 46440 13530
rect 46388 13466 46440 13472
rect 45560 13320 45612 13326
rect 45560 13262 45612 13268
rect 44916 12912 44968 12918
rect 44916 12854 44968 12860
rect 44272 11824 44324 11830
rect 44272 11766 44324 11772
rect 44548 11824 44600 11830
rect 44548 11766 44600 11772
rect 44928 11762 44956 12854
rect 45572 12306 45600 13262
rect 45744 13252 45796 13258
rect 45744 13194 45796 13200
rect 45652 12844 45704 12850
rect 45652 12786 45704 12792
rect 45560 12300 45612 12306
rect 45560 12242 45612 12248
rect 45664 11914 45692 12786
rect 45480 11898 45692 11914
rect 45756 11898 45784 13194
rect 46768 12986 46796 13874
rect 47596 13870 47624 14350
rect 47584 13864 47636 13870
rect 47584 13806 47636 13812
rect 47952 13728 48004 13734
rect 47952 13670 48004 13676
rect 47964 13326 47992 13670
rect 47952 13320 48004 13326
rect 47952 13262 48004 13268
rect 46756 12980 46808 12986
rect 46756 12922 46808 12928
rect 45836 12300 45888 12306
rect 45836 12242 45888 12248
rect 45468 11892 45692 11898
rect 45520 11886 45692 11892
rect 45744 11892 45796 11898
rect 45468 11834 45520 11840
rect 45744 11834 45796 11840
rect 41880 11756 41932 11762
rect 41880 11698 41932 11704
rect 42524 11756 42576 11762
rect 42524 11698 42576 11704
rect 44916 11756 44968 11762
rect 44916 11698 44968 11704
rect 41892 11354 41920 11698
rect 41880 11348 41932 11354
rect 41880 11290 41932 11296
rect 45848 11082 45876 12242
rect 47768 12096 47820 12102
rect 47768 12038 47820 12044
rect 47780 11150 47808 12038
rect 47964 11354 47992 13262
rect 47952 11348 48004 11354
rect 47952 11290 48004 11296
rect 47768 11144 47820 11150
rect 47768 11086 47820 11092
rect 41788 11076 41840 11082
rect 41788 11018 41840 11024
rect 45836 11076 45888 11082
rect 45836 11018 45888 11024
rect 41800 10810 41828 11018
rect 41788 10804 41840 10810
rect 41788 10746 41840 10752
rect 45848 10690 45876 11018
rect 47768 11008 47820 11014
rect 47768 10950 47820 10956
rect 47780 10742 47808 10950
rect 48148 10810 48176 15506
rect 49068 15094 49096 15846
rect 52012 15502 52040 16050
rect 55416 15978 55444 16458
rect 55508 16182 55536 16934
rect 55956 16584 56008 16590
rect 55956 16526 56008 16532
rect 55496 16176 55548 16182
rect 55496 16118 55548 16124
rect 55968 16046 55996 16526
rect 57348 16250 57376 17546
rect 57336 16244 57388 16250
rect 57336 16186 57388 16192
rect 55956 16040 56008 16046
rect 55956 15982 56008 15988
rect 55404 15972 55456 15978
rect 55404 15914 55456 15920
rect 55968 15502 55996 15982
rect 52000 15496 52052 15502
rect 52000 15438 52052 15444
rect 55956 15496 56008 15502
rect 55956 15438 56008 15444
rect 56416 15496 56468 15502
rect 56416 15438 56468 15444
rect 51448 15428 51500 15434
rect 51448 15370 51500 15376
rect 49516 15360 49568 15366
rect 49516 15302 49568 15308
rect 49056 15088 49108 15094
rect 49056 15030 49108 15036
rect 49148 15020 49200 15026
rect 49148 14962 49200 14968
rect 49056 14816 49108 14822
rect 49056 14758 49108 14764
rect 49068 14414 49096 14758
rect 49056 14408 49108 14414
rect 49056 14350 49108 14356
rect 48964 14272 49016 14278
rect 48964 14214 49016 14220
rect 48976 14006 49004 14214
rect 49160 14074 49188 14962
rect 49528 14958 49556 15302
rect 50294 15260 50602 15280
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15184 50602 15204
rect 49516 14952 49568 14958
rect 49516 14894 49568 14900
rect 49148 14068 49200 14074
rect 49148 14010 49200 14016
rect 48964 14000 49016 14006
rect 48964 13942 49016 13948
rect 49528 13938 49556 14894
rect 49792 14816 49844 14822
rect 49792 14758 49844 14764
rect 49700 14340 49752 14346
rect 49700 14282 49752 14288
rect 49516 13932 49568 13938
rect 49516 13874 49568 13880
rect 49712 13530 49740 14282
rect 49700 13524 49752 13530
rect 49700 13466 49752 13472
rect 49804 13326 49832 14758
rect 50294 14172 50602 14192
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14096 50602 14116
rect 51172 13728 51224 13734
rect 51172 13670 51224 13676
rect 51184 13326 51212 13670
rect 51460 13530 51488 15370
rect 52012 15026 52040 15438
rect 53288 15428 53340 15434
rect 53288 15370 53340 15376
rect 52092 15360 52144 15366
rect 52092 15302 52144 15308
rect 53104 15360 53156 15366
rect 53104 15302 53156 15308
rect 52000 15020 52052 15026
rect 52000 14962 52052 14968
rect 52012 14482 52040 14962
rect 52000 14476 52052 14482
rect 52000 14418 52052 14424
rect 51540 14272 51592 14278
rect 51540 14214 51592 14220
rect 51552 14006 51580 14214
rect 51540 14000 51592 14006
rect 51540 13942 51592 13948
rect 51448 13524 51500 13530
rect 51448 13466 51500 13472
rect 52012 13394 52040 14418
rect 52104 14414 52132 15302
rect 52092 14408 52144 14414
rect 52092 14350 52144 14356
rect 53116 13938 53144 15302
rect 53104 13932 53156 13938
rect 53104 13874 53156 13880
rect 53300 13530 53328 15370
rect 53748 15360 53800 15366
rect 53748 15302 53800 15308
rect 53656 14816 53708 14822
rect 53656 14758 53708 14764
rect 53380 14272 53432 14278
rect 53380 14214 53432 14220
rect 53288 13524 53340 13530
rect 53288 13466 53340 13472
rect 52000 13388 52052 13394
rect 52000 13330 52052 13336
rect 49792 13320 49844 13326
rect 49792 13262 49844 13268
rect 51172 13320 51224 13326
rect 51172 13262 51224 13268
rect 51172 13184 51224 13190
rect 51172 13126 51224 13132
rect 50294 13084 50602 13104
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13008 50602 13028
rect 48228 12844 48280 12850
rect 48228 12786 48280 12792
rect 50620 12844 50672 12850
rect 50620 12786 50672 12792
rect 48240 12306 48268 12786
rect 50068 12640 50120 12646
rect 50068 12582 50120 12588
rect 48228 12300 48280 12306
rect 48228 12242 48280 12248
rect 49608 11756 49660 11762
rect 49608 11698 49660 11704
rect 48596 11688 48648 11694
rect 48596 11630 48648 11636
rect 48412 11552 48464 11558
rect 48412 11494 48464 11500
rect 48136 10804 48188 10810
rect 48136 10746 48188 10752
rect 45756 10674 45876 10690
rect 47768 10736 47820 10742
rect 47768 10678 47820 10684
rect 41880 10668 41932 10674
rect 41880 10610 41932 10616
rect 45744 10668 45876 10674
rect 45796 10662 45876 10668
rect 45744 10610 45796 10616
rect 41892 9722 41920 10610
rect 43352 10464 43404 10470
rect 43352 10406 43404 10412
rect 43364 9994 43392 10406
rect 45756 10062 45784 10610
rect 47860 10260 47912 10266
rect 47860 10202 47912 10208
rect 45744 10056 45796 10062
rect 45744 9998 45796 10004
rect 43352 9988 43404 9994
rect 43352 9930 43404 9936
rect 45652 9988 45704 9994
rect 45652 9930 45704 9936
rect 45376 9920 45428 9926
rect 45376 9862 45428 9868
rect 41880 9716 41932 9722
rect 41880 9658 41932 9664
rect 42064 9580 42116 9586
rect 42064 9522 42116 9528
rect 43904 9580 43956 9586
rect 43904 9522 43956 9528
rect 42076 9178 42104 9522
rect 43812 9376 43864 9382
rect 43812 9318 43864 9324
rect 42064 9172 42116 9178
rect 42064 9114 42116 9120
rect 41880 8900 41932 8906
rect 41880 8842 41932 8848
rect 41972 8900 42024 8906
rect 41972 8842 42024 8848
rect 41696 7880 41748 7886
rect 41696 7822 41748 7828
rect 41892 7546 41920 8842
rect 41420 7540 41472 7546
rect 41420 7482 41472 7488
rect 41880 7540 41932 7546
rect 41880 7482 41932 7488
rect 40500 7472 40552 7478
rect 40500 7414 40552 7420
rect 40408 7336 40460 7342
rect 40460 7296 40632 7324
rect 40408 7278 40460 7284
rect 40604 6866 40632 7296
rect 40592 6860 40644 6866
rect 40592 6802 40644 6808
rect 40604 6118 40632 6802
rect 41984 6662 42012 8842
rect 43628 8356 43680 8362
rect 43628 8298 43680 8304
rect 42800 8288 42852 8294
rect 42800 8230 42852 8236
rect 42812 8090 42840 8230
rect 42800 8084 42852 8090
rect 42800 8026 42852 8032
rect 42812 7342 42840 8026
rect 43536 7404 43588 7410
rect 43536 7346 43588 7352
rect 42800 7336 42852 7342
rect 42800 7278 42852 7284
rect 41972 6656 42024 6662
rect 41972 6598 42024 6604
rect 41696 6316 41748 6322
rect 41696 6258 41748 6264
rect 40224 6112 40276 6118
rect 40224 6054 40276 6060
rect 40592 6112 40644 6118
rect 40592 6054 40644 6060
rect 40236 5778 40264 6054
rect 41708 5914 41736 6258
rect 41512 5908 41564 5914
rect 41512 5850 41564 5856
rect 41696 5908 41748 5914
rect 41696 5850 41748 5856
rect 40224 5772 40276 5778
rect 40224 5714 40276 5720
rect 41236 5636 41288 5642
rect 41236 5578 41288 5584
rect 39212 5296 39264 5302
rect 39212 5238 39264 5244
rect 39856 5296 39908 5302
rect 39856 5238 39908 5244
rect 39488 5228 39540 5234
rect 39488 5170 39540 5176
rect 37740 5160 37792 5166
rect 37740 5102 37792 5108
rect 36728 4820 36780 4826
rect 36728 4762 36780 4768
rect 36544 4616 36596 4622
rect 36544 4558 36596 4564
rect 37752 4214 37780 5102
rect 38844 4548 38896 4554
rect 38844 4490 38896 4496
rect 38568 4480 38620 4486
rect 38568 4422 38620 4428
rect 37740 4208 37792 4214
rect 37740 4150 37792 4156
rect 37280 4140 37332 4146
rect 37280 4082 37332 4088
rect 35992 4004 36044 4010
rect 35992 3946 36044 3952
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 32588 3596 32640 3602
rect 32588 3538 32640 3544
rect 34612 3596 34664 3602
rect 34612 3538 34664 3544
rect 29736 3528 29788 3534
rect 29736 3470 29788 3476
rect 31116 3528 31168 3534
rect 31116 3470 31168 3476
rect 29644 3188 29696 3194
rect 29644 3130 29696 3136
rect 32600 3058 32628 3538
rect 33508 3460 33560 3466
rect 33508 3402 33560 3408
rect 34060 3460 34112 3466
rect 34060 3402 34112 3408
rect 32588 3052 32640 3058
rect 32588 2994 32640 3000
rect 33520 2650 33548 3402
rect 33968 3392 34020 3398
rect 33968 3334 34020 3340
rect 33980 3126 34008 3334
rect 34072 3194 34100 3402
rect 34060 3188 34112 3194
rect 34060 3130 34112 3136
rect 33968 3120 34020 3126
rect 33968 3062 34020 3068
rect 34624 3058 34652 3538
rect 35900 3460 35952 3466
rect 35900 3402 35952 3408
rect 35912 3194 35940 3402
rect 36084 3392 36136 3398
rect 36084 3334 36136 3340
rect 36452 3392 36504 3398
rect 36452 3334 36504 3340
rect 35900 3188 35952 3194
rect 35900 3130 35952 3136
rect 36096 3126 36124 3334
rect 36084 3120 36136 3126
rect 36084 3062 36136 3068
rect 34612 3052 34664 3058
rect 34612 2994 34664 3000
rect 33508 2644 33560 2650
rect 33508 2586 33560 2592
rect 34624 2514 34652 2994
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 34612 2508 34664 2514
rect 34612 2450 34664 2456
rect 36464 2446 36492 3334
rect 37292 3058 37320 4082
rect 37280 3052 37332 3058
rect 37280 2994 37332 3000
rect 37556 3052 37608 3058
rect 37556 2994 37608 3000
rect 37292 2514 37320 2994
rect 37568 2650 37596 2994
rect 37556 2644 37608 2650
rect 37556 2586 37608 2592
rect 37280 2508 37332 2514
rect 37280 2450 37332 2456
rect 38580 2446 38608 4422
rect 38752 4140 38804 4146
rect 38752 4082 38804 4088
rect 38660 3936 38712 3942
rect 38660 3878 38712 3884
rect 38672 3126 38700 3878
rect 38660 3120 38712 3126
rect 38660 3062 38712 3068
rect 38764 2650 38792 4082
rect 38856 2922 38884 4490
rect 39500 3738 39528 5170
rect 39948 5024 40000 5030
rect 39948 4966 40000 4972
rect 39960 4622 39988 4966
rect 41248 4826 41276 5578
rect 41236 4820 41288 4826
rect 41236 4762 41288 4768
rect 39856 4616 39908 4622
rect 39856 4558 39908 4564
rect 39948 4616 40000 4622
rect 39948 4558 40000 4564
rect 39868 4214 39896 4558
rect 41524 4554 41552 5850
rect 42812 5710 42840 7278
rect 43076 6792 43128 6798
rect 43076 6734 43128 6740
rect 43088 6322 43116 6734
rect 43076 6316 43128 6322
rect 43076 6258 43128 6264
rect 43352 6112 43404 6118
rect 43352 6054 43404 6060
rect 43364 5710 43392 6054
rect 42800 5704 42852 5710
rect 42800 5646 42852 5652
rect 43352 5704 43404 5710
rect 43352 5646 43404 5652
rect 42708 5568 42760 5574
rect 42708 5510 42760 5516
rect 41696 5160 41748 5166
rect 41696 5102 41748 5108
rect 41708 4622 41736 5102
rect 41696 4616 41748 4622
rect 41696 4558 41748 4564
rect 42432 4616 42484 4622
rect 42432 4558 42484 4564
rect 41512 4548 41564 4554
rect 41512 4490 41564 4496
rect 39856 4208 39908 4214
rect 39856 4150 39908 4156
rect 39488 3732 39540 3738
rect 39488 3674 39540 3680
rect 39868 3602 39896 4150
rect 40408 4140 40460 4146
rect 40408 4082 40460 4088
rect 39856 3596 39908 3602
rect 39856 3538 39908 3544
rect 39868 3058 39896 3538
rect 40420 3194 40448 4082
rect 42444 4078 42472 4558
rect 42432 4072 42484 4078
rect 42432 4014 42484 4020
rect 40500 3936 40552 3942
rect 40500 3878 40552 3884
rect 40512 3534 40540 3878
rect 40500 3528 40552 3534
rect 40500 3470 40552 3476
rect 40408 3188 40460 3194
rect 40408 3130 40460 3136
rect 42444 3058 42472 4014
rect 42720 3126 42748 5510
rect 42812 3738 42840 5646
rect 43076 4480 43128 4486
rect 43076 4422 43128 4428
rect 42800 3732 42852 3738
rect 42800 3674 42852 3680
rect 43088 3534 43116 4422
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 43548 3194 43576 7346
rect 43640 6798 43668 8298
rect 43824 7478 43852 9318
rect 43916 9178 43944 9522
rect 43904 9172 43956 9178
rect 43904 9114 43956 9120
rect 44180 8900 44232 8906
rect 44180 8842 44232 8848
rect 44192 7546 44220 8842
rect 45388 7818 45416 9862
rect 45664 9722 45692 9930
rect 45652 9716 45704 9722
rect 45652 9658 45704 9664
rect 45652 9580 45704 9586
rect 45652 9522 45704 9528
rect 45664 8634 45692 9522
rect 45756 8974 45784 9998
rect 45744 8968 45796 8974
rect 45744 8910 45796 8916
rect 46848 8968 46900 8974
rect 46848 8910 46900 8916
rect 45652 8628 45704 8634
rect 45652 8570 45704 8576
rect 45756 8498 45784 8910
rect 46388 8832 46440 8838
rect 46388 8774 46440 8780
rect 46400 8566 46428 8774
rect 46388 8560 46440 8566
rect 46388 8502 46440 8508
rect 46860 8498 46888 8910
rect 47124 8900 47176 8906
rect 47124 8842 47176 8848
rect 45744 8492 45796 8498
rect 45744 8434 45796 8440
rect 46848 8492 46900 8498
rect 46848 8434 46900 8440
rect 45756 7886 45784 8434
rect 46860 7954 46888 8434
rect 47136 8090 47164 8842
rect 47400 8832 47452 8838
rect 47400 8774 47452 8780
rect 47124 8084 47176 8090
rect 47124 8026 47176 8032
rect 46848 7948 46900 7954
rect 46848 7890 46900 7896
rect 45744 7880 45796 7886
rect 45744 7822 45796 7828
rect 45376 7812 45428 7818
rect 45376 7754 45428 7760
rect 44180 7540 44232 7546
rect 44180 7482 44232 7488
rect 43812 7472 43864 7478
rect 43812 7414 43864 7420
rect 46860 7342 46888 7890
rect 47412 7886 47440 8774
rect 47400 7880 47452 7886
rect 47400 7822 47452 7828
rect 47124 7404 47176 7410
rect 47124 7346 47176 7352
rect 45652 7336 45704 7342
rect 45652 7278 45704 7284
rect 46848 7336 46900 7342
rect 46848 7278 46900 7284
rect 45664 6798 45692 7278
rect 47136 7002 47164 7346
rect 47492 7336 47544 7342
rect 47492 7278 47544 7284
rect 47124 6996 47176 7002
rect 47124 6938 47176 6944
rect 47504 6798 47532 7278
rect 47676 7200 47728 7206
rect 47676 7142 47728 7148
rect 43628 6792 43680 6798
rect 43628 6734 43680 6740
rect 43904 6792 43956 6798
rect 43904 6734 43956 6740
rect 45652 6792 45704 6798
rect 45652 6734 45704 6740
rect 47492 6792 47544 6798
rect 47492 6734 47544 6740
rect 43916 6322 43944 6734
rect 45284 6724 45336 6730
rect 45284 6666 45336 6672
rect 44456 6656 44508 6662
rect 44456 6598 44508 6604
rect 43904 6316 43956 6322
rect 43904 6258 43956 6264
rect 43916 5710 43944 6258
rect 43904 5704 43956 5710
rect 43904 5646 43956 5652
rect 43812 5636 43864 5642
rect 43812 5578 43864 5584
rect 43824 3738 43852 5578
rect 43916 5234 43944 5646
rect 44272 5568 44324 5574
rect 44272 5510 44324 5516
rect 43904 5228 43956 5234
rect 43904 5170 43956 5176
rect 44284 4146 44312 5510
rect 44468 5370 44496 6598
rect 44456 5364 44508 5370
rect 44456 5306 44508 5312
rect 44272 4140 44324 4146
rect 44272 4082 44324 4088
rect 45296 4010 45324 6666
rect 47504 6322 47532 6734
rect 45376 6316 45428 6322
rect 45376 6258 45428 6264
rect 47400 6316 47452 6322
rect 47400 6258 47452 6264
rect 47492 6316 47544 6322
rect 47492 6258 47544 6264
rect 45388 5370 45416 6258
rect 46848 6112 46900 6118
rect 46848 6054 46900 6060
rect 47032 6112 47084 6118
rect 47032 6054 47084 6060
rect 46388 5568 46440 5574
rect 46388 5510 46440 5516
rect 45376 5364 45428 5370
rect 45376 5306 45428 5312
rect 46400 5302 46428 5510
rect 46388 5296 46440 5302
rect 46388 5238 46440 5244
rect 46860 4162 46888 6054
rect 46860 4134 46980 4162
rect 47044 4146 47072 6054
rect 47412 4826 47440 6258
rect 47400 4820 47452 4826
rect 47400 4762 47452 4768
rect 47688 4622 47716 7142
rect 47872 6798 47900 10202
rect 48148 10062 48176 10746
rect 48424 10674 48452 11494
rect 48608 11082 48636 11630
rect 49620 11354 49648 11698
rect 49608 11348 49660 11354
rect 49608 11290 49660 11296
rect 50080 11150 50108 12582
rect 50160 12164 50212 12170
rect 50160 12106 50212 12112
rect 50172 11898 50200 12106
rect 50294 11996 50602 12016
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11920 50602 11940
rect 50160 11892 50212 11898
rect 50160 11834 50212 11840
rect 50068 11144 50120 11150
rect 50068 11086 50120 11092
rect 48596 11076 48648 11082
rect 48596 11018 48648 11024
rect 48412 10668 48464 10674
rect 48412 10610 48464 10616
rect 48608 10266 48636 11018
rect 50294 10908 50602 10928
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10832 50602 10852
rect 50632 10810 50660 12786
rect 51184 12646 51212 13126
rect 52012 12850 52040 13330
rect 53392 13326 53420 14214
rect 53380 13320 53432 13326
rect 53380 13262 53432 13268
rect 52000 12844 52052 12850
rect 52000 12786 52052 12792
rect 52368 12844 52420 12850
rect 52368 12786 52420 12792
rect 51172 12640 51224 12646
rect 51172 12582 51224 12588
rect 51184 12238 51212 12582
rect 52380 12306 52408 12786
rect 52368 12300 52420 12306
rect 52368 12242 52420 12248
rect 51172 12232 51224 12238
rect 51172 12174 51224 12180
rect 51184 11830 51212 12174
rect 51172 11824 51224 11830
rect 51172 11766 51224 11772
rect 51184 11642 51212 11766
rect 52092 11756 52144 11762
rect 52092 11698 52144 11704
rect 51092 11614 51212 11642
rect 51092 10810 51120 11614
rect 51172 11552 51224 11558
rect 51172 11494 51224 11500
rect 50620 10804 50672 10810
rect 50620 10746 50672 10752
rect 51080 10804 51132 10810
rect 51080 10746 51132 10752
rect 50160 10668 50212 10674
rect 50160 10610 50212 10616
rect 48964 10600 49016 10606
rect 48964 10542 49016 10548
rect 48596 10260 48648 10266
rect 48596 10202 48648 10208
rect 48136 10056 48188 10062
rect 48136 9998 48188 10004
rect 48148 6914 48176 9998
rect 48976 9586 49004 10542
rect 50172 9722 50200 10610
rect 50294 9820 50602 9840
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9744 50602 9764
rect 50160 9716 50212 9722
rect 50160 9658 50212 9664
rect 51184 9654 51212 11494
rect 51540 10056 51592 10062
rect 51540 9998 51592 10004
rect 51172 9648 51224 9654
rect 51172 9590 51224 9596
rect 48964 9580 49016 9586
rect 48964 9522 49016 9528
rect 51552 9382 51580 9998
rect 52104 9450 52132 11698
rect 52380 11370 52408 12242
rect 53668 12238 53696 14758
rect 53760 12918 53788 15302
rect 54852 15020 54904 15026
rect 54852 14962 54904 14968
rect 54864 12986 54892 14962
rect 54944 14952 54996 14958
rect 54944 14894 54996 14900
rect 54956 14006 54984 14894
rect 56428 14414 56456 15438
rect 57336 15428 57388 15434
rect 57336 15370 57388 15376
rect 57348 15162 57376 15370
rect 57336 15156 57388 15162
rect 57336 15098 57388 15104
rect 57336 15020 57388 15026
rect 57336 14962 57388 14968
rect 55956 14408 56008 14414
rect 55956 14350 56008 14356
rect 56416 14408 56468 14414
rect 56416 14350 56468 14356
rect 55588 14340 55640 14346
rect 55588 14282 55640 14288
rect 54944 14000 54996 14006
rect 54944 13942 54996 13948
rect 54852 12980 54904 12986
rect 54852 12922 54904 12928
rect 53748 12912 53800 12918
rect 53748 12854 53800 12860
rect 55496 12844 55548 12850
rect 55496 12786 55548 12792
rect 55404 12776 55456 12782
rect 55404 12718 55456 12724
rect 55416 12238 55444 12718
rect 53656 12232 53708 12238
rect 53656 12174 53708 12180
rect 55404 12232 55456 12238
rect 55404 12174 55456 12180
rect 52920 12164 52972 12170
rect 52920 12106 52972 12112
rect 52380 11354 52500 11370
rect 52932 11354 52960 12106
rect 53656 12096 53708 12102
rect 53656 12038 53708 12044
rect 54392 12096 54444 12102
rect 54392 12038 54444 12044
rect 53288 11688 53340 11694
rect 53288 11630 53340 11636
rect 52380 11348 52512 11354
rect 52380 11342 52460 11348
rect 52460 11290 52512 11296
rect 52920 11348 52972 11354
rect 52920 11290 52972 11296
rect 53300 11150 53328 11630
rect 53288 11144 53340 11150
rect 53288 11086 53340 11092
rect 53300 10674 53328 11086
rect 52920 10668 52972 10674
rect 52920 10610 52972 10616
rect 53288 10668 53340 10674
rect 53288 10610 53340 10616
rect 52184 10464 52236 10470
rect 52184 10406 52236 10412
rect 52092 9444 52144 9450
rect 52092 9386 52144 9392
rect 51172 9376 51224 9382
rect 51172 9318 51224 9324
rect 51540 9376 51592 9382
rect 51540 9318 51592 9324
rect 51184 9042 51212 9318
rect 51172 9036 51224 9042
rect 51172 8978 51224 8984
rect 52196 8974 52224 10406
rect 52932 10266 52960 10610
rect 52920 10260 52972 10266
rect 52920 10202 52972 10208
rect 53300 10130 53328 10610
rect 53288 10124 53340 10130
rect 53288 10066 53340 10072
rect 53668 9654 53696 12038
rect 54404 11150 54432 12038
rect 55416 11762 55444 12174
rect 55404 11756 55456 11762
rect 55404 11698 55456 11704
rect 54392 11144 54444 11150
rect 54392 11086 54444 11092
rect 53748 11076 53800 11082
rect 53748 11018 53800 11024
rect 53760 10266 53788 11018
rect 54760 11008 54812 11014
rect 54760 10950 54812 10956
rect 53748 10260 53800 10266
rect 53748 10202 53800 10208
rect 54772 10062 54800 10950
rect 55508 10810 55536 12786
rect 55600 11898 55628 14282
rect 55968 13870 55996 14350
rect 57348 14074 57376 14962
rect 56692 14068 56744 14074
rect 56692 14010 56744 14016
rect 57336 14068 57388 14074
rect 57336 14010 57388 14016
rect 55956 13864 56008 13870
rect 55956 13806 56008 13812
rect 55968 12782 55996 13806
rect 56704 13326 56732 14010
rect 56692 13320 56744 13326
rect 56692 13262 56744 13268
rect 57244 13184 57296 13190
rect 57244 13126 57296 13132
rect 55956 12776 56008 12782
rect 55956 12718 56008 12724
rect 56600 12640 56652 12646
rect 56600 12582 56652 12588
rect 56612 12238 56640 12582
rect 57256 12306 57284 13126
rect 56876 12300 56928 12306
rect 56876 12242 56928 12248
rect 57244 12300 57296 12306
rect 57244 12242 57296 12248
rect 56600 12232 56652 12238
rect 56600 12174 56652 12180
rect 56784 12096 56836 12102
rect 56784 12038 56836 12044
rect 55588 11892 55640 11898
rect 55588 11834 55640 11840
rect 56796 11830 56824 12038
rect 56784 11824 56836 11830
rect 56784 11766 56836 11772
rect 55956 11552 56008 11558
rect 55956 11494 56008 11500
rect 55496 10804 55548 10810
rect 55496 10746 55548 10752
rect 55968 10742 55996 11494
rect 56888 11218 56916 12242
rect 57532 12238 57560 59162
rect 58624 58880 58676 58886
rect 58624 58822 58676 58828
rect 58636 58614 58664 58822
rect 58624 58608 58676 58614
rect 58624 58550 58676 58556
rect 58440 57860 58492 57866
rect 58440 57802 58492 57808
rect 58452 57050 58480 57802
rect 58440 57044 58492 57050
rect 58440 56986 58492 56992
rect 57704 53508 57756 53514
rect 57704 53450 57756 53456
rect 57716 52698 57744 53450
rect 58164 53440 58216 53446
rect 58164 53382 58216 53388
rect 58176 53174 58204 53382
rect 58164 53168 58216 53174
rect 58164 53110 58216 53116
rect 57704 52692 57756 52698
rect 57704 52634 57756 52640
rect 58532 51400 58584 51406
rect 58532 51342 58584 51348
rect 58544 49434 58572 51342
rect 58532 49428 58584 49434
rect 58532 49370 58584 49376
rect 58532 44736 58584 44742
rect 58532 44678 58584 44684
rect 58544 43790 58572 44678
rect 58532 43784 58584 43790
rect 58532 43726 58584 43732
rect 57888 43648 57940 43654
rect 57888 43590 57940 43596
rect 57900 42702 57928 43590
rect 58164 43308 58216 43314
rect 58164 43250 58216 43256
rect 58176 42906 58204 43250
rect 58164 42900 58216 42906
rect 58164 42842 58216 42848
rect 57888 42696 57940 42702
rect 57888 42638 57940 42644
rect 58440 33924 58492 33930
rect 58440 33866 58492 33872
rect 58452 33114 58480 33866
rect 58532 33856 58584 33862
rect 58532 33798 58584 33804
rect 58440 33108 58492 33114
rect 58440 33050 58492 33056
rect 58544 32502 58572 33798
rect 58532 32496 58584 32502
rect 58532 32438 58584 32444
rect 57888 32428 57940 32434
rect 57888 32370 57940 32376
rect 57900 32026 57928 32370
rect 57888 32020 57940 32026
rect 57888 31962 57940 31968
rect 58532 31816 58584 31822
rect 58532 31758 58584 31764
rect 58544 30938 58572 31758
rect 58532 30932 58584 30938
rect 58532 30874 58584 30880
rect 57888 27328 57940 27334
rect 57888 27270 57940 27276
rect 57900 27062 57928 27270
rect 57888 27056 57940 27062
rect 57888 26998 57940 27004
rect 58164 25900 58216 25906
rect 58164 25842 58216 25848
rect 58176 25498 58204 25842
rect 58164 25492 58216 25498
rect 58164 25434 58216 25440
rect 58532 24064 58584 24070
rect 58532 24006 58584 24012
rect 58544 23798 58572 24006
rect 58532 23792 58584 23798
rect 58532 23734 58584 23740
rect 58440 23044 58492 23050
rect 58440 22986 58492 22992
rect 58452 21146 58480 22986
rect 58532 22976 58584 22982
rect 58532 22918 58584 22924
rect 58544 22710 58572 22918
rect 58532 22704 58584 22710
rect 58532 22646 58584 22652
rect 58440 21140 58492 21146
rect 58440 21082 58492 21088
rect 58440 20868 58492 20874
rect 58440 20810 58492 20816
rect 58452 20058 58480 20810
rect 58440 20052 58492 20058
rect 58440 19994 58492 20000
rect 58072 18624 58124 18630
rect 58072 18566 58124 18572
rect 58084 18358 58112 18566
rect 58072 18352 58124 18358
rect 58072 18294 58124 18300
rect 58164 17536 58216 17542
rect 58164 17478 58216 17484
rect 58176 17270 58204 17478
rect 58164 17264 58216 17270
rect 58164 17206 58216 17212
rect 57796 16516 57848 16522
rect 57796 16458 57848 16464
rect 57808 15706 57836 16458
rect 57888 16448 57940 16454
rect 57888 16390 57940 16396
rect 57900 16182 57928 16390
rect 57888 16176 57940 16182
rect 57888 16118 57940 16124
rect 57796 15700 57848 15706
rect 57796 15642 57848 15648
rect 58072 14272 58124 14278
rect 58072 14214 58124 14220
rect 58084 14006 58112 14214
rect 58072 14000 58124 14006
rect 58072 13942 58124 13948
rect 57520 12232 57572 12238
rect 57520 12174 57572 12180
rect 58440 12096 58492 12102
rect 58440 12038 58492 12044
rect 58452 11830 58480 12038
rect 58440 11824 58492 11830
rect 58440 11766 58492 11772
rect 58622 11792 58678 11801
rect 57244 11756 57296 11762
rect 58622 11727 58624 11736
rect 57244 11698 57296 11704
rect 58676 11727 58678 11736
rect 58624 11698 58676 11704
rect 56876 11212 56928 11218
rect 56876 11154 56928 11160
rect 55956 10736 56008 10742
rect 55956 10678 56008 10684
rect 56888 10470 56916 11154
rect 57256 10810 57284 11698
rect 57336 11076 57388 11082
rect 57336 11018 57388 11024
rect 57244 10804 57296 10810
rect 57244 10746 57296 10752
rect 56876 10464 56928 10470
rect 56876 10406 56928 10412
rect 56888 10130 56916 10406
rect 56876 10124 56928 10130
rect 56876 10066 56928 10072
rect 54760 10056 54812 10062
rect 54760 9998 54812 10004
rect 53748 9988 53800 9994
rect 53748 9930 53800 9936
rect 53656 9648 53708 9654
rect 53656 9590 53708 9596
rect 52552 9580 52604 9586
rect 52552 9522 52604 9528
rect 52564 9178 52592 9522
rect 53012 9512 53064 9518
rect 53012 9454 53064 9460
rect 52552 9172 52604 9178
rect 52552 9114 52604 9120
rect 53024 8974 53052 9454
rect 53760 9382 53788 9930
rect 55312 9512 55364 9518
rect 55312 9454 55364 9460
rect 53748 9376 53800 9382
rect 53748 9318 53800 9324
rect 55324 8974 55352 9454
rect 57348 9450 57376 11018
rect 58256 11008 58308 11014
rect 58256 10950 58308 10956
rect 58268 10742 58296 10950
rect 58256 10736 58308 10742
rect 58256 10678 58308 10684
rect 58256 9920 58308 9926
rect 58256 9862 58308 9868
rect 58268 9654 58296 9862
rect 58256 9648 58308 9654
rect 58256 9590 58308 9596
rect 57336 9444 57388 9450
rect 57336 9386 57388 9392
rect 52184 8968 52236 8974
rect 52184 8910 52236 8916
rect 53012 8968 53064 8974
rect 53012 8910 53064 8916
rect 55312 8968 55364 8974
rect 55312 8910 55364 8916
rect 52644 8900 52696 8906
rect 52644 8842 52696 8848
rect 54116 8900 54168 8906
rect 54116 8842 54168 8848
rect 50294 8732 50602 8752
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8656 50602 8676
rect 48228 8492 48280 8498
rect 48228 8434 48280 8440
rect 50160 8492 50212 8498
rect 50160 8434 50212 8440
rect 48240 8090 48268 8434
rect 48228 8084 48280 8090
rect 48228 8026 48280 8032
rect 50172 7954 50200 8434
rect 50804 8288 50856 8294
rect 50804 8230 50856 8236
rect 50160 7948 50212 7954
rect 50160 7890 50212 7896
rect 50172 7342 50200 7890
rect 50620 7812 50672 7818
rect 50620 7754 50672 7760
rect 50294 7644 50602 7664
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7568 50602 7588
rect 50632 7546 50660 7754
rect 50620 7540 50672 7546
rect 50620 7482 50672 7488
rect 50816 7478 50844 8230
rect 52656 7954 52684 8842
rect 54128 8634 54156 8842
rect 54392 8832 54444 8838
rect 54392 8774 54444 8780
rect 54116 8628 54168 8634
rect 54116 8570 54168 8576
rect 53840 8560 53892 8566
rect 53840 8502 53892 8508
rect 52736 8492 52788 8498
rect 52736 8434 52788 8440
rect 52644 7948 52696 7954
rect 52644 7890 52696 7896
rect 51172 7744 51224 7750
rect 51172 7686 51224 7692
rect 50804 7472 50856 7478
rect 50804 7414 50856 7420
rect 50160 7336 50212 7342
rect 50160 7278 50212 7284
rect 48056 6886 48176 6914
rect 47860 6792 47912 6798
rect 47860 6734 47912 6740
rect 48056 5778 48084 6886
rect 50172 6798 50200 7278
rect 51184 6798 51212 7686
rect 52656 7478 52684 7890
rect 52644 7472 52696 7478
rect 52644 7414 52696 7420
rect 51540 7404 51592 7410
rect 51540 7346 51592 7352
rect 51552 7002 51580 7346
rect 52184 7200 52236 7206
rect 52184 7142 52236 7148
rect 51540 6996 51592 7002
rect 51540 6938 51592 6944
rect 49792 6792 49844 6798
rect 49792 6734 49844 6740
rect 50160 6792 50212 6798
rect 50160 6734 50212 6740
rect 51172 6792 51224 6798
rect 51172 6734 51224 6740
rect 49332 6724 49384 6730
rect 49332 6666 49384 6672
rect 48964 6656 49016 6662
rect 48964 6598 49016 6604
rect 48976 6390 49004 6598
rect 49344 6458 49372 6666
rect 49332 6452 49384 6458
rect 49332 6394 49384 6400
rect 48964 6384 49016 6390
rect 48964 6326 49016 6332
rect 49804 6322 49832 6734
rect 50294 6556 50602 6576
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6480 50602 6500
rect 52196 6390 52224 7142
rect 52184 6384 52236 6390
rect 52184 6326 52236 6332
rect 49792 6316 49844 6322
rect 49792 6258 49844 6264
rect 51172 6112 51224 6118
rect 51172 6054 51224 6060
rect 48044 5772 48096 5778
rect 48044 5714 48096 5720
rect 48056 5642 48084 5714
rect 49608 5704 49660 5710
rect 49608 5646 49660 5652
rect 48044 5636 48096 5642
rect 48044 5578 48096 5584
rect 48228 5568 48280 5574
rect 48228 5510 48280 5516
rect 47676 4616 47728 4622
rect 47676 4558 47728 4564
rect 48240 4554 48268 5510
rect 48228 4548 48280 4554
rect 48228 4490 48280 4496
rect 46952 4078 46980 4134
rect 47032 4140 47084 4146
rect 47032 4082 47084 4088
rect 46940 4072 46992 4078
rect 46940 4014 46992 4020
rect 45284 4004 45336 4010
rect 45284 3946 45336 3952
rect 43812 3732 43864 3738
rect 43812 3674 43864 3680
rect 48240 3534 48268 4490
rect 48964 3936 49016 3942
rect 48964 3878 49016 3884
rect 48976 3534 49004 3878
rect 49620 3738 49648 5646
rect 50294 5468 50602 5488
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5392 50602 5412
rect 51184 5302 51212 6054
rect 51172 5296 51224 5302
rect 51172 5238 51224 5244
rect 52656 5234 52684 7414
rect 52748 7410 52776 8434
rect 52736 7404 52788 7410
rect 52736 7346 52788 7352
rect 52748 6866 52776 7346
rect 52736 6860 52788 6866
rect 52736 6802 52788 6808
rect 52748 6254 52776 6802
rect 52736 6248 52788 6254
rect 52736 6190 52788 6196
rect 52748 5914 52776 6190
rect 52736 5908 52788 5914
rect 52736 5850 52788 5856
rect 52644 5228 52696 5234
rect 52644 5170 52696 5176
rect 50160 5160 50212 5166
rect 50160 5102 50212 5108
rect 50172 4622 50200 5102
rect 50436 5024 50488 5030
rect 50436 4966 50488 4972
rect 50448 4622 50476 4966
rect 52748 4622 52776 5850
rect 53852 5710 53880 8502
rect 54116 8492 54168 8498
rect 54116 8434 54168 8440
rect 54128 8090 54156 8434
rect 54116 8084 54168 8090
rect 54116 8026 54168 8032
rect 54024 7812 54076 7818
rect 54024 7754 54076 7760
rect 54036 7546 54064 7754
rect 54024 7540 54076 7546
rect 54024 7482 54076 7488
rect 54404 7478 54432 8774
rect 55324 8294 55352 8910
rect 56600 8900 56652 8906
rect 56600 8842 56652 8848
rect 58440 8900 58492 8906
rect 58440 8842 58492 8848
rect 55864 8832 55916 8838
rect 55864 8774 55916 8780
rect 55312 8288 55364 8294
rect 55312 8230 55364 8236
rect 55324 7886 55352 8230
rect 55312 7880 55364 7886
rect 55312 7822 55364 7828
rect 54392 7472 54444 7478
rect 54392 7414 54444 7420
rect 55324 7410 55352 7822
rect 54208 7404 54260 7410
rect 54208 7346 54260 7352
rect 55312 7404 55364 7410
rect 55312 7346 55364 7352
rect 54220 7002 54248 7346
rect 54208 6996 54260 7002
rect 54208 6938 54260 6944
rect 55324 6798 55352 7346
rect 55876 6798 55904 8774
rect 56612 8090 56640 8842
rect 58452 8090 58480 8842
rect 58532 8832 58584 8838
rect 58532 8774 58584 8780
rect 56600 8084 56652 8090
rect 56600 8026 56652 8032
rect 58440 8084 58492 8090
rect 58440 8026 58492 8032
rect 55956 7812 56008 7818
rect 55956 7754 56008 7760
rect 56784 7812 56836 7818
rect 56784 7754 56836 7760
rect 55968 7546 55996 7754
rect 55956 7540 56008 7546
rect 55956 7482 56008 7488
rect 56796 7002 56824 7754
rect 56784 6996 56836 7002
rect 56784 6938 56836 6944
rect 58544 6798 58572 8774
rect 55312 6792 55364 6798
rect 55312 6734 55364 6740
rect 55864 6792 55916 6798
rect 55864 6734 55916 6740
rect 58532 6792 58584 6798
rect 58532 6734 58584 6740
rect 54668 6724 54720 6730
rect 54668 6666 54720 6672
rect 54680 6458 54708 6666
rect 54668 6452 54720 6458
rect 54668 6394 54720 6400
rect 54116 6316 54168 6322
rect 54116 6258 54168 6264
rect 53840 5704 53892 5710
rect 53840 5646 53892 5652
rect 54128 5370 54156 6258
rect 54116 5364 54168 5370
rect 54116 5306 54168 5312
rect 54024 5228 54076 5234
rect 54024 5170 54076 5176
rect 50160 4616 50212 4622
rect 50160 4558 50212 4564
rect 50436 4616 50488 4622
rect 50436 4558 50488 4564
rect 52736 4616 52788 4622
rect 52736 4558 52788 4564
rect 50172 4162 50200 4558
rect 51540 4480 51592 4486
rect 51540 4422 51592 4428
rect 50294 4380 50602 4400
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4304 50602 4324
rect 49988 4146 50200 4162
rect 51552 4146 51580 4422
rect 52748 4146 52776 4558
rect 53564 4548 53616 4554
rect 53564 4490 53616 4496
rect 53380 4480 53432 4486
rect 53380 4422 53432 4428
rect 53392 4214 53420 4422
rect 53380 4208 53432 4214
rect 53380 4150 53432 4156
rect 49976 4140 50200 4146
rect 50028 4134 50200 4140
rect 49976 4082 50028 4088
rect 49608 3732 49660 3738
rect 49608 3674 49660 3680
rect 50172 3534 50200 4134
rect 51540 4140 51592 4146
rect 51540 4082 51592 4088
rect 52736 4140 52788 4146
rect 52736 4082 52788 4088
rect 50620 3936 50672 3942
rect 50620 3878 50672 3884
rect 50632 3534 50660 3878
rect 52748 3534 52776 4082
rect 53576 3738 53604 4490
rect 53564 3732 53616 3738
rect 53564 3674 53616 3680
rect 48228 3528 48280 3534
rect 48228 3470 48280 3476
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50620 3528 50672 3534
rect 50620 3470 50672 3476
rect 52736 3528 52788 3534
rect 52736 3470 52788 3476
rect 43536 3188 43588 3194
rect 43536 3130 43588 3136
rect 42708 3120 42760 3126
rect 42708 3062 42760 3068
rect 48240 3058 48268 3470
rect 52276 3460 52328 3466
rect 52276 3402 52328 3408
rect 51724 3392 51776 3398
rect 51724 3334 51776 3340
rect 50294 3292 50602 3312
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3216 50602 3236
rect 51736 3126 51764 3334
rect 52288 3194 52316 3402
rect 52276 3188 52328 3194
rect 52276 3130 52328 3136
rect 51724 3120 51776 3126
rect 51724 3062 51776 3068
rect 52748 3058 52776 3470
rect 39856 3052 39908 3058
rect 39856 2994 39908 3000
rect 42432 3052 42484 3058
rect 42432 2994 42484 3000
rect 48228 3052 48280 3058
rect 48228 2994 48280 3000
rect 52736 3052 52788 3058
rect 52736 2994 52788 3000
rect 54036 2922 54064 5170
rect 54116 3936 54168 3942
rect 54116 3878 54168 3884
rect 54128 3126 54156 3878
rect 54116 3120 54168 3126
rect 54116 3062 54168 3068
rect 38844 2916 38896 2922
rect 38844 2858 38896 2864
rect 54024 2916 54076 2922
rect 54024 2858 54076 2864
rect 38752 2644 38804 2650
rect 38752 2586 38804 2592
rect 34244 2440 34296 2446
rect 34244 2382 34296 2388
rect 36452 2440 36504 2446
rect 36452 2382 36504 2388
rect 38568 2440 38620 2446
rect 38568 2382 38620 2388
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 28540 2372 28592 2378
rect 28540 2314 28592 2320
rect 32 800 60 2314
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 34256 800 34284 2382
rect 50294 2204 50602 2224
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2128 50602 2148
rect 18 0 74 800
rect 34242 0 34298 800
<< via2 >>
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 34940 60410 34996 60412
rect 35020 60410 35076 60412
rect 35100 60410 35156 60412
rect 35180 60410 35236 60412
rect 34940 60358 34986 60410
rect 34986 60358 34996 60410
rect 35020 60358 35050 60410
rect 35050 60358 35062 60410
rect 35062 60358 35076 60410
rect 35100 60358 35114 60410
rect 35114 60358 35126 60410
rect 35126 60358 35156 60410
rect 35180 60358 35190 60410
rect 35190 60358 35236 60410
rect 34940 60356 34996 60358
rect 35020 60356 35076 60358
rect 35100 60356 35156 60358
rect 35180 60356 35236 60358
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 3698 50632 3754 50688
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 19580 59866 19636 59868
rect 19660 59866 19716 59868
rect 19740 59866 19796 59868
rect 19820 59866 19876 59868
rect 19580 59814 19626 59866
rect 19626 59814 19636 59866
rect 19660 59814 19690 59866
rect 19690 59814 19702 59866
rect 19702 59814 19716 59866
rect 19740 59814 19754 59866
rect 19754 59814 19766 59866
rect 19766 59814 19796 59866
rect 19820 59814 19830 59866
rect 19830 59814 19876 59866
rect 19580 59812 19636 59814
rect 19660 59812 19716 59814
rect 19740 59812 19796 59814
rect 19820 59812 19876 59814
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 19580 58778 19636 58780
rect 19660 58778 19716 58780
rect 19740 58778 19796 58780
rect 19820 58778 19876 58780
rect 19580 58726 19626 58778
rect 19626 58726 19636 58778
rect 19660 58726 19690 58778
rect 19690 58726 19702 58778
rect 19702 58726 19716 58778
rect 19740 58726 19754 58778
rect 19754 58726 19766 58778
rect 19766 58726 19796 58778
rect 19820 58726 19830 58778
rect 19830 58726 19876 58778
rect 19580 58724 19636 58726
rect 19660 58724 19716 58726
rect 19740 58724 19796 58726
rect 19820 58724 19876 58726
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 34940 59322 34996 59324
rect 35020 59322 35076 59324
rect 35100 59322 35156 59324
rect 35180 59322 35236 59324
rect 34940 59270 34986 59322
rect 34986 59270 34996 59322
rect 35020 59270 35050 59322
rect 35050 59270 35062 59322
rect 35062 59270 35076 59322
rect 35100 59270 35114 59322
rect 35114 59270 35126 59322
rect 35126 59270 35156 59322
rect 35180 59270 35190 59322
rect 35190 59270 35236 59322
rect 34940 59268 34996 59270
rect 35020 59268 35076 59270
rect 35100 59268 35156 59270
rect 35180 59268 35236 59270
rect 34940 58234 34996 58236
rect 35020 58234 35076 58236
rect 35100 58234 35156 58236
rect 35180 58234 35236 58236
rect 34940 58182 34986 58234
rect 34986 58182 34996 58234
rect 35020 58182 35050 58234
rect 35050 58182 35062 58234
rect 35062 58182 35076 58234
rect 35100 58182 35114 58234
rect 35114 58182 35126 58234
rect 35126 58182 35156 58234
rect 35180 58182 35190 58234
rect 35190 58182 35236 58234
rect 34940 58180 34996 58182
rect 35020 58180 35076 58182
rect 35100 58180 35156 58182
rect 35180 58180 35236 58182
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 50300 59866 50356 59868
rect 50380 59866 50436 59868
rect 50460 59866 50516 59868
rect 50540 59866 50596 59868
rect 50300 59814 50346 59866
rect 50346 59814 50356 59866
rect 50380 59814 50410 59866
rect 50410 59814 50422 59866
rect 50422 59814 50436 59866
rect 50460 59814 50474 59866
rect 50474 59814 50486 59866
rect 50486 59814 50516 59866
rect 50540 59814 50550 59866
rect 50550 59814 50596 59866
rect 50300 59812 50356 59814
rect 50380 59812 50436 59814
rect 50460 59812 50516 59814
rect 50540 59812 50596 59814
rect 50300 58778 50356 58780
rect 50380 58778 50436 58780
rect 50460 58778 50516 58780
rect 50540 58778 50596 58780
rect 50300 58726 50346 58778
rect 50346 58726 50356 58778
rect 50380 58726 50410 58778
rect 50410 58726 50422 58778
rect 50422 58726 50436 58778
rect 50460 58726 50474 58778
rect 50474 58726 50486 58778
rect 50486 58726 50516 58778
rect 50540 58726 50550 58778
rect 50550 58726 50596 58778
rect 50300 58724 50356 58726
rect 50380 58724 50436 58726
rect 50460 58724 50516 58726
rect 50540 58724 50596 58726
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 58622 11756 58678 11792
rect 58622 11736 58624 11756
rect 58624 11736 58676 11756
rect 58676 11736 58678 11756
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
<< metal3 >>
rect 4208 60416 4528 60417
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 60351 4528 60352
rect 34928 60416 35248 60417
rect 34928 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35248 60416
rect 34928 60351 35248 60352
rect 19568 59872 19888 59873
rect 19568 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19888 59872
rect 19568 59807 19888 59808
rect 50288 59872 50608 59873
rect 50288 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50608 59872
rect 50288 59807 50608 59808
rect 4208 59328 4528 59329
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 59263 4528 59264
rect 34928 59328 35248 59329
rect 34928 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35248 59328
rect 34928 59263 35248 59264
rect 19568 58784 19888 58785
rect 19568 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19888 58784
rect 19568 58719 19888 58720
rect 50288 58784 50608 58785
rect 50288 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50608 58784
rect 50288 58719 50608 58720
rect 4208 58240 4528 58241
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 58175 4528 58176
rect 34928 58240 35248 58241
rect 34928 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35248 58240
rect 34928 58175 35248 58176
rect 19568 57696 19888 57697
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 57631 19888 57632
rect 50288 57696 50608 57697
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 57631 50608 57632
rect 4208 57152 4528 57153
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 57087 4528 57088
rect 34928 57152 35248 57153
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 57087 35248 57088
rect 19568 56608 19888 56609
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 56543 19888 56544
rect 50288 56608 50608 56609
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 56543 50608 56544
rect 4208 56064 4528 56065
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 55999 4528 56000
rect 34928 56064 35248 56065
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 55999 35248 56000
rect 19568 55520 19888 55521
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 55455 19888 55456
rect 50288 55520 50608 55521
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 55455 50608 55456
rect 4208 54976 4528 54977
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 54911 4528 54912
rect 34928 54976 35248 54977
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 54911 35248 54912
rect 19568 54432 19888 54433
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 54367 19888 54368
rect 50288 54432 50608 54433
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 54367 50608 54368
rect 4208 53888 4528 53889
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 53823 4528 53824
rect 34928 53888 35248 53889
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 53823 35248 53824
rect 19568 53344 19888 53345
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 53279 19888 53280
rect 50288 53344 50608 53345
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 53279 50608 53280
rect 4208 52800 4528 52801
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 52735 4528 52736
rect 34928 52800 35248 52801
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 52735 35248 52736
rect 19568 52256 19888 52257
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 52191 19888 52192
rect 50288 52256 50608 52257
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 52191 50608 52192
rect 4208 51712 4528 51713
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 51647 4528 51648
rect 34928 51712 35248 51713
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 51647 35248 51648
rect 19568 51168 19888 51169
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 51103 19888 51104
rect 50288 51168 50608 51169
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 51103 50608 51104
rect 0 50690 800 50720
rect 3693 50690 3759 50693
rect 0 50688 3759 50690
rect 0 50632 3698 50688
rect 3754 50632 3759 50688
rect 0 50630 3759 50632
rect 0 50600 800 50630
rect 3693 50627 3759 50630
rect 4208 50624 4528 50625
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 50559 4528 50560
rect 34928 50624 35248 50625
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 50559 35248 50560
rect 19568 50080 19888 50081
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 50015 19888 50016
rect 50288 50080 50608 50081
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 50015 50608 50016
rect 4208 49536 4528 49537
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 49471 4528 49472
rect 34928 49536 35248 49537
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 49471 35248 49472
rect 19568 48992 19888 48993
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 48927 19888 48928
rect 50288 48992 50608 48993
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 48927 50608 48928
rect 4208 48448 4528 48449
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 48383 4528 48384
rect 34928 48448 35248 48449
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 48383 35248 48384
rect 19568 47904 19888 47905
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 47839 19888 47840
rect 50288 47904 50608 47905
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 47839 50608 47840
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 50288 46816 50608 46817
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 46751 50608 46752
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 50288 45728 50608 45729
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 45663 50608 45664
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 50288 44640 50608 44641
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 44575 50608 44576
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 50288 43552 50608 43553
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 43487 50608 43488
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 50288 42464 50608 42465
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 42399 50608 42400
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 50288 41376 50608 41377
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 41311 50608 41312
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 50288 40288 50608 40289
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 40223 50608 40224
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 50288 39200 50608 39201
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 39135 50608 39136
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 50288 38112 50608 38113
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 38047 50608 38048
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 50288 37024 50608 37025
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 36959 50608 36960
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 50288 35936 50608 35937
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 35871 50608 35872
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 50288 34848 50608 34849
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 34783 50608 34784
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 50288 33760 50608 33761
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 33695 50608 33696
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 50288 32672 50608 32673
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 32607 50608 32608
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 50288 31584 50608 31585
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 31519 50608 31520
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 50288 30496 50608 30497
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 30431 50608 30432
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 50288 29408 50608 29409
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 29343 50608 29344
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 50288 28320 50608 28321
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 28255 50608 28256
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 50288 27232 50608 27233
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 27167 50608 27168
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 50288 26144 50608 26145
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 26079 50608 26080
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 50288 25056 50608 25057
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 24991 50608 24992
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 50288 23968 50608 23969
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 23903 50608 23904
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 50288 22880 50608 22881
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 22815 50608 22816
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 50288 21792 50608 21793
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 21727 50608 21728
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 50288 20704 50608 20705
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 20639 50608 20640
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 50288 19616 50608 19617
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 19551 50608 19552
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 50288 18528 50608 18529
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 18463 50608 18464
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 50288 17440 50608 17441
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 17375 50608 17376
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 50288 16352 50608 16353
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 16287 50608 16288
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 50288 15264 50608 15265
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 15199 50608 15200
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 50288 14176 50608 14177
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 14111 50608 14112
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 50288 13088 50608 13089
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 13023 50608 13024
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 50288 12000 50608 12001
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 11935 50608 11936
rect 58617 11794 58683 11797
rect 59716 11794 60516 11824
rect 58617 11792 60516 11794
rect 58617 11736 58622 11792
rect 58678 11736 60516 11792
rect 58617 11734 60516 11736
rect 58617 11731 58683 11734
rect 59716 11704 60516 11734
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 50288 10912 50608 10913
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 10847 50608 10848
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 50288 9824 50608 9825
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 9759 50608 9760
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 50288 8736 50608 8737
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 8671 50608 8672
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 50288 7648 50608 7649
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 7583 50608 7584
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 50288 6560 50608 6561
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 6495 50608 6496
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 50288 5472 50608 5473
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 5407 50608 5408
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 50288 4384 50608 4385
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 4319 50608 4320
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 50288 3296 50608 3297
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 3231 50608 3232
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 50288 2208 50608 2209
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2143 50608 2144
<< via3 >>
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 34936 60412 35000 60416
rect 34936 60356 34940 60412
rect 34940 60356 34996 60412
rect 34996 60356 35000 60412
rect 34936 60352 35000 60356
rect 35016 60412 35080 60416
rect 35016 60356 35020 60412
rect 35020 60356 35076 60412
rect 35076 60356 35080 60412
rect 35016 60352 35080 60356
rect 35096 60412 35160 60416
rect 35096 60356 35100 60412
rect 35100 60356 35156 60412
rect 35156 60356 35160 60412
rect 35096 60352 35160 60356
rect 35176 60412 35240 60416
rect 35176 60356 35180 60412
rect 35180 60356 35236 60412
rect 35236 60356 35240 60412
rect 35176 60352 35240 60356
rect 19576 59868 19640 59872
rect 19576 59812 19580 59868
rect 19580 59812 19636 59868
rect 19636 59812 19640 59868
rect 19576 59808 19640 59812
rect 19656 59868 19720 59872
rect 19656 59812 19660 59868
rect 19660 59812 19716 59868
rect 19716 59812 19720 59868
rect 19656 59808 19720 59812
rect 19736 59868 19800 59872
rect 19736 59812 19740 59868
rect 19740 59812 19796 59868
rect 19796 59812 19800 59868
rect 19736 59808 19800 59812
rect 19816 59868 19880 59872
rect 19816 59812 19820 59868
rect 19820 59812 19876 59868
rect 19876 59812 19880 59868
rect 19816 59808 19880 59812
rect 50296 59868 50360 59872
rect 50296 59812 50300 59868
rect 50300 59812 50356 59868
rect 50356 59812 50360 59868
rect 50296 59808 50360 59812
rect 50376 59868 50440 59872
rect 50376 59812 50380 59868
rect 50380 59812 50436 59868
rect 50436 59812 50440 59868
rect 50376 59808 50440 59812
rect 50456 59868 50520 59872
rect 50456 59812 50460 59868
rect 50460 59812 50516 59868
rect 50516 59812 50520 59868
rect 50456 59808 50520 59812
rect 50536 59868 50600 59872
rect 50536 59812 50540 59868
rect 50540 59812 50596 59868
rect 50596 59812 50600 59868
rect 50536 59808 50600 59812
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 34936 59324 35000 59328
rect 34936 59268 34940 59324
rect 34940 59268 34996 59324
rect 34996 59268 35000 59324
rect 34936 59264 35000 59268
rect 35016 59324 35080 59328
rect 35016 59268 35020 59324
rect 35020 59268 35076 59324
rect 35076 59268 35080 59324
rect 35016 59264 35080 59268
rect 35096 59324 35160 59328
rect 35096 59268 35100 59324
rect 35100 59268 35156 59324
rect 35156 59268 35160 59324
rect 35096 59264 35160 59268
rect 35176 59324 35240 59328
rect 35176 59268 35180 59324
rect 35180 59268 35236 59324
rect 35236 59268 35240 59324
rect 35176 59264 35240 59268
rect 19576 58780 19640 58784
rect 19576 58724 19580 58780
rect 19580 58724 19636 58780
rect 19636 58724 19640 58780
rect 19576 58720 19640 58724
rect 19656 58780 19720 58784
rect 19656 58724 19660 58780
rect 19660 58724 19716 58780
rect 19716 58724 19720 58780
rect 19656 58720 19720 58724
rect 19736 58780 19800 58784
rect 19736 58724 19740 58780
rect 19740 58724 19796 58780
rect 19796 58724 19800 58780
rect 19736 58720 19800 58724
rect 19816 58780 19880 58784
rect 19816 58724 19820 58780
rect 19820 58724 19876 58780
rect 19876 58724 19880 58780
rect 19816 58720 19880 58724
rect 50296 58780 50360 58784
rect 50296 58724 50300 58780
rect 50300 58724 50356 58780
rect 50356 58724 50360 58780
rect 50296 58720 50360 58724
rect 50376 58780 50440 58784
rect 50376 58724 50380 58780
rect 50380 58724 50436 58780
rect 50436 58724 50440 58780
rect 50376 58720 50440 58724
rect 50456 58780 50520 58784
rect 50456 58724 50460 58780
rect 50460 58724 50516 58780
rect 50516 58724 50520 58780
rect 50456 58720 50520 58724
rect 50536 58780 50600 58784
rect 50536 58724 50540 58780
rect 50540 58724 50596 58780
rect 50596 58724 50600 58780
rect 50536 58720 50600 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 34936 58236 35000 58240
rect 34936 58180 34940 58236
rect 34940 58180 34996 58236
rect 34996 58180 35000 58236
rect 34936 58176 35000 58180
rect 35016 58236 35080 58240
rect 35016 58180 35020 58236
rect 35020 58180 35076 58236
rect 35076 58180 35080 58236
rect 35016 58176 35080 58180
rect 35096 58236 35160 58240
rect 35096 58180 35100 58236
rect 35100 58180 35156 58236
rect 35156 58180 35160 58236
rect 35096 58176 35160 58180
rect 35176 58236 35240 58240
rect 35176 58180 35180 58236
rect 35180 58180 35236 58236
rect 35236 58180 35240 58236
rect 35176 58176 35240 58180
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 60416 4528 60432
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36212 4528 36416
rect 4208 35976 4250 36212
rect 4486 35976 4528 36212
rect 4208 35392 4528 35976
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5576 4528 5952
rect 4208 5340 4250 5576
rect 4486 5340 4528 5576
rect 4208 4928 4528 5340
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 59872 19888 60432
rect 19568 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19888 59872
rect 19568 58784 19888 59808
rect 19568 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19888 58784
rect 19568 57696 19888 58720
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51530 19888 52192
rect 19568 51294 19610 51530
rect 19846 51294 19888 51530
rect 19568 51168 19888 51294
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20894 19888 21728
rect 19568 20704 19610 20894
rect 19846 20704 19888 20894
rect 19568 20640 19576 20704
rect 19640 20640 19656 20658
rect 19720 20640 19736 20658
rect 19800 20640 19816 20658
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 60416 35248 60432
rect 34928 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35248 60416
rect 34928 59328 35248 60352
rect 34928 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35248 59328
rect 34928 58240 35248 59264
rect 34928 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35248 58240
rect 34928 57152 35248 58176
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36212 35248 36416
rect 34928 35976 34970 36212
rect 35206 35976 35248 36212
rect 34928 35392 35248 35976
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5576 35248 5952
rect 34928 5340 34970 5576
rect 35206 5340 35248 5576
rect 34928 4928 35248 5340
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 59872 50608 60432
rect 50288 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50608 59872
rect 50288 58784 50608 59808
rect 50288 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50608 58784
rect 50288 57696 50608 58720
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51530 50608 52192
rect 50288 51294 50330 51530
rect 50566 51294 50608 51530
rect 50288 51168 50608 51294
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20894 50608 21728
rect 50288 20704 50330 20894
rect 50566 20704 50608 20894
rect 50288 20640 50296 20704
rect 50360 20640 50376 20658
rect 50440 20640 50456 20658
rect 50520 20640 50536 20658
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
<< via4 >>
rect 4250 35976 4486 36212
rect 4250 5340 4486 5576
rect 19610 51294 19846 51530
rect 19610 20704 19846 20894
rect 19610 20658 19640 20704
rect 19640 20658 19656 20704
rect 19656 20658 19720 20704
rect 19720 20658 19736 20704
rect 19736 20658 19800 20704
rect 19800 20658 19816 20704
rect 19816 20658 19846 20704
rect 34970 35976 35206 36212
rect 34970 5340 35206 5576
rect 50330 51294 50566 51530
rect 50330 20704 50566 20894
rect 50330 20658 50360 20704
rect 50360 20658 50376 20704
rect 50376 20658 50440 20704
rect 50440 20658 50456 20704
rect 50456 20658 50520 20704
rect 50520 20658 50536 20704
rect 50536 20658 50566 20704
<< metal5 >>
rect 1104 51530 59340 51572
rect 1104 51294 19610 51530
rect 19846 51294 50330 51530
rect 50566 51294 59340 51530
rect 1104 51252 59340 51294
rect 1104 36212 59340 36254
rect 1104 35976 4250 36212
rect 4486 35976 34970 36212
rect 35206 35976 59340 36212
rect 1104 35934 59340 35976
rect 1104 20894 59340 20936
rect 1104 20658 19610 20894
rect 19846 20658 50330 20894
rect 50566 20658 59340 20894
rect 1104 20616 59340 20658
rect 1104 5576 59340 5618
rect 1104 5340 4250 5576
rect 4486 5340 34970 5576
rect 35206 5340 59340 5576
rect 1104 5298 59340 5340
use sky130_fd_sc_hd__diode_2  ANTENNA_0 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform -1 0 1748 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1632082664
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_11
timestamp 1632082664
transform 1 0 2116 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output2 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform -1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1632082664
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1632082664
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1632082664
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1632082664
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1632082664
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1632082664
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1632082664
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1632082664
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1632082664
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1632082664
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1632082664
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1632082664
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_81
timestamp 1632082664
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1632082664
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1632082664
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1632082664
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1632082664
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_97
timestamp 1632082664
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1632082664
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1632082664
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1632082664
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1383_ sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 11684 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1382_
timestamp 1632082664
transform 1 0 11500 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1632082664
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1632082664
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1632082664
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1632082664
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1386_
timestamp 1632082664
transform 1 0 13340 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1632082664
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1632082664
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1632082664
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_129
timestamp 1632082664
transform 1 0 12972 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1632082664
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_149
timestamp 1632082664
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1632082664
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1632082664
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_169
timestamp 1632082664
transform 1 0 16652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1395_
timestamp 1632082664
transform 1 0 17204 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1393_
timestamp 1632082664
transform 1 0 16652 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1632082664
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1632082664
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1632082664
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_185
timestamp 1632082664
transform 1 0 18124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_197
timestamp 1632082664
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1397_
timestamp 1632082664
transform 1 0 19872 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1396_
timestamp 1632082664
transform 1 0 18492 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_1_205
timestamp 1632082664
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1632082664
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_203
timestamp 1632082664
transform 1 0 19780 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1632082664
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1632082664
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_225
timestamp 1632082664
transform 1 0 21804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1632082664
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1398_
timestamp 1632082664
transform 1 0 21804 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1632082664
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1632082664
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1632082664
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1632082664
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_241
timestamp 1632082664
transform 1 0 23276 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1741_
timestamp 1632082664
transform 1 0 22448 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_1_231
timestamp 1632082664
transform 1 0 22356 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_248
timestamp 1632082664
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1632082664
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_269
timestamp 1632082664
transform 1 0 25852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1739_
timestamp 1632082664
transform 1 0 24380 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1737_
timestamp 1632082664
transform 1 0 24288 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_1_268
timestamp 1632082664
transform 1 0 25760 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1632082664
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1735_
timestamp 1632082664
transform 1 0 26956 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1734_
timestamp 1632082664
transform 1 0 26956 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1632082664
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1632082664
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1632082664
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_297
timestamp 1632082664
transform 1 0 28428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1742_
timestamp 1632082664
transform 1 0 28796 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_0_309
timestamp 1632082664
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1632082664
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_297
timestamp 1632082664
transform 1 0 28428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1632082664
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1632082664
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_317
timestamp 1632082664
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_321
timestamp 1632082664
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1632082664
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_337
timestamp 1632082664
transform 1 0 32108 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_349
timestamp 1632082664
transform 1 0 33212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1767_
timestamp 1632082664
transform 1 0 32660 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1632082664
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1632082664
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1632082664
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1632082664
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1 sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 33948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1811_
timestamp 1632082664
transform 1 0 34684 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1789_
timestamp 1632082664
transform 1 0 34500 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1632082664
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_359
timestamp 1632082664
transform 1 0 34132 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1632082664
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_381
timestamp 1632082664
transform 1 0 36156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1844_
timestamp 1632082664
transform 1 0 37260 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1822_
timestamp 1632082664
transform 1 0 37260 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_1_379
timestamp 1632082664
transform 1 0 35972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1632082664
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1632082664
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1632082664
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1632082664
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_409
timestamp 1632082664
transform 1 0 38732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1866_
timestamp 1632082664
transform 1 0 39100 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_1_409
timestamp 1632082664
transform 1 0 38732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_429
timestamp 1632082664
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_433
timestamp 1632082664
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_421
timestamp 1632082664
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1632082664
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1632082664
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1632082664
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1987_
timestamp 1632082664
transform 1 0 42412 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_0_449
timestamp 1632082664
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1632082664
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1632082664
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1632082664
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1632082664
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_477
timestamp 1632082664
transform 1 0 44988 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_465
timestamp 1632082664
transform 1 0 43884 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_477
timestamp 1632082664
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_461
timestamp 1632082664
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1632082664
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1632082664
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_489
timestamp 1632082664
transform 1 0 46092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_489
timestamp 1632082664
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_517
timestamp 1632082664
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_505
timestamp 1632082664
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_517
timestamp 1632082664
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_505
timestamp 1632082664
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1632082664
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1632082664
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_501
timestamp 1632082664
transform 1 0 47196 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1632082664
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_529
timestamp 1632082664
transform 1 0 49772 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1508_
timestamp 1632082664
transform 1 0 50784 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_0_533
timestamp 1632082664
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1632082664
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_537
timestamp 1632082664
transform 1 0 50508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1632082664
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1512_
timestamp 1632082664
transform 1 0 52716 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_0_561
timestamp 1632082664
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_545
timestamp 1632082664
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1632082664
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1632082664
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_556
timestamp 1632082664
transform 1 0 52256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1632082664
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_577
timestamp 1632082664
transform 1 0 54188 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_573
timestamp 1632082664
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_601
timestamp 1632082664
transform 1 0 56396 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_589
timestamp 1632082664
transform 1 0 55292 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_601
timestamp 1632082664
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_589
timestamp 1632082664
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1632082664
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1632082664
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_617
timestamp 1632082664
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_617
timestamp 1632082664
transform 1 0 57868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1632082664
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1632082664
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_613
timestamp 1632082664
transform 1 0 57500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1632082664
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_629
timestamp 1632082664
transform 1 0 58972 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_629
timestamp 1632082664
transform 1 0 58972 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1632082664
transform -1 0 59340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1632082664
transform -1 0 59340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1632082664
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1632082664
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1632082664
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_29
timestamp 1632082664
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1366_
timestamp 1632082664
transform 1 0 4600 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1632082664
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_37
timestamp 1632082664
transform 1 0 4508 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1632082664
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_54
timestamp 1632082664
transform 1 0 6072 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp 1632082664
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_66
timestamp 1632082664
transform 1 0 7176 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1380_
timestamp 1632082664
transform 1 0 10396 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1632082664
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1632082664
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1632082664
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1632082664
transform 1 0 11868 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_129
timestamp 1632082664
transform 1 0 12972 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1387_
timestamp 1632082664
transform 1 0 14076 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1632082664
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1632082664
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1391_
timestamp 1632082664
transform 1 0 15916 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_157
timestamp 1632082664
transform 1 0 15548 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_177
timestamp 1632082664
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1632082664
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1394_
timestamp 1632082664
transform 1 0 19228 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1632082664
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1632082664
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1399_
timestamp 1632082664
transform 1 0 21068 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_213
timestamp 1632082664
transform 1 0 20700 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1632082664
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1632082664
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1736_
timestamp 1632082664
transform 1 0 24840 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1632082664
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_257
timestamp 1632082664
transform 1 0 24748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1632082664
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_253
timestamp 1632082664
transform 1 0 24380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1733_
timestamp 1632082664
transform 1 0 26680 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_274
timestamp 1632082664
transform 1 0 26312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1632082664
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1725_
timestamp 1632082664
transform 1 0 29624 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_2_294
timestamp 1632082664
transform 1 0 28152 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1632082664
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_309
timestamp 1632082664
transform 1 0 29532 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_326
timestamp 1632082664
transform 1 0 31096 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1756_
timestamp 1632082664
transform 1 0 32568 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_338
timestamp 1632082664
transform 1 0 32200 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_358
timestamp 1632082664
transform 1 0 34040 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1778_
timestamp 1632082664
transform 1 0 34684 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1632082664
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1800_
timestamp 1632082664
transform 1 0 36524 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_381
timestamp 1632082664
transform 1 0 36156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1632082664
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_401
timestamp 1632082664
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1888_
timestamp 1632082664
transform 1 0 39836 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_2_437
timestamp 1632082664
transform 1 0 41308 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1632082664
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1632082664
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1965_
timestamp 1632082664
transform 1 0 42412 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_2_465
timestamp 1632082664
transform 1 0 43884 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_477
timestamp 1632082664
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1632082664
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_473
timestamp 1632082664
transform 1 0 44620 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_489
timestamp 1632082664
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_501
timestamp 1632082664
transform 1 0 47196 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1605_
timestamp 1632082664
transform 1 0 48208 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_2_509
timestamp 1632082664
transform 1 0 47932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_533
timestamp 1632082664
transform 1 0 50140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1507_
timestamp 1632082664
transform 1 0 50324 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1632082664
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_528
timestamp 1632082664
transform 1 0 49680 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1509_
timestamp 1632082664
transform 1 0 52164 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_551
timestamp 1632082664
transform 1 0 51796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_571
timestamp 1632082664
transform 1 0 53636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_583
timestamp 1632082664
transform 1 0 54740 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_601
timestamp 1632082664
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_589
timestamp 1632082664
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1632082664
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1632082664
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_613
timestamp 1632082664
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_625
timestamp 1632082664
transform 1 0 58604 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_629
timestamp 1632082664
transform 1 0 58972 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1632082664
transform -1 0 59340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1632082664
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1632082664
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1632082664
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1364_
timestamp 1632082664
transform 1 0 3680 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_3_27
timestamp 1632082664
transform 1 0 3588 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1369_
timestamp 1632082664
transform 1 0 6348 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1632082664
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1632082664
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_73
timestamp 1632082664
transform 1 0 7820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_97
timestamp 1632082664
transform 1 0 10028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_85
timestamp 1632082664
transform 1 0 8924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1381_
timestamp 1632082664
transform 1 0 11500 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1632082664
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp 1632082664
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1384_
timestamp 1632082664
transform 1 0 13340 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_129
timestamp 1632082664
transform 1 0 12972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1632082664
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1632082664
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1390_
timestamp 1632082664
transform 1 0 16652 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1632082664
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1632082664
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_185
timestamp 1632082664
transform 1 0 18124 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_115_clk sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 18584 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1632082664
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1632082664
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1401_
timestamp 1632082664
transform 1 0 21804 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_3_210
timestamp 1632082664
transform 1 0 20424 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1632082664
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_241
timestamp 1632082664
transform 1 0 23276 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1738_
timestamp 1632082664
transform 1 0 24012 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_3_265
timestamp 1632082664
transform 1 0 25484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1732_
timestamp 1632082664
transform 1 0 26956 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1632082664
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_277
timestamp 1632082664
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_309
timestamp 1632082664
transform 1 0 29532 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1724_
timestamp 1632082664
transform 1 0 29716 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_3_297
timestamp 1632082664
transform 1 0 28428 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_327
timestamp 1632082664
transform 1 0 31188 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_337
timestamp 1632082664
transform 1 0 32108 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1719_
timestamp 1632082664
transform 1 0 32752 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1632082664
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_343
timestamp 1632082664
transform 1 0 32660 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1632082664
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 1632082664
transform 1 0 34592 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_360
timestamp 1632082664
transform 1 0 34224 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1855_
timestamp 1632082664
transform 1 0 37260 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_3_380
timestamp 1632082664
transform 1 0 36064 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1632082664
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1877_
timestamp 1632082664
transform 1 0 39100 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_409
timestamp 1632082664
transform 1 0 38732 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_429
timestamp 1632082664
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1632082664
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_449
timestamp 1632082664
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1632082664
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1632082664
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1610_
timestamp 1632082664
transform 1 0 43976 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_3_465
timestamp 1632082664
transform 1 0 43884 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_461
timestamp 1632082664
transform 1 0 43516 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_494
timestamp 1632082664
transform 1 0 46552 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_482
timestamp 1632082664
transform 1 0 45448 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_502
timestamp 1632082664
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1604_
timestamp 1632082664
transform 1 0 47564 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1632082664
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_521
timestamp 1632082664
transform 1 0 49036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1506_
timestamp 1632082664
transform 1 0 49864 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_3_529
timestamp 1632082664
transform 1 0 49772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_558
timestamp 1632082664
transform 1 0 52440 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1511_
timestamp 1632082664
transform 1 0 52716 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_3_546
timestamp 1632082664
transform 1 0 51336 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1632082664
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_577
timestamp 1632082664
transform 1 0 54188 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_601
timestamp 1632082664
transform 1 0 56396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_589
timestamp 1632082664
transform 1 0 55292 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_617
timestamp 1632082664
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1632082664
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_613
timestamp 1632082664
transform 1 0 57500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_629
timestamp 1632082664
transform 1 0 58972 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1632082664
transform -1 0 59340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1632082664
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1632082664
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1632082664
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1363_
timestamp 1632082664
transform 1 0 3772 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1632082664
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1632082664
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1365_
timestamp 1632082664
transform 1 0 5612 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_45
timestamp 1632082664
transform 1 0 5244 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1632082664
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1632082664
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1632082664
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1632082664
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1378_
timestamp 1632082664
transform 1 0 9752 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1632082664
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_93
timestamp 1632082664
transform 1 0 9660 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1379_
timestamp 1632082664
transform 1 0 11592 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_110
timestamp 1632082664
transform 1 0 11224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_130
timestamp 1632082664
transform 1 0 13064 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1632082664
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1388_
timestamp 1632082664
transform 1 0 14076 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1632082664
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1392_
timestamp 1632082664
transform 1 0 15916 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_157
timestamp 1632082664
transform 1 0 15548 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1632082664
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1632082664
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_197
timestamp 1632082664
transform 1 0 19228 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1400_
timestamp 1632082664
transform 1 0 20056 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1632082664
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_205
timestamp 1632082664
transform 1 0 19964 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1632082664
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1402_
timestamp 1632082664
transform 1 0 21896 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_222
timestamp 1632082664
transform 1 0 21528 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_242
timestamp 1632082664
transform 1 0 23368 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1632082664
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_253
timestamp 1632082664
transform 1 0 24380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1731_
timestamp 1632082664
transform 1 0 25116 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1632082664
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1730_
timestamp 1632082664
transform 1 0 26956 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_277
timestamp 1632082664
transform 1 0 26588 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_297
timestamp 1632082664
transform 1 0 28428 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1632082664
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_309
timestamp 1632082664
transform 1 0 29532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp 1632082664
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1723_
timestamp 1632082664
transform 1 0 29992 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_4_330
timestamp 1632082664
transform 1 0 31464 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_313
timestamp 1632082664
transform 1 0 29900 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_342
timestamp 1632082664
transform 1 0 32568 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1718_
timestamp 1632082664
transform 1 0 32752 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_4_365
timestamp 1632082664
transform 1 0 34684 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1613_
timestamp 1632082664
transform 1 0 35328 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1632082664
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_371
timestamp 1632082664
transform 1 0 35236 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_360
timestamp 1632082664
transform 1 0 34224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1833_
timestamp 1632082664
transform 1 0 37168 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_388
timestamp 1632082664
transform 1 0 36800 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_408
timestamp 1632082664
transform 1 0 38640 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1910_
timestamp 1632082664
transform 1 0 39836 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1632082664
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_437
timestamp 1632082664
transform 1 0 41308 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1954_
timestamp 1632082664
transform 1 0 41676 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_4_457
timestamp 1632082664
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1632082664
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1632082664
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1632082664
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1632082664
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_489
timestamp 1632082664
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1602_
timestamp 1632082664
transform 1 0 47564 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_501
timestamp 1632082664
transform 1 0 47196 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_521
timestamp 1632082664
transform 1 0 49036 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1505_
timestamp 1632082664
transform 1 0 50140 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1632082664
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_529
timestamp 1632082664
transform 1 0 49772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1510_
timestamp 1632082664
transform 1 0 51980 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_549
timestamp 1632082664
transform 1 0 51612 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1632082664
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_569
timestamp 1632082664
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_601
timestamp 1632082664
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_589
timestamp 1632082664
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1632082664
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1632082664
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_613
timestamp 1632082664
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_625
timestamp 1632082664
transform 1 0 58604 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_629
timestamp 1632082664
transform 1 0 58972 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1632082664
transform -1 0 59340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3
timestamp 1632082664
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1361_
timestamp 1632082664
transform 1 0 2392 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1632082664
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_11
timestamp 1632082664
transform 1 0 2116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1362_
timestamp 1632082664
transform 1 0 4232 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_30
timestamp 1632082664
transform 1 0 3864 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_50
timestamp 1632082664
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1368_
timestamp 1632082664
transform 1 0 6348 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1632082664
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_73
timestamp 1632082664
transform 1 0 7820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_104
timestamp 1632082664
transform 1 0 10672 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1376_
timestamp 1632082664
transform 1 0 9200 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_5_85
timestamp 1632082664
transform 1 0 8924 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_119_clk
timestamp 1632082664
transform 1 0 11960 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1632082664
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_117
timestamp 1632082664
transform 1 0 11868 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_113
timestamp 1632082664
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1385_
timestamp 1632082664
transform 1 0 14168 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_138
timestamp 1632082664
transform 1 0 13800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_158
timestamp 1632082664
transform 1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1632082664
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1632082664
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1632082664
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1632082664
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_193
timestamp 1632082664
transform 1 0 18860 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1740_
timestamp 1632082664
transform 1 0 19872 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_5_201
timestamp 1632082664
transform 1 0 19596 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1632082664
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1632082664
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1632082664
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_114_clk
timestamp 1632082664
transform 1 0 23368 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_5_241
timestamp 1632082664
transform 1 0 23276 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_237
timestamp 1632082664
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_262
timestamp 1632082664
transform 1 0 25208 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_274
timestamp 1632082664
transform 1 0 26312 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1632082664
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1632082664
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_113_clk
timestamp 1632082664
transform 1 0 28152 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_5_293
timestamp 1632082664
transform 1 0 28060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_326
timestamp 1632082664
transform 1 0 31096 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_314
timestamp 1632082664
transform 1 0 29992 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp 1632082664
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1717_
timestamp 1632082664
transform 1 0 32476 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1632082664
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_337
timestamp 1632082664
transform 1 0 32108 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1612_
timestamp 1632082664
transform 1 0 35144 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_5_357
timestamp 1632082664
transform 1 0 33948 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_369
timestamp 1632082664
transform 1 0 35052 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_386
timestamp 1632082664
transform 1 0 36616 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1632082664
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_393
timestamp 1632082664
transform 1 0 37260 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1899_
timestamp 1632082664
transform 1 0 37720 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_397
timestamp 1632082664
transform 1 0 37628 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_414
timestamp 1632082664
transform 1 0 39192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_97_clk
timestamp 1632082664
transform 1 0 39560 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_5_438
timestamp 1632082664
transform 1 0 41400 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_446
timestamp 1632082664
transform 1 0 42136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1632082664
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1632082664
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1607_
timestamp 1632082664
transform 1 0 43976 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_465
timestamp 1632082664
transform 1 0 43884 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_461
timestamp 1632082664
transform 1 0 43516 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_494
timestamp 1632082664
transform 1 0 46552 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_482
timestamp 1632082664
transform 1 0 45448 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_505
timestamp 1632082664
transform 1 0 47564 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1632082664
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1504_
timestamp 1632082664
transform 1 0 48300 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1632082664
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1503_
timestamp 1632082664
transform 1 0 50140 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_529
timestamp 1632082664
transform 1 0 49772 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_549
timestamp 1632082664
transform 1 0 51612 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1513_
timestamp 1632082664
transform 1 0 52808 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1632082664
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_561
timestamp 1632082664
transform 1 0 52716 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_557
timestamp 1632082664
transform 1 0 52348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_578
timestamp 1632082664
transform 1 0 54280 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_602
timestamp 1632082664
transform 1 0 56488 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_590
timestamp 1632082664
transform 1 0 55384 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_614
timestamp 1632082664
transform 1 0 57592 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_617
timestamp 1632082664
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1632082664
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_629
timestamp 1632082664
transform 1 0 58972 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1632082664
transform -1 0 59340 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1632082664
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1359_
timestamp 1632082664
transform 1 0 2024 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1632082664
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1632082664
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_9
timestamp 1632082664
transform 1 0 1932 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1632082664
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1632082664
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1632082664
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1360_
timestamp 1632082664
transform 1 0 3956 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1357_
timestamp 1632082664
transform 1 0 3864 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1632082664
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1632082664
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_26
timestamp 1632082664
transform 1 0 3496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_57
timestamp 1632082664
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_46
timestamp 1632082664
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1632082664
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1367_
timestamp 1632082664
transform 1 0 5796 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1632082664
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_47
timestamp 1632082664
transform 1 0 5428 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_120_clk
timestamp 1632082664
transform 1 0 7176 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_6_67
timestamp 1632082664
transform 1 0 7268 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_65
timestamp 1632082664
transform 1 0 7084 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1632082664
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1632082664
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1374_
timestamp 1632082664
transform 1 0 8924 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1372_
timestamp 1632082664
transform 1 0 9384 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1632082664
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_86
timestamp 1632082664
transform 1 0 9016 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_101
timestamp 1632082664
transform 1 0 10396 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_106
timestamp 1632082664
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1762_
timestamp 1632082664
transform 1 0 11868 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1377_
timestamp 1632082664
transform 1 0 10764 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1632082664
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1632082664
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 1632082664
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1632082664
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1389_
timestamp 1632082664
transform 1 0 14444 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_7_133
timestamp 1632082664
transform 1 0 13340 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1632082664
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1632082664
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1632082664
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_145
timestamp 1632082664
transform 1 0 14444 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1757_
timestamp 1632082664
transform 1 0 14720 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1754_
timestamp 1632082664
transform 1 0 16284 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1632082664
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_161
timestamp 1632082664
transform 1 0 15916 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1750_
timestamp 1632082664
transform 1 0 16928 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_6_181
timestamp 1632082664
transform 1 0 17756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1632082664
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_169
timestamp 1632082664
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1744_
timestamp 1632082664
transform 1 0 19504 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1743_
timestamp 1632082664
transform 1 0 19228 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_7_188
timestamp 1632082664
transform 1 0 18400 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1632082664
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 1632082664
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_216
timestamp 1632082664
transform 1 0 20976 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1404_
timestamp 1632082664
transform 1 0 22080 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1403_
timestamp 1632082664
transform 1 0 21804 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_6_213
timestamp 1632082664
transform 1 0 20700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1632082664
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp 1632082664
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_244
timestamp 1632082664
transform 1 0 23552 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_241
timestamp 1632082664
transform 1 0 23276 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1632082664
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp 1632082664
transform 1 0 25852 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1729_
timestamp 1632082664
transform 1 0 25760 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1406_
timestamp 1632082664
transform 1 0 24380 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1632082664
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1632082664
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_252
timestamp 1632082664
transform 1 0 24288 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_265
timestamp 1632082664
transform 1 0 25484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1728_
timestamp 1632082664
transform 1 0 26956 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1727_
timestamp 1632082664
transform 1 0 27600 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1632082664
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_284
timestamp 1632082664
transform 1 0 27232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_277
timestamp 1632082664
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_309
timestamp 1632082664
transform 1 0 29532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1722_
timestamp 1632082664
transform 1 0 29716 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1721_
timestamp 1632082664
transform 1 0 29532 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_7_297
timestamp 1632082664
transform 1 0 28428 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1632082664
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_304
timestamp 1632082664
transform 1 0 29072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_327
timestamp 1632082664
transform 1 0 31188 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_325
timestamp 1632082664
transform 1 0 31004 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_337
timestamp 1632082664
transform 1 0 32108 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1716_
timestamp 1632082664
transform 1 0 32660 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 1632082664
transform 1 0 32108 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_7_353
timestamp 1632082664
transform 1 0 33580 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1632082664
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1632082664
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_98_clk
timestamp 1632082664
transform 1 0 35052 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_7_365
timestamp 1632082664
transform 1 0 34684 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1614_
timestamp 1632082664
transform 1 0 35328 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1632082664
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_371
timestamp 1632082664
transform 1 0 35236 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1632082664
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_365
timestamp 1632082664
transform 1 0 34684 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_359
timestamp 1632082664
transform 1 0 34132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_393
timestamp 1632082664
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_389
timestamp 1632082664
transform 1 0 36892 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1632082664
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_388
timestamp 1632082664
transform 1 0 36800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1976_
timestamp 1632082664
transform 1 0 37904 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1943_
timestamp 1632082664
transform 1 0 37996 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_416
timestamp 1632082664
transform 1 0 39376 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_397
timestamp 1632082664
transform 1 0 37628 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_437
timestamp 1632082664
transform 1 0 41308 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1932_
timestamp 1632082664
transform 1 0 39836 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1921_
timestamp 1632082664
transform 1 0 40296 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1632082664
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_425
timestamp 1632082664
transform 1 0 40204 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_417
timestamp 1632082664
transform 1 0 39468 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_421
timestamp 1632082664
transform 1 0 39836 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_454
timestamp 1632082664
transform 1 0 42872 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1609_
timestamp 1632082664
transform 1 0 43056 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1632082664
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_442
timestamp 1632082664
transform 1 0 41768 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1632082664
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_445
timestamp 1632082664
transform 1 0 42044 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1608_
timestamp 1632082664
transform 1 0 43792 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1606_
timestamp 1632082664
transform 1 0 44988 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1632082664
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_472
timestamp 1632082664
transform 1 0 44528 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_461
timestamp 1632082664
transform 1 0 43516 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_93_clk
timestamp 1632082664
transform 1 0 46828 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1603_
timestamp 1632082664
transform 1 0 45632 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_7_500
timestamp 1632082664
transform 1 0 47104 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_480
timestamp 1632082664
transform 1 0 45264 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_493
timestamp 1632082664
transform 1 0 46460 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1599_
timestamp 1632082664
transform 1 0 47932 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_6_517
timestamp 1632082664
transform 1 0 48668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1632082664
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_505
timestamp 1632082664
transform 1 0 47564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1502_
timestamp 1632082664
transform 1 0 49772 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_6_533
timestamp 1632082664
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1632082664
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_525
timestamp 1632082664
transform 1 0 49404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_529
timestamp 1632082664
transform 1 0 49772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_92_clk
timestamp 1632082664
transform 1 0 51428 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_7_561
timestamp 1632082664
transform 1 0 52716 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_545
timestamp 1632082664
transform 1 0 51244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_545
timestamp 1632082664
transform 1 0 51244 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1632082664
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_557
timestamp 1632082664
transform 1 0 52348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_579
timestamp 1632082664
transform 1 0 54372 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1514_
timestamp 1632082664
transform 1 0 53268 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_7_583
timestamp 1632082664
transform 1 0 54740 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_567
timestamp 1632082664
transform 1 0 53268 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_595
timestamp 1632082664
transform 1 0 55844 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_601
timestamp 1632082664
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_589
timestamp 1632082664
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1632082664
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1632082664
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_607
timestamp 1632082664
transform 1 0 56948 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_617
timestamp 1632082664
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_613
timestamp 1632082664
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1632082664
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1632082664
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_625
timestamp 1632082664
transform 1 0 58604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_629
timestamp 1632082664
transform 1 0 58972 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_629
timestamp 1632082664
transform 1 0 58972 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1632082664
transform -1 0 59340 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1632082664
transform -1 0 59340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1358_
timestamp 1632082664
transform 1 0 1840 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp 1632082664
transform 1 0 1748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1632082664
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1632082664
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1632082664
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1632082664
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1632082664
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp 1632082664
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1353_
timestamp 1632082664
transform 1 0 5152 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_60
timestamp 1632082664
transform 1 0 6624 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1370_
timestamp 1632082664
transform 1 0 6992 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1632082664
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1375_
timestamp 1632082664
transform 1 0 8924 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_8_101
timestamp 1632082664
transform 1 0 10396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1632082664
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_113
timestamp 1632082664
transform 1 0 11500 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1760_
timestamp 1632082664
transform 1 0 12144 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_119
timestamp 1632082664
transform 1 0 12052 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_141
timestamp 1632082664
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1632082664
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1632082664
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1753_
timestamp 1632082664
transform 1 0 15088 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_8_149
timestamp 1632082664
transform 1 0 14812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_168
timestamp 1632082664
transform 1 0 16560 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1749_
timestamp 1632082664
transform 1 0 17296 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_8_197
timestamp 1632082664
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1745_
timestamp 1632082664
transform 1 0 19780 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1632082664
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1632082664
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_219
timestamp 1632082664
transform 1 0 21252 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1405_
timestamp 1632082664
transform 1 0 22448 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_231
timestamp 1632082664
transform 1 0 22356 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1632082664
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1407_
timestamp 1632082664
transform 1 0 24380 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_8_269
timestamp 1632082664
transform 1 0 25852 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1632082664
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_281
timestamp 1632082664
transform 1 0 26956 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1726_
timestamp 1632082664
transform 1 0 27600 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_287
timestamp 1632082664
transform 1 0 27508 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1632082664
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1632082664
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_304
timestamp 1632082664
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_321
timestamp 1632082664
transform 1 0 30636 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1713_
timestamp 1632082664
transform 1 0 30820 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 1632082664
transform 1 0 32660 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_339
timestamp 1632082664
transform 1 0 32292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1632082664
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1632082664
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1632082664
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_359
timestamp 1632082664
transform 1 0 34132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_377
timestamp 1632082664
transform 1 0 35788 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1615_
timestamp 1632082664
transform 1 0 35972 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_395
timestamp 1632082664
transform 1 0 37444 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1616_
timestamp 1632082664
transform 1 0 37812 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_415
timestamp 1632082664
transform 1 0 39284 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_421
timestamp 1632082664
transform 1 0 39836 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1485_
timestamp 1632082664
transform 1 0 40572 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1632082664
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1632082664
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_445
timestamp 1632082664
transform 1 0 42044 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1611_
timestamp 1632082664
transform 1 0 43056 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_8_453
timestamp 1632082664
transform 1 0 42780 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_477
timestamp 1632082664
transform 1 0 44988 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1632082664
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_472
timestamp 1632082664
transform 1 0 44528 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1600_
timestamp 1632082664
transform 1 0 45724 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1598_
timestamp 1632082664
transform 1 0 47564 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_501
timestamp 1632082664
transform 1 0 47196 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_521
timestamp 1632082664
transform 1 0 49036 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1500_
timestamp 1632082664
transform 1 0 50140 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1632082664
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_529
timestamp 1632082664
transform 1 0 49772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1515_
timestamp 1632082664
transform 1 0 52808 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_8_549
timestamp 1632082664
transform 1 0 51612 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_561
timestamp 1632082664
transform 1 0 52716 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_578
timestamp 1632082664
transform 1 0 54280 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_586
timestamp 1632082664
transform 1 0 55016 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1523_
timestamp 1632082664
transform 1 0 55292 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1632082664
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1526_
timestamp 1632082664
transform 1 0 57132 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_625
timestamp 1632082664
transform 1 0 58604 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_605
timestamp 1632082664
transform 1 0 56764 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_629
timestamp 1632082664
transform 1 0 58972 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1632082664
transform -1 0 59340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1632082664
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1356_
timestamp 1632082664
transform 1 0 2024 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_9
timestamp 1632082664
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1632082664
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_121_clk
timestamp 1632082664
transform 1 0 4048 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_9_26
timestamp 1632082664
transform 1 0 3496 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1371_
timestamp 1632082664
transform 1 0 6716 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1632082664
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1632082664
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1632082664
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1373_
timestamp 1632082664
transform 1 0 8556 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_77
timestamp 1632082664
transform 1 0 8188 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_97
timestamp 1632082664
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1632082664
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1632082664
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_125
timestamp 1632082664
transform 1 0 12604 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1632082664
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1759_
timestamp 1632082664
transform 1 0 12880 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_144
timestamp 1632082664
transform 1 0 14352 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1752_
timestamp 1632082664
transform 1 0 14720 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1632082664
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1748_
timestamp 1632082664
transform 1 0 17848 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1632082664
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1632082664
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_181
timestamp 1632082664
transform 1 0 17756 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1746_
timestamp 1632082664
transform 1 0 19688 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_198
timestamp 1632082664
transform 1 0 19320 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_218
timestamp 1632082664
transform 1 0 21160 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1632082664
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1632082664
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_237
timestamp 1632082664
transform 1 0 22908 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_245
timestamp 1632082664
transform 1 0 23644 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1408_
timestamp 1632082664
transform 1 0 23828 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_263
timestamp 1632082664
transform 1 0 25300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1704_
timestamp 1632082664
transform 1 0 26956 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1632082664
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1632082664
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp 1632082664
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1709_
timestamp 1632082664
transform 1 0 29532 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_297
timestamp 1632082664
transform 1 0 28428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_325
timestamp 1632082664
transform 1 0 31004 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 1632082664
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1712_
timestamp 1632082664
transform 1 0 32108 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_353
timestamp 1632082664
transform 1 0 33580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1632082664
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_365
timestamp 1632082664
transform 1 0 34684 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1617_
timestamp 1632082664
transform 1 0 35328 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_371
timestamp 1632082664
transform 1 0 35236 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1632082664
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1632082664
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_388
timestamp 1632082664
transform 1 0 36800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1483_
timestamp 1632082664
transform 1 0 38640 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_9_405
timestamp 1632082664
transform 1 0 38364 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0000_
timestamp 1632082664
transform 1 0 40480 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_424
timestamp 1632082664
transform 1 0 40112 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1488_
timestamp 1632082664
transform 1 0 42780 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1632082664
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_449
timestamp 1632082664
transform 1 0 42412 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_444
timestamp 1632082664
transform 1 0 41952 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_469
timestamp 1632082664
transform 1 0 44252 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1601_
timestamp 1632082664
transform 1 0 45632 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_500
timestamp 1632082664
transform 1 0 47104 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_481
timestamp 1632082664
transform 1 0 45356 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1498_
timestamp 1632082664
transform 1 0 48944 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_505
timestamp 1632082664
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1632082664
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_517
timestamp 1632082664
transform 1 0 48668 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1501_
timestamp 1632082664
transform 1 0 50784 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_536
timestamp 1632082664
transform 1 0 50416 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1516_
timestamp 1632082664
transform 1 0 52716 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1632082664
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_556
timestamp 1632082664
transform 1 0 52256 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1520_
timestamp 1632082664
transform 1 0 54556 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_577
timestamp 1632082664
transform 1 0 54188 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_597
timestamp 1632082664
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1632082664
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_617
timestamp 1632082664
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1632082664
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1632082664
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_629
timestamp 1632082664
transform 1 0 58972 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1632082664
transform -1 0 59340 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1355_
timestamp 1632082664
transform 1 0 1840 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1632082664
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1632082664
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1632082664
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1354_
timestamp 1632082664
transform 1 0 4048 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1632082664
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1632082664
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 1632082664
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1350_
timestamp 1632082664
transform 1 0 5888 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_48
timestamp 1632082664
transform 1 0 5520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1632082664
transform 1 0 7360 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1632082664
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1763_
timestamp 1632082664
transform 1 0 10304 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1632082664
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1632082664
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_97
timestamp 1632082664
transform 1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1761_
timestamp 1632082664
transform 1 0 12144 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_116
timestamp 1632082664
transform 1 0 11776 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1755_
timestamp 1632082664
transform 1 0 14444 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1632082664
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1632082664
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1632082664
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1751_
timestamp 1632082664
transform 1 0 16284 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_161
timestamp 1632082664
transform 1 0 15916 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_181
timestamp 1632082664
transform 1 0 17756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1747_
timestamp 1632082664
transform 1 0 19320 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1632082664
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_197
timestamp 1632082664
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1632082664
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_214
timestamp 1632082664
transform 1 0 20792 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1414_
timestamp 1632082664
transform 1 0 21620 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_222
timestamp 1632082664
transform 1 0 21528 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1632082664
transform 1 0 23092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1409_
timestamp 1632082664
transform 1 0 24380 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1632082664
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1632082664
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_269
timestamp 1632082664
transform 1 0 25852 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1701_
timestamp 1632082664
transform 1 0 26220 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1632082664
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1632082664
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1707_
timestamp 1632082664
transform 1 0 29532 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1632082664
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1632082664
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_325
timestamp 1632082664
transform 1 0 31004 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_353
timestamp 1632082664
transform 1 0 33580 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1711_
timestamp 1632082664
transform 1 0 32108 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1477_
timestamp 1632082664
transform 1 0 34684 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1632082664
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_361
timestamp 1632082664
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_393
timestamp 1632082664
transform 1 0 37260 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1481_
timestamp 1632082664
transform 1 0 37444 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_10_381
timestamp 1632082664
transform 1 0 36156 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_411
timestamp 1632082664
transform 1 0 38916 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_433
timestamp 1632082664
transform 1 0 40940 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1632082664
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1632082664
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1632082664
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_96_clk
timestamp 1632082664
transform 1 0 41768 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_10_441
timestamp 1632082664
transform 1 0 41676 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_474
timestamp 1632082664
transform 1 0 44712 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1493_
timestamp 1632082664
transform 1 0 44988 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_10_462
timestamp 1632082664
transform 1 0 43608 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1632082664
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1495_
timestamp 1632082664
transform 1 0 46828 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_493
timestamp 1632082664
transform 1 0 46460 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_513
timestamp 1632082664
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1632082664
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1499_
timestamp 1632082664
transform 1 0 50140 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1632082664
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1632082664
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1517_
timestamp 1632082664
transform 1 0 52716 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_10_549
timestamp 1632082664
transform 1 0 51612 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_577
timestamp 1632082664
transform 1 0 54188 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1521_
timestamp 1632082664
transform 1 0 55292 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1632082664
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_585
timestamp 1632082664
transform 1 0 54924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1524_
timestamp 1632082664
transform 1 0 57132 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_625
timestamp 1632082664
transform 1 0 58604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_605
timestamp 1632082664
transform 1 0 56764 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_629
timestamp 1632082664
transform 1 0 58972 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1632082664
transform -1 0 59340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1632082664
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1632082664
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1632082664
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_27
timestamp 1632082664
transform 1 0 3588 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1352_
timestamp 1632082664
transform 1 0 4416 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_35
timestamp 1632082664
transform 1 0 4324 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1349_
timestamp 1632082664
transform 1 0 6348 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1632082664
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1632082664
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_73
timestamp 1632082664
transform 1 0 7820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_102
timestamp 1632082664
transform 1 0 10488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1343_
timestamp 1632082664
transform 1 0 9016 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_85
timestamp 1632082664
transform 1 0 8924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1632082664
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1632082664
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1345_
timestamp 1632082664
transform 1 0 12236 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1632082664
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_137
timestamp 1632082664
transform 1 0 13708 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1758_
timestamp 1632082664
transform 1 0 14260 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_11_159
timestamp 1632082664
transform 1 0 15732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1632082664
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1632082664
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1632082664
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1632082664
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1416_
timestamp 1632082664
transform 1 0 19136 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_11_193
timestamp 1632082664
transform 1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1632082664
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1412_
timestamp 1632082664
transform 1 0 21988 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_11_212
timestamp 1632082664
transform 1 0 20608 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1632082664
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1410_
timestamp 1632082664
transform 1 0 23828 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_243
timestamp 1632082664
transform 1 0 23460 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_263
timestamp 1632082664
transform 1 0 25300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1702_
timestamp 1632082664
transform 1 0 26956 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1632082664
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1632082664
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_275
timestamp 1632082664
transform 1 0 26404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1703_
timestamp 1632082664
transform 1 0 28796 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_297
timestamp 1632082664
transform 1 0 28428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1632082664
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1632082664
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_349
timestamp 1632082664
transform 1 0 33212 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1475_
timestamp 1632082664
transform 1 0 33396 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1632082664
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1632082664
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1632082664
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1478_
timestamp 1632082664
transform 1 0 35236 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_367
timestamp 1632082664
transform 1 0 34868 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1480_
timestamp 1632082664
transform 1 0 37260 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1632082664
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1632082664
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_387
timestamp 1632082664
transform 1 0 36708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1482_
timestamp 1632082664
transform 1 0 39100 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_409
timestamp 1632082664
transform 1 0 38732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1632082664
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1632082664
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1484_
timestamp 1632082664
transform 1 0 42412 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1632082664
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1632082664
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1490_
timestamp 1632082664
transform 1 0 44252 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_465
timestamp 1632082664
transform 1 0 43884 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1632082664
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1632082664
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1496_
timestamp 1632082664
transform 1 0 47564 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1632082664
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1632082664
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1497_
timestamp 1632082664
transform 1 0 49404 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_11_541
timestamp 1632082664
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_521
timestamp 1632082664
transform 1 0 49036 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1632082664
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1518_
timestamp 1632082664
transform 1 0 52716 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1632082664
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1632082664
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_577
timestamp 1632082664
transform 1 0 54188 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_583
timestamp 1632082664
transform 1 0 54740 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_91_clk
timestamp 1632082664
transform 1 0 54832 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_11_604
timestamp 1632082664
transform 1 0 56672 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_617
timestamp 1632082664
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1632082664
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_629
timestamp 1632082664
transform 1 0 58972 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1632082664
transform -1 0 59340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1632082664
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1632082664
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1632082664
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1351_
timestamp 1632082664
transform 1 0 4048 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1632082664
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1632082664
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_29
timestamp 1632082664
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1347_
timestamp 1632082664
transform 1 0 5888 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_48
timestamp 1632082664
transform 1 0 5520 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1632082664
transform 1 0 7360 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1632082664
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1341_
timestamp 1632082664
transform 1 0 8924 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1632082664
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_101
timestamp 1632082664
transform 1 0 10396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1344_
timestamp 1632082664
transform 1 0 10764 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1632082664
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1632082664
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1765_
timestamp 1632082664
transform 1 0 14076 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1632082664
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1632082664
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_157
timestamp 1632082664
transform 1 0 15548 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_181
timestamp 1632082664
transform 1 0 17756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_169
timestamp 1632082664
transform 1 0 16652 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1632082664
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1632082664
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_193
timestamp 1632082664
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1415_
timestamp 1632082664
transform 1 0 20332 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1413_
timestamp 1632082664
transform 1 0 22172 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_225
timestamp 1632082664
transform 1 0 21804 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1632082664
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1697_
timestamp 1632082664
transform 1 0 24380 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1632082664
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1632082664
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_269
timestamp 1632082664
transform 1 0 25852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1699_
timestamp 1632082664
transform 1 0 26220 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1632082664
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1632082664
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1708_
timestamp 1632082664
transform 1 0 29532 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1632082664
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1632082664
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_325
timestamp 1632082664
transform 1 0 31004 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_99_clk
timestamp 1632082664
transform 1 0 32384 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_12_337
timestamp 1632082664
transform 1 0 32108 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1476_
timestamp 1632082664
transform 1 0 34684 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1632082664
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_360
timestamp 1632082664
transform 1 0 34224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1479_
timestamp 1632082664
transform 1 0 36524 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_381
timestamp 1632082664
transform 1 0 36156 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1632082664
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1632082664
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_421
timestamp 1632082664
transform 1 0 39836 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0011_
timestamp 1632082664
transform 1 0 40664 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1632082664
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_429
timestamp 1632082664
transform 1 0 40572 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1632082664
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1486_
timestamp 1632082664
transform 1 0 42504 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_446
timestamp 1632082664
transform 1 0 42136 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_466
timestamp 1632082664
transform 1 0 43976 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_474
timestamp 1632082664
transform 1 0 44712 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1489_
timestamp 1632082664
transform 1 0 44988 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1632082664
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1494_
timestamp 1632082664
transform 1 0 46828 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_493
timestamp 1632082664
transform 1 0 46460 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_513
timestamp 1632082664
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1632082664
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_533
timestamp 1632082664
transform 1 0 50140 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1632082664
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1632082664
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_541
timestamp 1632082664
transform 1 0 50876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1583_
timestamp 1632082664
transform 1 0 51152 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_560
timestamp 1632082664
transform 1 0 52624 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_580
timestamp 1632082664
transform 1 0 54464 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1519_
timestamp 1632082664
transform 1 0 52992 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1522_
timestamp 1632082664
transform 1 0 55292 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1632082664
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1525_
timestamp 1632082664
transform 1 0 57132 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_625
timestamp 1632082664
transform 1 0 58604 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_605
timestamp 1632082664
transform 1 0 56764 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_629
timestamp 1632082664
transform 1 0 58972 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1632082664
transform -1 0 59340 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1632082664
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1632082664
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1632082664
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1632082664
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1632082664
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1632082664
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1632082664
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1632082664
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1632082664
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1632082664
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1632082664
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1632082664
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1348_
timestamp 1632082664
transform 1 0 6072 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1346_
timestamp 1632082664
transform 1 0 6348 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1632082664
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_53
timestamp 1632082664
transform 1 0 5980 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1632082664
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1632082664
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1632082664
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_70
timestamp 1632082664
transform 1 0 7544 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_73
timestamp 1632082664
transform 1 0 7820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_102
timestamp 1632082664
transform 1 0 10488 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1632082664
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1340_
timestamp 1632082664
transform 1 0 9016 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1339_
timestamp 1632082664
transform 1 0 9108 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1632082664
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_85
timestamp 1632082664
transform 1 0 8924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_103
timestamp 1632082664
transform 1 0 10580 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1632082664
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1342_
timestamp 1632082664
transform 1 0 10948 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_14_123
timestamp 1632082664
transform 1 0 12420 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1632082664
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1632082664
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_125
timestamp 1632082664
transform 1 0 12604 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_118_clk
timestamp 1632082664
transform 1 0 12880 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_14_141
timestamp 1632082664
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1632082664
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1632082664
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_135
timestamp 1632082664
transform 1 0 13524 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp 1632082664
transform 1 0 15824 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1766_
timestamp 1632082664
transform 1 0 14720 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_13_148
timestamp 1632082664
transform 1 0 14720 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_147
timestamp 1632082664
transform 1 0 14628 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_164
timestamp 1632082664
transform 1 0 16192 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1780_
timestamp 1632082664
transform 1 0 16652 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1777_
timestamp 1632082664
transform 1 0 16560 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_14_184
timestamp 1632082664
transform 1 0 18032 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_185
timestamp 1632082664
transform 1 0 18124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1632082664
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_116_clk
timestamp 1632082664
transform 1 0 19596 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1417_
timestamp 1632082664
transform 1 0 19320 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1632082664
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_197
timestamp 1632082664
transform 1 0 19228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1632082664
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_214
timestamp 1632082664
transform 1 0 20792 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1632082664
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1632082664
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1632082664
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1632082664
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1632082664
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1411_
timestamp 1632082664
transform 1 0 23184 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1632082664
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_237
timestamp 1632082664
transform 1 0 22908 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_269
timestamp 1632082664
transform 1 0 25852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1698_
timestamp 1632082664
transform 1 0 25024 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1696_
timestamp 1632082664
transform 1 0 24380 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1632082664
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1632082664
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_256
timestamp 1632082664
transform 1 0 24656 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_112_clk
timestamp 1632082664
transform 1 0 26680 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1700_
timestamp 1632082664
transform 1 0 26956 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1632082664
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_277
timestamp 1632082664
transform 1 0 26588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1632082664
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_298
timestamp 1632082664
transform 1 0 28520 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1632082664
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1710_
timestamp 1632082664
transform 1 0 29532 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1705_
timestamp 1632082664
transform 1 0 28796 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1632082664
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_297
timestamp 1632082664
transform 1 0 28428 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1632082664
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_325
timestamp 1632082664
transform 1 0 31004 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1632082664
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_337
timestamp 1632082664
transform 1 0 32108 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_349
timestamp 1632082664
transform 1 0 33212 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1474_
timestamp 1632082664
transform 1 0 32752 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1632082664
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1632082664
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_343
timestamp 1632082664
transform 1 0 32660 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1632082664
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1473_
timestamp 1632082664
transform 1 0 33764 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1632082664
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_371
timestamp 1632082664
transform 1 0 35236 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1632082664
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_360
timestamp 1632082664
transform 1 0 34224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_383
timestamp 1632082664
transform 1 0 36340 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1619_
timestamp 1632082664
transform 1 0 37168 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1618_
timestamp 1632082664
transform 1 0 37260 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1632082664
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1632082664
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1632082664
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_389
timestamp 1632082664
transform 1 0 36892 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_408
timestamp 1632082664
transform 1 0 38640 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_409
timestamp 1632082664
transform 1 0 38732 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_421
timestamp 1632082664
transform 1 0 39836 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0022_
timestamp 1632082664
transform 1 0 40480 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1632082664
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1632082664
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1632082664
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_427
timestamp 1632082664
transform 1 0 40388 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_445
timestamp 1632082664
transform 1 0 42044 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1597_
timestamp 1632082664
transform 1 0 43056 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1487_
timestamp 1632082664
transform 1 0 42412 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1632082664
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_444
timestamp 1632082664
transform 1 0 41952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_453
timestamp 1632082664
transform 1 0 42780 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1492_
timestamp 1632082664
transform 1 0 44988 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1491_
timestamp 1632082664
transform 1 0 44252 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1632082664
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_472
timestamp 1632082664
transform 1 0 44528 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_465
timestamp 1632082664
transform 1 0 43884 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1632082664
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_493
timestamp 1632082664
transform 1 0 46460 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1632082664
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_94_clk
timestamp 1632082664
transform 1 0 47288 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1586_
timestamp 1632082664
transform 1 0 48944 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_13_505
timestamp 1632082664
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1632082664
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_501
timestamp 1632082664
transform 1 0 47196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1632082664
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_517
timestamp 1632082664
transform 1 0 48668 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_522
timestamp 1632082664
transform 1 0 49128 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_530
timestamp 1632082664
transform 1 0 49864 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1584_
timestamp 1632082664
transform 1 0 50784 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_14_533
timestamp 1632082664
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1632082664
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_536
timestamp 1632082664
transform 1 0 50416 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_561
timestamp 1632082664
transform 1 0 52716 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1581_
timestamp 1632082664
transform 1 0 51520 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1632082664
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_556
timestamp 1632082664
transform 1 0 52256 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_545
timestamp 1632082664
transform 1 0 51244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1580_
timestamp 1632082664
transform 1 0 53360 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1577_
timestamp 1632082664
transform 1 0 53360 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_13_567
timestamp 1632082664
transform 1 0 53268 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_564
timestamp 1632082664
transform 1 0 52992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1528_
timestamp 1632082664
transform 1 0 55936 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_14_589
timestamp 1632082664
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_584
timestamp 1632082664
transform 1 0 54832 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1632082664
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_601
timestamp 1632082664
transform 1 0 56396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_584
timestamp 1632082664
transform 1 0 54832 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_622
timestamp 1632082664
transform 1 0 58328 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1527_
timestamp 1632082664
transform 1 0 56856 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_13_617
timestamp 1632082664
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1632082664
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_605
timestamp 1632082664
transform 1 0 56764 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_612
timestamp 1632082664
transform 1 0 57408 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_629
timestamp 1632082664
transform 1 0 58972 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1632082664
transform -1 0 59340 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1632082664
transform -1 0 59340 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1632082664
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1632082664
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1632082664
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1632082664
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1632082664
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1632082664
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1632082664
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1632082664
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1632082664
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_81
timestamp 1632082664
transform 1 0 8556 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1632082664
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1338_
timestamp 1632082664
transform 1 0 9292 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1632082664
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1764_
timestamp 1632082664
transform 1 0 11500 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1632082664
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1632082664
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1769_
timestamp 1632082664
transform 1 0 14076 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_15_129
timestamp 1632082664
transform 1 0 12972 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_157
timestamp 1632082664
transform 1 0 15548 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 1632082664
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_185
timestamp 1632082664
transform 1 0 18124 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1776_
timestamp 1632082664
transform 1 0 16652 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1632082664
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_clk
timestamp 1632082664
transform 1 0 18952 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1418_
timestamp 1632082664
transform 1 0 19596 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_193
timestamp 1632082664
transform 1 0 18860 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_197
timestamp 1632082664
transform 1 0 19228 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1632082664
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1421_
timestamp 1632082664
transform 1 0 21804 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1632082664
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1632082664
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_241
timestamp 1632082664
transform 1 0 23276 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1695_
timestamp 1632082664
transform 1 0 24012 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_15_265
timestamp 1632082664
transform 1 0 25484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_281
timestamp 1632082664
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1706_
timestamp 1632082664
transform 1 0 27600 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1632082664
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_287
timestamp 1632082664
transform 1 0 27508 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1632082664
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_304
timestamp 1632082664
transform 1 0 29072 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_328
timestamp 1632082664
transform 1 0 31280 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_316
timestamp 1632082664
transform 1 0 30176 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1676_
timestamp 1632082664
transform 1 0 32384 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1632082664
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_337
timestamp 1632082664
transform 1 0 32108 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1472_
timestamp 1632082664
transform 1 0 34224 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_356
timestamp 1632082664
transform 1 0 33856 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1620_
timestamp 1632082664
transform 1 0 37260 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_15_376
timestamp 1632082664
transform 1 0 35696 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1632082664
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_388
timestamp 1632082664
transform 1 0 36800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_409
timestamp 1632082664
transform 1 0 38732 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_421
timestamp 1632082664
transform 1 0 39836 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0033_
timestamp 1632082664
transform 1 0 40480 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_427
timestamp 1632082664
transform 1 0 40388 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1632082664
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1632082664
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_444
timestamp 1632082664
transform 1 0 41952 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1596_
timestamp 1632082664
transform 1 0 43792 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_15_461
timestamp 1632082664
transform 1 0 43516 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1595_
timestamp 1632082664
transform 1 0 45632 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1632082664
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_480
timestamp 1632082664
transform 1 0 45264 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_clk
timestamp 1632082664
transform 1 0 48208 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_505
timestamp 1632082664
transform 1 0 47564 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1587_
timestamp 1632082664
transform 1 0 48944 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1632082664
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_519
timestamp 1632082664
transform 1 0 48852 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_511
timestamp 1632082664
transform 1 0 48116 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_515
timestamp 1632082664
transform 1 0 48484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1582_
timestamp 1632082664
transform 1 0 50784 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_536
timestamp 1632082664
transform 1 0 50416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_561
timestamp 1632082664
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1632082664
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_556
timestamp 1632082664
transform 1 0 52256 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1532_
timestamp 1632082664
transform 1 0 54096 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_15_573
timestamp 1632082664
transform 1 0 53820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1530_
timestamp 1632082664
transform 1 0 55936 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_592
timestamp 1632082664
transform 1 0 55568 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_617
timestamp 1632082664
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1632082664
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_612
timestamp 1632082664
transform 1 0 57408 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_629
timestamp 1632082664
transform 1 0 58972 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1632082664
transform -1 0 59340 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1632082664
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1632082664
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1632082664
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_29
timestamp 1632082664
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1287_
timestamp 1632082664
transform 1 0 4416 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1632082664
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_35
timestamp 1632082664
transform 1 0 4324 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1632082664
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_52
timestamp 1632082664
transform 1 0 5888 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_76
timestamp 1632082664
transform 1 0 8096 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_64
timestamp 1632082664
transform 1 0 6992 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1337_
timestamp 1632082664
transform 1 0 9384 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1632082664
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_89
timestamp 1632082664
transform 1 0 9292 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1632082664
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_clk
timestamp 1632082664
transform 1 0 11500 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_106
timestamp 1632082664
transform 1 0 10856 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1768_
timestamp 1632082664
transform 1 0 12144 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_112
timestamp 1632082664
transform 1 0 11408 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_116
timestamp 1632082664
transform 1 0 11776 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1770_
timestamp 1632082664
transform 1 0 14076 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1632082664
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1632082664
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1773_
timestamp 1632082664
transform 1 0 15916 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_157
timestamp 1632082664
transform 1 0 15548 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1632082664
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_197
timestamp 1632082664
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1632082664
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1419_
timestamp 1632082664
transform 1 0 19872 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1632082664
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_203
timestamp 1632082664
transform 1 0 19780 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1632082664
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_220
timestamp 1632082664
transform 1 0 21344 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1422_
timestamp 1632082664
transform 1 0 22080 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_16_244
timestamp 1632082664
transform 1 0 23552 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1694_
timestamp 1632082664
transform 1 0 24380 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_16_269
timestamp 1632082664
transform 1 0 25852 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1632082664
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_281
timestamp 1632082664
transform 1 0 26956 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_309
timestamp 1632082664
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_293
timestamp 1632082664
transform 1 0 28060 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1632082664
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_305
timestamp 1632082664
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1463_
timestamp 1632082664
transform 1 0 30544 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_317
timestamp 1632082664
transform 1 0 30268 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1467_
timestamp 1632082664
transform 1 0 32384 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_336
timestamp 1632082664
transform 1 0 32016 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_356
timestamp 1632082664
transform 1 0 33856 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1470_
timestamp 1632082664
transform 1 0 34684 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1632082664
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1621_
timestamp 1632082664
transform 1 0 37352 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_16_381
timestamp 1632082664
transform 1 0 36156 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_393
timestamp 1632082664
transform 1 0 37260 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_410
timestamp 1632082664
transform 1 0 38824 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_clk
timestamp 1632082664
transform 1 0 39836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_418
timestamp 1632082664
transform 1 0 39560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0044_
timestamp 1632082664
transform 1 0 40480 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1632082664
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_424
timestamp 1632082664
transform 1 0 40112 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_456
timestamp 1632082664
transform 1 0 43056 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_444
timestamp 1632082664
transform 1 0 41952 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_468
timestamp 1632082664
transform 1 0 44160 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1632082664
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1632082664
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1594_
timestamp 1632082664
transform 1 0 46368 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_489
timestamp 1632082664
transform 1 0 46092 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1590_
timestamp 1632082664
transform 1 0 48208 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_508
timestamp 1632082664
transform 1 0 47840 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_533
timestamp 1632082664
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1632082664
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_528
timestamp 1632082664
transform 1 0 49680 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1578_
timestamp 1632082664
transform 1 0 51520 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_545
timestamp 1632082664
transform 1 0 51244 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1576_
timestamp 1632082664
transform 1 0 53360 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_564
timestamp 1632082664
transform 1 0 52992 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_589
timestamp 1632082664
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1632082664
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_601
timestamp 1632082664
transform 1 0 56396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_584
timestamp 1632082664
transform 1 0 54832 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_622
timestamp 1632082664
transform 1 0 58328 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1529_
timestamp 1632082664
transform 1 0 56856 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_605
timestamp 1632082664
transform 1 0 56764 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1632082664
transform -1 0 59340 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1284_
timestamp 1632082664
transform 1 0 2852 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1632082664
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_15
timestamp 1632082664
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1632082664
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_35
timestamp 1632082664
transform 1 0 4324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1632082664
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1289_
timestamp 1632082664
transform 1 0 6348 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1632082664
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1632082664
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_73
timestamp 1632082664
transform 1 0 7820 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1336_
timestamp 1632082664
transform 1 0 9384 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_89
timestamp 1632082664
transform 1 0 9292 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_85
timestamp 1632082664
transform 1 0 8924 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1632082664
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_106
timestamp 1632082664
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1771_
timestamp 1632082664
transform 1 0 12144 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1632082664
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_119
timestamp 1632082664
transform 1 0 12052 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1772_
timestamp 1632082664
transform 1 0 13984 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_136
timestamp 1632082664
transform 1 0 13616 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_156
timestamp 1632082664
transform 1 0 15456 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1775_
timestamp 1632082664
transform 1 0 16652 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_17_185
timestamp 1632082664
transform 1 0 18124 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1632082664
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_197
timestamp 1632082664
transform 1 0 19228 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1420_
timestamp 1632082664
transform 1 0 19872 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_203
timestamp 1632082664
transform 1 0 19780 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1782_
timestamp 1632082664
transform 1 0 21804 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1632082664
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1632082664
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_241
timestamp 1632082664
transform 1 0 23276 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1693_
timestamp 1632082664
transform 1 0 24104 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_249
timestamp 1632082664
transform 1 0 24012 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_266
timestamp 1632082664
transform 1 0 25576 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_281
timestamp 1632082664
transform 1 0 26956 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_289
timestamp 1632082664
transform 1 0 27692 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1632082664
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1458_
timestamp 1632082664
transform 1 0 27876 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1632082664
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1461_
timestamp 1632082664
transform 1 0 29716 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_307
timestamp 1632082664
transform 1 0 29348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_327
timestamp 1632082664
transform 1 0 31188 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1465_
timestamp 1632082664
transform 1 0 32108 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1632082664
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1632082664
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_353
timestamp 1632082664
transform 1 0 33580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1469_
timestamp 1632082664
transform 1 0 33948 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1632082664
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1632082664
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1632082664
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1622_
timestamp 1632082664
transform 1 0 37444 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1632082664
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1632082664
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_411
timestamp 1632082664
transform 1 0 38916 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0055_
timestamp 1632082664
transform 1 0 40480 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_427
timestamp 1632082664
transform 1 0 40388 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_423
timestamp 1632082664
transform 1 0 40020 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0110_
timestamp 1632082664
transform 1 0 42412 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1632082664
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_444
timestamp 1632082664
transform 1 0 41952 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0143_
timestamp 1632082664
transform 1 0 44252 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_465
timestamp 1632082664
transform 1 0 43884 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1632082664
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1632082664
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1591_
timestamp 1632082664
transform 1 0 48944 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_17_505
timestamp 1632082664
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1632082664
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1632082664
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_517
timestamp 1632082664
transform 1 0 48668 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1585_
timestamp 1632082664
transform 1 0 50784 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_536
timestamp 1632082664
transform 1 0 50416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_561
timestamp 1632082664
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1632082664
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_556
timestamp 1632082664
transform 1 0 52256 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1535_
timestamp 1632082664
transform 1 0 54096 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_573
timestamp 1632082664
transform 1 0 53820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1531_
timestamp 1632082664
transform 1 0 55936 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_592
timestamp 1632082664
transform 1 0 55568 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1632082664
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output5
timestamp 1632082664
transform 1 0 58328 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_621
timestamp 1632082664
transform 1 0 58236 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_617
timestamp 1632082664
transform 1 0 57868 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_612
timestamp 1632082664
transform 1 0 57408 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_626
timestamp 1632082664
transform 1 0 58696 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1632082664
transform -1 0 59340 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1632082664
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1632082664
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1632082664
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1285_
timestamp 1632082664
transform 1 0 3772 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1632082664
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1632082664
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1286_
timestamp 1632082664
transform 1 0 5612 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_45
timestamp 1632082664
transform 1 0 5244 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1632082664
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1632082664
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1632082664
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1335_
timestamp 1632082664
transform 1 0 9384 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1632082664
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_89
timestamp 1632082664
transform 1 0 9292 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1632082664
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_118
timestamp 1632082664
transform 1 0 11960 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_106
timestamp 1632082664
transform 1 0 10856 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_130
timestamp 1632082664
transform 1 0 13064 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1632082664
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1326_
timestamp 1632082664
transform 1 0 14076 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1632082664
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1774_
timestamp 1632082664
transform 1 0 15916 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_157
timestamp 1632082664
transform 1 0 15548 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1632082664
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1632082664
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1632082664
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1632082664
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1632082664
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_209
timestamp 1632082664
transform 1 0 20332 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1423_
timestamp 1632082664
transform 1 0 20884 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_243
timestamp 1632082664
transform 1 0 23460 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_231
timestamp 1632082664
transform 1 0 22356 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1692_
timestamp 1632082664
transform 1 0 24380 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_18_269
timestamp 1632082664
transform 1 0 25852 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1632082664
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1632082664
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1456_
timestamp 1632082664
transform 1 0 27416 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_285
timestamp 1632082664
transform 1 0 27324 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_281
timestamp 1632082664
transform 1 0 26956 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_302
timestamp 1632082664
transform 1 0 28888 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1460_
timestamp 1632082664
transform 1 0 29532 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1632082664
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1462_
timestamp 1632082664
transform 1 0 31372 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_325
timestamp 1632082664
transform 1 0 31004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1632082664
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1632082664
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1471_
timestamp 1632082664
transform 1 0 34684 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1632082664
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1632082664
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_381
timestamp 1632082664
transform 1 0 36156 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_393
timestamp 1632082664
transform 1 0 37260 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_412
timestamp 1632082664
transform 1 0 39008 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1623_
timestamp 1632082664
transform 1 0 37536 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_421
timestamp 1632082664
transform 1 0 39836 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0066_
timestamp 1632082664
transform 1 0 40664 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1632082664
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_429
timestamp 1632082664
transform 1 0 40572 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0077_
timestamp 1632082664
transform 1 0 42504 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_446
timestamp 1632082664
transform 1 0 42136 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_466
timestamp 1632082664
transform 1 0 43976 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_474
timestamp 1632082664
transform 1 0 44712 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1632082664
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1632082664
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1593_
timestamp 1632082664
transform 1 0 46368 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_489
timestamp 1632082664
transform 1 0 46092 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1592_
timestamp 1632082664
transform 1 0 48208 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_508
timestamp 1632082664
transform 1 0 47840 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_533
timestamp 1632082664
transform 1 0 50140 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1632082664
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_528
timestamp 1632082664
transform 1 0 49680 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_541
timestamp 1632082664
transform 1 0 50876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1579_
timestamp 1632082664
transform 1 0 51152 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_560
timestamp 1632082664
transform 1 0 52624 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_580
timestamp 1632082664
transform 1 0 54464 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1575_
timestamp 1632082664
transform 1 0 52992 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1534_
timestamp 1632082664
transform 1 0 55384 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1632082664
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_589
timestamp 1632082664
transform 1 0 55292 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1183_
timestamp 1632082664
transform 1 0 57224 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_606
timestamp 1632082664
transform 1 0 56856 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_626
timestamp 1632082664
transform 1 0 58696 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1632082664
transform -1 0 59340 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1632082664
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1282_
timestamp 1632082664
transform 1 0 2116 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1281_
timestamp 1632082664
transform 1 0 1840 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1632082664
transform 1 0 1748 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1632082664
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1632082664
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1632082664
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1283_
timestamp 1632082664
transform 1 0 3956 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1632082664
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1632082664
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_41
timestamp 1632082664
transform 1 0 4876 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1632082664
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_27
timestamp 1632082664
transform 1 0 3588 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1632082664
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1291_
timestamp 1632082664
transform 1 0 6808 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1290_
timestamp 1632082664
transform 1 0 6348 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1288_
timestamp 1632082664
transform 1 0 4968 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1632082664
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1632082664
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_58
timestamp 1632082664
transform 1 0 6440 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_78
timestamp 1632082664
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_73
timestamp 1632082664
transform 1 0 7820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_85
timestamp 1632082664
transform 1 0 8924 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1333_
timestamp 1632082664
transform 1 0 9568 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1332_
timestamp 1632082664
transform 1 0 8924 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1632082664
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_91
timestamp 1632082664
transform 1 0 9476 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_101
timestamp 1632082664
transform 1 0 10396 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1330_
timestamp 1632082664
transform 1 0 10764 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1632082664
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1632082664
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1632082664
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1632082664
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1632082664
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1632082664
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1324_
timestamp 1632082664
transform 1 0 13800 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1632082664
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1632082664
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1632082664
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_137
timestamp 1632082664
transform 1 0 13708 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_117_clk
timestamp 1632082664
transform 1 0 15548 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1632082664
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_154
timestamp 1632082664
transform 1 0 15272 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_153
timestamp 1632082664
transform 1 0 15180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1779_
timestamp 1632082664
transform 1 0 16652 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1632082664
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_185
timestamp 1632082664
transform 1 0 18124 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1632082664
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1632082664
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_197
timestamp 1632082664
transform 1 0 19228 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1425_
timestamp 1632082664
transform 1 0 19872 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1632082664
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1632082664
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1632082664
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_203
timestamp 1632082664
transform 1 0 19780 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1424_
timestamp 1632082664
transform 1 0 20700 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_229
timestamp 1632082664
transform 1 0 22172 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1632082664
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1632082664
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_209
timestamp 1632082664
transform 1 0 20332 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1632082664
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_241
timestamp 1632082664
transform 1 0 23276 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_237
timestamp 1632082664
transform 1 0 22908 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1691_
timestamp 1632082664
transform 1 0 23736 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_19_245
timestamp 1632082664
transform 1 0 23644 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1632082664
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_253
timestamp 1632082664
transform 1 0 24380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_261
timestamp 1632082664
transform 1 0 25116 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1689_
timestamp 1632082664
transform 1 0 25300 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_19_262
timestamp 1632082664
transform 1 0 25208 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1632082664
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1632082664
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1455_
timestamp 1632082664
transform 1 0 27232 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1454_
timestamp 1632082664
transform 1 0 27140 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1632082664
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_279
timestamp 1632082664
transform 1 0 26772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_281
timestamp 1632082664
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_299
timestamp 1632082664
transform 1 0 28612 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1457_
timestamp 1632082664
transform 1 0 29072 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1632082664
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1632082664
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1632082664
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_300
timestamp 1632082664
transform 1 0 28704 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1464_
timestamp 1632082664
transform 1 0 30912 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_19_320
timestamp 1632082664
transform 1 0 30544 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_332
timestamp 1632082664
transform 1 0 31648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_321
timestamp 1632082664
transform 1 0 30636 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1468_
timestamp 1632082664
transform 1 0 32752 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1466_
timestamp 1632082664
transform 1 0 32108 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_19_353
timestamp 1632082664
transform 1 0 33580 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1632082664
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_340
timestamp 1632082664
transform 1 0 32384 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1673_
timestamp 1632082664
transform 1 0 34684 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1671_
timestamp 1632082664
transform 1 0 34960 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1632082664
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1632082664
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_365
timestamp 1632082664
transform 1 0 34684 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_381
timestamp 1632082664
transform 1 0 36156 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_384
timestamp 1632082664
transform 1 0 36432 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1632082664
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_393
timestamp 1632082664
transform 1 0 37260 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_389
timestamp 1632082664
transform 1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_412
timestamp 1632082664
transform 1 0 39008 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1625_
timestamp 1632082664
transform 1 0 37536 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1624_
timestamp 1632082664
transform 1 0 37536 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_19_412
timestamp 1632082664
transform 1 0 39008 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1632082664
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_436
timestamp 1632082664
transform 1 0 41216 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_424
timestamp 1632082664
transform 1 0 40112 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1632082664
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_437
timestamp 1632082664
transform 1 0 41308 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_433
timestamp 1632082664
transform 1 0 40940 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_95_clk
timestamp 1632082664
transform 1 0 43148 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_19_449
timestamp 1632082664
transform 1 0 42412 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0088_
timestamp 1632082664
transform 1 0 41400 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_454
timestamp 1632082664
transform 1 0 42872 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1632082664
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_466
timestamp 1632082664
transform 1 0 43976 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_474
timestamp 1632082664
transform 1 0 44712 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0154_
timestamp 1632082664
transform 1 0 44988 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1632082664
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_477
timestamp 1632082664
transform 1 0 44988 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1632082664
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0121_
timestamp 1632082664
transform 1 0 45356 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_493
timestamp 1632082664
transform 1 0 46460 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1589_
timestamp 1632082664
transform 1 0 48668 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1565_
timestamp 1632082664
transform 1 0 47932 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_19_505
timestamp 1632082664
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1632082664
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1632082664
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_505
timestamp 1632082664
transform 1 0 47564 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1632082664
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1588_
timestamp 1632082664
transform 1 0 50508 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1568_
timestamp 1632082664
transform 1 0 50140 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1632082664
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1632082664
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_533
timestamp 1632082664
transform 1 0 50140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1632082664
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_561
timestamp 1632082664
transform 1 0 52716 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1571_
timestamp 1632082664
transform 1 0 51980 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1632082664
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1632082664
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_549
timestamp 1632082664
transform 1 0 51612 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1632082664
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1573_
timestamp 1632082664
transform 1 0 53452 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_569
timestamp 1632082664
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_90_clk
timestamp 1632082664
transform 1 0 56672 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_19_585
timestamp 1632082664
transform 1 0 54924 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1533_
timestamp 1632082664
transform 1 0 55936 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_589
timestamp 1632082664
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1632082664
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1632082664
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_601
timestamp 1632082664
transform 1 0 56396 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_593
timestamp 1632082664
transform 1 0 55660 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_624
timestamp 1632082664
transform 1 0 58512 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_617
timestamp 1632082664
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1632082664
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_612
timestamp 1632082664
transform 1 0 57408 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_629
timestamp 1632082664
transform 1 0 58972 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1632082664
transform -1 0 59340 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1632082664
transform -1 0 59340 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1280_
timestamp 1632082664
transform 1 0 1656 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1632082664
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1632082664
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_34
timestamp 1632082664
transform 1 0 4232 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_22
timestamp 1632082664
transform 1 0 3128 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_46
timestamp 1632082664
transform 1 0 5336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1632082664
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1632082664
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1292_
timestamp 1632082664
transform 1 0 6532 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1632082664
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_75
timestamp 1632082664
transform 1 0 8004 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1329_
timestamp 1632082664
transform 1 0 9568 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_91
timestamp 1632082664
transform 1 0 9476 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_87
timestamp 1632082664
transform 1 0 9108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1328_
timestamp 1632082664
transform 1 0 11500 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1632082664
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1632082664
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1323_
timestamp 1632082664
transform 1 0 14076 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_21_129
timestamp 1632082664
transform 1 0 12972 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_157
timestamp 1632082664
transform 1 0 15548 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1632082664
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1781_
timestamp 1632082664
transform 1 0 16652 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_21_185
timestamp 1632082664
transform 1 0 18124 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1632082664
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_197
timestamp 1632082664
transform 1 0 19228 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1427_
timestamp 1632082664
transform 1 0 19872 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_203
timestamp 1632082664
transform 1 0 19780 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1428_
timestamp 1632082664
transform 1 0 21804 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1632082664
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1632082664
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_241
timestamp 1632082664
transform 1 0 23276 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_253
timestamp 1632082664
transform 1 0 24380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1688_
timestamp 1632082664
transform 1 0 25024 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_259
timestamp 1632082664
transform 1 0 24932 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1453_
timestamp 1632082664
transform 1 0 26956 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1632082664
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1632082664
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1459_
timestamp 1632082664
transform 1 0 28796 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_297
timestamp 1632082664
transform 1 0 28428 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1632082664
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1632082664
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_337
timestamp 1632082664
transform 1 0 32108 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1674_
timestamp 1632082664
transform 1 0 32752 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1632082664
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_343
timestamp 1632082664
transform 1 0 32660 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1632082664
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_360
timestamp 1632082664
transform 1 0 34224 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1670_
timestamp 1632082664
transform 1 0 34960 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_21_384
timestamp 1632082664
transform 1 0 36432 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1632082664
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_393
timestamp 1632082664
transform 1 0 37260 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1626_
timestamp 1632082664
transform 1 0 37536 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_21_412
timestamp 1632082664
transform 1 0 39008 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_436
timestamp 1632082664
transform 1 0 41216 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_424
timestamp 1632082664
transform 1 0 40112 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0099_
timestamp 1632082664
transform 1 0 42872 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1632082664
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_453
timestamp 1632082664
transform 1 0 42780 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_449
timestamp 1632082664
transform 1 0 42412 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0132_
timestamp 1632082664
transform 1 0 44712 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_470
timestamp 1632082664
transform 1 0 44344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_490
timestamp 1632082664
transform 1 0 46184 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_502
timestamp 1632082664
transform 1 0 47288 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1563_
timestamp 1632082664
transform 1 0 47656 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1632082664
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_505
timestamp 1632082664
transform 1 0 47564 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_522
timestamp 1632082664
transform 1 0 49128 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1567_
timestamp 1632082664
transform 1 0 49772 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_528
timestamp 1632082664
transform 1 0 49680 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_545
timestamp 1632082664
transform 1 0 51244 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1632082664
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_561
timestamp 1632082664
transform 1 0 52716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_557
timestamp 1632082664
transform 1 0 52348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_89_clk
timestamp 1632082664
transform 1 0 53084 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_21_585
timestamp 1632082664
transform 1 0 54924 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1537_
timestamp 1632082664
transform 1 0 55936 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_21_593
timestamp 1632082664
transform 1 0 55660 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_617
timestamp 1632082664
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1632082664
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_612
timestamp 1632082664
transform 1 0 57408 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_629
timestamp 1632082664
transform 1 0 58972 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1632082664
transform -1 0 59340 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1279_
timestamp 1632082664
transform 1 0 1656 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1632082664
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1632082664
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_clk
timestamp 1632082664
transform 1 0 4508 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_22_22
timestamp 1632082664
transform 1 0 3128 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_29
timestamp 1632082664
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1632082664
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1293_
timestamp 1632082664
transform 1 0 6716 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_57
timestamp 1632082664
transform 1 0 6348 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1632082664
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1632082664
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_clk
timestamp 1632082664
transform 1 0 9844 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1632082664
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1632082664
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1632082664
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1325_
timestamp 1632082664
transform 1 0 12144 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_119
timestamp 1632082664
transform 1 0 12052 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_115
timestamp 1632082664
transform 1 0 11684 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1322_
timestamp 1632082664
transform 1 0 14076 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1632082664
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1632082664
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_157
timestamp 1632082664
transform 1 0 15548 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1783_
timestamp 1632082664
transform 1 0 17112 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_173
timestamp 1632082664
transform 1 0 17020 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_169
timestamp 1632082664
transform 1 0 16652 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_190
timestamp 1632082664
transform 1 0 18584 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1632082664
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1632082664
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1426_
timestamp 1632082664
transform 1 0 20424 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_209
timestamp 1632082664
transform 1 0 20332 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_226
timestamp 1632082664
transform 1 0 21896 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_246
timestamp 1632082664
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1429_
timestamp 1632082664
transform 1 0 22264 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_111_clk
timestamp 1632082664
transform 1 0 25944 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1632082664
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1632082664
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_269
timestamp 1632082664
transform 1 0 25852 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_265
timestamp 1632082664
transform 1 0 25484 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_290
timestamp 1632082664
transform 1 0 27784 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_302
timestamp 1632082664
transform 1 0 28888 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_309
timestamp 1632082664
transform 1 0 29532 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1632082664
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_317
timestamp 1632082664
transform 1 0 30268 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1678_
timestamp 1632082664
transform 1 0 30452 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_100_clk
timestamp 1632082664
transform 1 0 32292 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_22_335
timestamp 1632082664
transform 1 0 31924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1632082664
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1669_
timestamp 1632082664
transform 1 0 34868 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1632082664
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1632082664
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_359
timestamp 1632082664
transform 1 0 34132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_383
timestamp 1632082664
transform 1 0 36340 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_395
timestamp 1632082664
transform 1 0 37444 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_101_clk
timestamp 1632082664
transform 1 0 37536 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_22_416
timestamp 1632082664
transform 1 0 39376 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1634_
timestamp 1632082664
transform 1 0 39836 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_22_437
timestamp 1632082664
transform 1 0 41308 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1632082664
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_449
timestamp 1632082664
transform 1 0 42412 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_461
timestamp 1632082664
transform 1 0 43516 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1632082664
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_477
timestamp 1632082664
transform 1 0 44988 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_473
timestamp 1632082664
transform 1 0 44620 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_496
timestamp 1632082664
transform 1 0 46736 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0165_
timestamp 1632082664
transform 1 0 45264 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1562_
timestamp 1632082664
transform 1 0 47564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_504
timestamp 1632082664
transform 1 0 47472 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_521
timestamp 1632082664
transform 1 0 49036 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1566_
timestamp 1632082664
transform 1 0 50140 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1632082664
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_529
timestamp 1632082664
transform 1 0 49772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1570_
timestamp 1632082664
transform 1 0 51980 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_549
timestamp 1632082664
transform 1 0 51612 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1632082664
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_569
timestamp 1632082664
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1536_
timestamp 1632082664
transform 1 0 56672 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_22_589
timestamp 1632082664
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1632082664
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1632082664
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_601
timestamp 1632082664
transform 1 0 56396 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_620
timestamp 1632082664
transform 1 0 58144 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_628
timestamp 1632082664
transform 1 0 58880 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1632082664
transform -1 0 59340 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1278_
timestamp 1632082664
transform 1 0 1656 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1632082664
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1632082664
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_34
timestamp 1632082664
transform 1 0 4232 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_22
timestamp 1632082664
transform 1 0 3128 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_46
timestamp 1632082664
transform 1 0 5336 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1632082664
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1632082664
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1294_
timestamp 1632082664
transform 1 0 6532 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1632082664
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1334_
timestamp 1632082664
transform 1 0 8464 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_23_79
timestamp 1632082664
transform 1 0 8372 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_75
timestamp 1632082664
transform 1 0 8004 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_96
timestamp 1632082664
transform 1 0 9936 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1632082664
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1327_
timestamp 1632082664
transform 1 0 12236 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1632082664
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1632082664
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_137
timestamp 1632082664
transform 1 0 13708 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1321_
timestamp 1632082664
transform 1 0 14260 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_23_159
timestamp 1632082664
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1632082664
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1784_
timestamp 1632082664
transform 1 0 17388 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1632082664
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1632082664
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1787_
timestamp 1632082664
transform 1 0 19228 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_193
timestamp 1632082664
transform 1 0 18860 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_213
timestamp 1632082664
transform 1 0 20700 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1632082664
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1632082664
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 1632082664
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_237
timestamp 1632082664
transform 1 0 22908 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1690_
timestamp 1632082664
transform 1 0 23092 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1449_
timestamp 1632082664
transform 1 0 24932 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_255
timestamp 1632082664
transform 1 0 24564 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1452_
timestamp 1632082664
transform 1 0 26956 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1632082664
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1632082664
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_275
timestamp 1632082664
transform 1 0 26404 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1687_
timestamp 1632082664
transform 1 0 28796 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_297
timestamp 1632082664
transform 1 0 28428 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1632082664
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1632082664
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_337
timestamp 1632082664
transform 1 0 32108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1672_
timestamp 1632082664
transform 1 0 32844 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1632082664
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1632082664
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1668_
timestamp 1632082664
transform 1 0 34684 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_361
timestamp 1632082664
transform 1 0 34316 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_381
timestamp 1632082664
transform 1 0 36156 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1632082664
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_393
timestamp 1632082664
transform 1 0 37260 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_389
timestamp 1632082664
transform 1 0 36892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1627_
timestamp 1632082664
transform 1 0 37536 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_23_416
timestamp 1632082664
transform 1 0 39376 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_412
timestamp 1632082664
transform 1 0 39008 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1630_
timestamp 1632082664
transform 1 0 39468 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_23_433
timestamp 1632082664
transform 1 0 40940 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1632082664
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1632082664
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_445
timestamp 1632082664
transform 1 0 42044 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0176_
timestamp 1632082664
transform 1 0 44988 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1632082664
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_473
timestamp 1632082664
transform 1 0 44620 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_493
timestamp 1632082664
transform 1 0 46460 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1561_
timestamp 1632082664
transform 1 0 47656 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1632082664
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_505
timestamp 1632082664
transform 1 0 47564 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_501
timestamp 1632082664
transform 1 0 47196 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1564_
timestamp 1632082664
transform 1 0 49496 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_522
timestamp 1632082664
transform 1 0 49128 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_554
timestamp 1632082664
transform 1 0 52072 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1574_
timestamp 1632082664
transform 1 0 52716 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_23_542
timestamp 1632082664
transform 1 0 50968 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1632082664
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_577
timestamp 1632082664
transform 1 0 54188 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_589
timestamp 1632082664
transform 1 0 55292 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1538_
timestamp 1632082664
transform 1 0 55936 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_23_595
timestamp 1632082664
transform 1 0 55844 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_617
timestamp 1632082664
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1632082664
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_612
timestamp 1632082664
transform 1 0 57408 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_629
timestamp 1632082664
transform 1 0 58972 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1632082664
transform -1 0 59340 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1277_
timestamp 1632082664
transform 1 0 1840 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1632082664
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1632082664
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1632082664
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_41
timestamp 1632082664
transform 1 0 4876 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1632082664
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1632082664
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1632082664
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1295_
timestamp 1632082664
transform 1 0 5520 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_24_47
timestamp 1632082664
transform 1 0 5428 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_76
timestamp 1632082664
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_64
timestamp 1632082664
transform 1 0 6992 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1331_
timestamp 1632082664
transform 1 0 10396 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1632082664
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1632082664
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_97
timestamp 1632082664
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1632082664
transform 1 0 11868 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_129
timestamp 1632082664
transform 1 0 12972 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1320_
timestamp 1632082664
transform 1 0 14352 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1632082664
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_141
timestamp 1632082664
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_137
timestamp 1632082664
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_160
timestamp 1632082664
transform 1 0 15824 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1785_
timestamp 1632082664
transform 1 0 17296 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_172
timestamp 1632082664
transform 1 0 16928 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_110_clk
timestamp 1632082664
transform 1 0 19872 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_24_197
timestamp 1632082664
transform 1 0 19228 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1632082664
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_203
timestamp 1632082664
transform 1 0 19780 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1632082664
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1430_
timestamp 1632082664
transform 1 0 22080 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_224
timestamp 1632082664
transform 1 0 21712 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_244
timestamp 1632082664
transform 1 0 23552 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_269
timestamp 1632082664
transform 1 0 25852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1447_
timestamp 1632082664
transform 1 0 24380 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1632082664
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_277
timestamp 1632082664
transform 1 0 26588 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1451_
timestamp 1632082664
transform 1 0 26772 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1632082664
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_295
timestamp 1632082664
transform 1 0 28244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1632082664
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1632082664
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1677_
timestamp 1632082664
transform 1 0 30728 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_24_321
timestamp 1632082664
transform 1 0 30636 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_338
timestamp 1632082664
transform 1 0 32200 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1675_
timestamp 1632082664
transform 1 0 32752 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1667_
timestamp 1632082664
transform 1 0 34684 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1632082664
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_360
timestamp 1632082664
transform 1 0 34224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_381
timestamp 1632082664
transform 1 0 36156 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_393
timestamp 1632082664
transform 1 0 37260 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1632082664
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1628_
timestamp 1632082664
transform 1 0 37628 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1632_
timestamp 1632082664
transform 1 0 39836 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1632082664
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1632082664
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_437
timestamp 1632082664
transform 1 0 41308 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1635_
timestamp 1632082664
transform 1 0 41676 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1632082664
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1632082664
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0187_
timestamp 1632082664
transform 1 0 44988 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1632082664
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1632082664
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_493
timestamp 1632082664
transform 1 0 46460 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_88_clk
timestamp 1632082664
transform 1 0 47840 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_24_505
timestamp 1632082664
transform 1 0 47564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1569_
timestamp 1632082664
transform 1 0 50140 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1632082664
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_528
timestamp 1632082664
transform 1 0 49680 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1572_
timestamp 1632082664
transform 1 0 51980 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_549
timestamp 1632082664
transform 1 0 51612 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1632082664
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_569
timestamp 1632082664
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1539_
timestamp 1632082664
transform 1 0 56396 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_24_589
timestamp 1632082664
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1632082664
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1632082664
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_617
timestamp 1632082664
transform 1 0 57868 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_629
timestamp 1632082664
transform 1 0 58972 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1632082664
transform -1 0 59340 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1276_
timestamp 1632082664
transform 1 0 1472 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1632082664
transform 1 0 1380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_20
timestamp 1632082664
transform 1 0 2944 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1632082664
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1275_
timestamp 1632082664
transform 1 0 3312 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_25_40
timestamp 1632082664
transform 1 0 4784 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1296_
timestamp 1632082664
transform 1 0 6348 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1632082664
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1632082664
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1300_
timestamp 1632082664
transform 1 0 8188 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_73
timestamp 1632082664
transform 1 0 7820 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1632082664
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1632082664
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1632082664
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1632082664
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1632082664
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1632082664
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_137
timestamp 1632082664
transform 1 0 13708 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1319_
timestamp 1632082664
transform 1 0 14352 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_25_143
timestamp 1632082664
transform 1 0 14260 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_160
timestamp 1632082664
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp 1632082664
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1786_
timestamp 1632082664
transform 1 0 17296 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1632082664
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_175
timestamp 1632082664
transform 1 0 17204 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1791_
timestamp 1632082664
transform 1 0 19136 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_192
timestamp 1632082664
transform 1 0 18768 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1432_
timestamp 1632082664
transform 1 0 21804 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_25_212
timestamp 1632082664
transform 1 0 20608 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1632082664
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_241
timestamp 1632082664
transform 1 0 23276 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_269
timestamp 1632082664
transform 1 0 25852 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1446_
timestamp 1632082664
transform 1 0 24380 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1450_
timestamp 1632082664
transform 1 0 26956 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1632082664
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_277
timestamp 1632082664
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_309
timestamp 1632082664
transform 1 0 29532 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_297
timestamp 1632082664
transform 1 0 28428 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1680_
timestamp 1632082664
transform 1 0 30176 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_25_315
timestamp 1632082664
transform 1 0 30084 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_332
timestamp 1632082664
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1683_
timestamp 1632082664
transform 1 0 32108 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_25_353
timestamp 1632082664
transform 1 0 33580 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1632082664
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1666_
timestamp 1632082664
transform 1 0 34684 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_25_393
timestamp 1632082664
transform 1 0 37260 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_381
timestamp 1632082664
transform 1 0 36156 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1632082664
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_389
timestamp 1632082664
transform 1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_415
timestamp 1632082664
transform 1 0 39284 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1629_
timestamp 1632082664
transform 1 0 37812 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1633_
timestamp 1632082664
transform 1 0 40112 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_25_423
timestamp 1632082664
transform 1 0 40020 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_440
timestamp 1632082664
transform 1 0 41584 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1637_
timestamp 1632082664
transform 1 0 42412 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1632082664
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0198_
timestamp 1632082664
transform 1 0 44988 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_25_465
timestamp 1632082664
transform 1 0 43884 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_493
timestamp 1632082664
transform 1 0 46460 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1560_
timestamp 1632082664
transform 1 0 47656 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1632082664
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_505
timestamp 1632082664
transform 1 0 47564 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_501
timestamp 1632082664
transform 1 0 47196 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1556_
timestamp 1632082664
transform 1 0 50324 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_25_522
timestamp 1632082664
transform 1 0 49128 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_534
timestamp 1632082664
transform 1 0 50232 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_551
timestamp 1632082664
transform 1 0 51796 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_561
timestamp 1632082664
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1632082664
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1632082664
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1547_
timestamp 1632082664
transform 1 0 54096 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_25_573
timestamp 1632082664
transform 1 0 53820 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1541_
timestamp 1632082664
transform 1 0 55936 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_592
timestamp 1632082664
transform 1 0 55568 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_617
timestamp 1632082664
transform 1 0 57868 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1632082664
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_612
timestamp 1632082664
transform 1 0 57408 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_629
timestamp 1632082664
transform 1 0 58972 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1632082664
transform -1 0 59340 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1271_
timestamp 1632082664
transform 1 0 2484 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1632082664
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1632082664
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1632082664
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1632082664
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1632082664
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1274_
timestamp 1632082664
transform 1 0 4324 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1273_
timestamp 1632082664
transform 1 0 3772 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1632082664
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1632082664
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_31
timestamp 1632082664
transform 1 0 3956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1298_
timestamp 1632082664
transform 1 0 6348 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1297_
timestamp 1632082664
transform 1 0 5612 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1632082664
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1632082664
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1632082664
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_45
timestamp 1632082664
transform 1 0 5244 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1632082664
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1301_
timestamp 1632082664
transform 1 0 8188 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1632082664
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1632082664
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_73
timestamp 1632082664
transform 1 0 7820 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1303_
timestamp 1632082664
transform 1 0 8924 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1632082664
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1632082664
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_101
timestamp 1632082664
transform 1 0 10396 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1632082664
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1307_
timestamp 1632082664
transform 1 0 11500 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1306_
timestamp 1632082664
transform 1 0 10764 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1632082664
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1632082664
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1632082664
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1632082664
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1317_
timestamp 1632082664
transform 1 0 14076 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1316_
timestamp 1632082664
transform 1 0 14076 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_27_129
timestamp 1632082664
transform 1 0 12972 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1632082664
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1632082664
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_157
timestamp 1632082664
transform 1 0 15548 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_157
timestamp 1632082664
transform 1 0 15548 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1632082664
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_169
timestamp 1632082664
transform 1 0 16652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1790_
timestamp 1632082664
transform 1 0 17204 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1788_
timestamp 1632082664
transform 1 0 17112 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1632082664
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_173
timestamp 1632082664
transform 1 0 17020 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_169
timestamp 1632082664
transform 1 0 16652 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_190
timestamp 1632082664
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1436_
timestamp 1632082664
transform 1 0 19872 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_27_191
timestamp 1632082664
transform 1 0 18676 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1632082664
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1632082664
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_203
timestamp 1632082664
transform 1 0 19780 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_209
timestamp 1632082664
transform 1 0 20332 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1433_
timestamp 1632082664
transform 1 0 21804 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1431_
timestamp 1632082664
transform 1 0 20884 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1632082664
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1632082664
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_243
timestamp 1632082664
transform 1 0 23460 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_241
timestamp 1632082664
transform 1 0 23276 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_231
timestamp 1632082664
transform 1 0 22356 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_269
timestamp 1632082664
transform 1 0 25852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1445_
timestamp 1632082664
transform 1 0 24380 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1444_
timestamp 1632082664
transform 1 0 24380 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1632082664
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1632082664
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_269
timestamp 1632082664
transform 1 0 25852 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1448_
timestamp 1632082664
transform 1 0 26220 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1632082664
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1632082664
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1632082664
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1632082664
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1632082664
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1684_
timestamp 1632082664
transform 1 0 28336 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1632082664
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1632082664
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1632082664
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_312
timestamp 1632082664
transform 1 0 29808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_293
timestamp 1632082664
transform 1 0 28060 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1682_
timestamp 1632082664
transform 1 0 30176 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1679_
timestamp 1632082664
transform 1 0 31004 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1632082664
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_321
timestamp 1632082664
transform 1 0 30636 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_353
timestamp 1632082664
transform 1 0 33580 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1686_
timestamp 1632082664
transform 1 0 32108 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_26_341
timestamp 1632082664
transform 1 0 32476 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1632082664
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_353
timestamp 1632082664
transform 1 0 33580 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1664_
timestamp 1632082664
transform 1 0 33948 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1632082664
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1632082664
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1632082664
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_361
timestamp 1632082664
transform 1 0 34316 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1632082664
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1663_
timestamp 1632082664
transform 1 0 36064 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1657_
timestamp 1632082664
transform 1 0 37352 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1632082664
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_393
timestamp 1632082664
transform 1 0 37260 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1632082664
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_377
timestamp 1632082664
transform 1 0 35788 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1997_
timestamp 1632082664
transform 1 0 39192 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1631_
timestamp 1632082664
transform 1 0 37904 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_27_410
timestamp 1632082664
transform 1 0 38824 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_416
timestamp 1632082664
transform 1 0 39376 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_396
timestamp 1632082664
transform 1 0 37536 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_421
timestamp 1632082664
transform 1 0 39836 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1636_
timestamp 1632082664
transform 1 0 40664 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_27_430
timestamp 1632082664
transform 1 0 40664 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1632082664
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_429
timestamp 1632082664
transform 1 0 40572 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_442
timestamp 1632082664
transform 1 0 41768 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1639_
timestamp 1632082664
transform 1 0 42412 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1638_
timestamp 1632082664
transform 1 0 42504 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1632082664
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_446
timestamp 1632082664
transform 1 0 42136 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_466
timestamp 1632082664
transform 1 0 43976 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_474
timestamp 1632082664
transform 1 0 44712 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0220_
timestamp 1632082664
transform 1 0 44988 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0209_
timestamp 1632082664
transform 1 0 44988 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_27_465
timestamp 1632082664
transform 1 0 43884 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1632082664
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_493
timestamp 1632082664
transform 1 0 46460 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_493
timestamp 1632082664
transform 1 0 46460 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_501
timestamp 1632082664
transform 1 0 47196 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1558_
timestamp 1632082664
transform 1 0 47380 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1557_
timestamp 1632082664
transform 1 0 48944 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_27_505
timestamp 1632082664
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_519
timestamp 1632082664
transform 1 0 48852 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1632082664
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_517
timestamp 1632082664
transform 1 0 48668 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_501
timestamp 1632082664
transform 1 0 47196 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1554_
timestamp 1632082664
transform 1 0 50784 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_26_533
timestamp 1632082664
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1632082664
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1632082664
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_536
timestamp 1632082664
transform 1 0 50416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1553_
timestamp 1632082664
transform 1 0 51520 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_27_561
timestamp 1632082664
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1632082664
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_556
timestamp 1632082664
transform 1 0 52256 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_545
timestamp 1632082664
transform 1 0 51244 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1548_
timestamp 1632082664
transform 1 0 53360 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1546_
timestamp 1632082664
transform 1 0 54096 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_26_564
timestamp 1632082664
transform 1 0 52992 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_573
timestamp 1632082664
transform 1 0 53820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1543_
timestamp 1632082664
transform 1 0 55936 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1540_
timestamp 1632082664
transform 1 0 56488 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_26_589
timestamp 1632082664
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1632082664
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_601
timestamp 1632082664
transform 1 0 56396 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_592
timestamp 1632082664
transform 1 0 55568 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_584
timestamp 1632082664
transform 1 0 54832 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_617
timestamp 1632082664
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_618
timestamp 1632082664
transform 1 0 57960 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1632082664
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_612
timestamp 1632082664
transform 1 0 57408 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_629
timestamp 1632082664
transform 1 0 58972 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1632082664
transform -1 0 59340 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1632082664
transform -1 0 59340 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1632082664
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1632082664
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1632082664
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1272_
timestamp 1632082664
transform 1 0 3772 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1632082664
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1632082664
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_45
timestamp 1632082664
transform 1 0 5244 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1299_
timestamp 1632082664
transform 1 0 6256 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_28_53
timestamp 1632082664
transform 1 0 5980 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_72
timestamp 1632082664
transform 1 0 7728 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1304_
timestamp 1632082664
transform 1 0 8924 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1632082664
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_101
timestamp 1632082664
transform 1 0 10396 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1305_
timestamp 1632082664
transform 1 0 10764 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1632082664
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1632082664
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1315_
timestamp 1632082664
transform 1 0 14076 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1632082664
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1632082664
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1318_
timestamp 1632082664
transform 1 0 15916 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_28_157
timestamp 1632082664
transform 1 0 15548 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1632082664
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1632082664
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1632082664
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1632082664
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1632082664
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_209
timestamp 1632082664
transform 1 0 20332 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1434_
timestamp 1632082664
transform 1 0 20884 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_28_243
timestamp 1632082664
transform 1 0 23460 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_231
timestamp 1632082664
transform 1 0 22356 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_253
timestamp 1632082664
transform 1 0 24380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1443_
timestamp 1632082664
transform 1 0 25116 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1632082664
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1632082664
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_277
timestamp 1632082664
transform 1 0 26588 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1685_
timestamp 1632082664
transform 1 0 27600 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_28_285
timestamp 1632082664
transform 1 0 27324 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1632082664
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1632082664
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1632082664
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1681_
timestamp 1632082664
transform 1 0 30912 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_28_321
timestamp 1632082664
transform 1 0 30636 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1665_
timestamp 1632082664
transform 1 0 32752 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_28_340
timestamp 1632082664
transform 1 0 32384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1632082664
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1632082664
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_360
timestamp 1632082664
transform 1 0 34224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1659_
timestamp 1632082664
transform 1 0 36064 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_28_377
timestamp 1632082664
transform 1 0 35788 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1654_
timestamp 1632082664
transform 1 0 37904 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_28_416
timestamp 1632082664
transform 1 0 39376 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_396
timestamp 1632082664
transform 1 0 37536 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1632082664
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1632082664
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1632082664
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1640_
timestamp 1632082664
transform 1 0 42136 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_28_445
timestamp 1632082664
transform 1 0 42044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_474
timestamp 1632082664
transform 1 0 44712 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0231_
timestamp 1632082664
transform 1 0 44988 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_28_462
timestamp 1632082664
transform 1 0 43608 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1632082664
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_493
timestamp 1632082664
transform 1 0 46460 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1559_
timestamp 1632082664
transform 1 0 47656 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_28_505
timestamp 1632082664
transform 1 0 47564 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_522
timestamp 1632082664
transform 1 0 49128 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_530
timestamp 1632082664
transform 1 0 49864 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_533
timestamp 1632082664
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1632082664
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1551_
timestamp 1632082664
transform 1 0 51244 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_28_561
timestamp 1632082664
transform 1 0 52716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1632082664
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1550_
timestamp 1632082664
transform 1 0 53084 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_28_589
timestamp 1632082664
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1632082664
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1632082664
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_601
timestamp 1632082664
transform 1 0 56396 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_621
timestamp 1632082664
transform 1 0 58236 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1542_
timestamp 1632082664
transform 1 0 56764 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_28_629
timestamp 1632082664
transform 1 0 58972 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1632082664
transform -1 0 59340 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1269_
timestamp 1632082664
transform 1 0 1748 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1632082664
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1632082664
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1270_
timestamp 1632082664
transform 1 0 3588 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_23
timestamp 1632082664
transform 1 0 3220 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1260_
timestamp 1632082664
transform 1 0 6348 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_29_43
timestamp 1632082664
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1632082664
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1632082664
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1302_
timestamp 1632082664
transform 1 0 8188 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_73
timestamp 1632082664
transform 1 0 7820 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1632082664
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1632082664
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1308_
timestamp 1632082664
transform 1 0 11500 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1632082664
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1632082664
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1312_
timestamp 1632082664
transform 1 0 13340 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_129
timestamp 1632082664
transform 1 0 12972 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1632082664
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1632082664
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1792_
timestamp 1632082664
transform 1 0 18032 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1632082664
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1632082664
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1632082664
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_181
timestamp 1632082664
transform 1 0 17756 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1437_
timestamp 1632082664
transform 1 0 19872 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_200
timestamp 1632082664
transform 1 0 19504 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1440_
timestamp 1632082664
transform 1 0 21804 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1632082664
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1632082664
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1442_
timestamp 1632082664
transform 1 0 23644 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_241
timestamp 1632082664
transform 1 0 23276 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_261
timestamp 1632082664
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_281
timestamp 1632082664
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1632082664
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0946_
timestamp 1632082664
transform 1 0 27508 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1632082664
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1632082664
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_303
timestamp 1632082664
transform 1 0 28980 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0902_
timestamp 1632082664
transform 1 0 29808 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_29_311
timestamp 1632082664
transform 1 0 29716 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_328
timestamp 1632082664
transform 1 0 31280 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1662_
timestamp 1632082664
transform 1 0 33488 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1632082664
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1632082664
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_349
timestamp 1632082664
transform 1 0 33212 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1660_
timestamp 1632082664
transform 1 0 35328 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_368
timestamp 1632082664
transform 1 0 34960 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_393
timestamp 1632082664
transform 1 0 37260 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1632082664
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_388
timestamp 1632082664
transform 1 0 36800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1652_
timestamp 1632082664
transform 1 0 38272 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_29_401
timestamp 1632082664
transform 1 0 37996 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_102_clk
timestamp 1632082664
transform 1 0 40112 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_29_420
timestamp 1632082664
transform 1 0 39744 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1641_
timestamp 1632082664
transform 1 0 42412 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1632082664
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_444
timestamp 1632082664
transform 1 0 41952 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0242_
timestamp 1632082664
transform 1 0 44988 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_29_465
timestamp 1632082664
transform 1 0 43884 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_493
timestamp 1632082664
transform 1 0 46460 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_517
timestamp 1632082664
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_505
timestamp 1632082664
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1632082664
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_501
timestamp 1632082664
transform 1 0 47196 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_529
timestamp 1632082664
transform 1 0 49772 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_537
timestamp 1632082664
transform 1 0 50508 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1555_
timestamp 1632082664
transform 1 0 50692 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_29_561
timestamp 1632082664
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1632082664
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1632082664
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_555
timestamp 1632082664
transform 1 0 52164 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1549_
timestamp 1632082664
transform 1 0 53912 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_29_573
timestamp 1632082664
transform 1 0 53820 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_590
timestamp 1632082664
transform 1 0 55384 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1545_
timestamp 1632082664
transform 1 0 55936 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_29_617
timestamp 1632082664
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1632082664
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_612
timestamp 1632082664
transform 1 0 57408 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_629
timestamp 1632082664
transform 1 0 58972 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1632082664
transform -1 0 59340 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1632082664
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1268_
timestamp 1632082664
transform 1 0 1564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1632082664
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1632082664
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1632082664
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1632082664
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1632082664
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1632082664
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1259_
timestamp 1632082664
transform 1 0 6348 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_30_53
timestamp 1632082664
transform 1 0 5980 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_73
timestamp 1632082664
transform 1 0 7820 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_81
timestamp 1632082664
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1265_
timestamp 1632082664
transform 1 0 8924 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_30_101
timestamp 1632082664
transform 1 0 10396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1632082664
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_clk
timestamp 1632082664
transform 1 0 11500 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1632082664
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1313_
timestamp 1632082664
transform 1 0 14076 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1632082664
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1632082664
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1314_
timestamp 1632082664
transform 1 0 15916 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_30_157
timestamp 1632082664
transform 1 0 15548 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1632082664
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1632082664
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1632082664
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1632082664
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1632082664
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1435_
timestamp 1632082664
transform 1 0 20700 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_30_229
timestamp 1632082664
transform 1 0 22172 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_209
timestamp 1632082664
transform 1 0 20332 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_241
timestamp 1632082664
transform 1 0 23276 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1632082664
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_108_clk
timestamp 1632082664
transform 1 0 25668 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_30_265
timestamp 1632082664
transform 1 0 25484 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1632082664
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1632082664
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_287
timestamp 1632082664
transform 1 0 27508 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_299
timestamp 1632082664
transform 1 0 28612 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1632082664
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1632082664
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1632082664
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0869_
timestamp 1632082664
transform 1 0 31096 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_30_325
timestamp 1632082664
transform 1 0 31004 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_321
timestamp 1632082664
transform 1 0 30636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_354
timestamp 1632082664
transform 1 0 33672 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_342
timestamp 1632082664
transform 1 0 32568 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 1632082664
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1632082664
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1632082664
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1656_
timestamp 1632082664
transform 1 0 36064 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_30_377
timestamp 1632082664
transform 1 0 35788 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1653_
timestamp 1632082664
transform 1 0 37904 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_30_416
timestamp 1632082664
transform 1 0 39376 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_396
timestamp 1632082664
transform 1 0 37536 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_437
timestamp 1632082664
transform 1 0 41308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1650_
timestamp 1632082664
transform 1 0 39836 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1632082664
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1642_
timestamp 1632082664
transform 1 0 42320 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_30_445
timestamp 1632082664
transform 1 0 42044 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0253_
timestamp 1632082664
transform 1 0 45080 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_30_464
timestamp 1632082664
transform 1 0 43792 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1632082664
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_477
timestamp 1632082664
transform 1 0 44988 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_494
timestamp 1632082664
transform 1 0 46552 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_518
timestamp 1632082664
transform 1 0 48760 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_506
timestamp 1632082664
transform 1 0 47656 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_530
timestamp 1632082664
transform 1 0 49864 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_533
timestamp 1632082664
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1632082664
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_545
timestamp 1632082664
transform 1 0 51244 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1552_
timestamp 1632082664
transform 1 0 51888 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_30_551
timestamp 1632082664
transform 1 0 51796 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_580
timestamp 1632082664
transform 1 0 54464 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_568
timestamp 1632082664
transform 1 0 53360 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1544_
timestamp 1632082664
transform 1 0 56672 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_30_589
timestamp 1632082664
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1632082664
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_601
timestamp 1632082664
transform 1 0 56396 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_620
timestamp 1632082664
transform 1 0 58144 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_628
timestamp 1632082664
transform 1 0 58880 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1632082664
transform -1 0 59340 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1632082664
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1267_
timestamp 1632082664
transform 1 0 1564 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1632082664
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_21
timestamp 1632082664
transform 1 0 3036 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1255_
timestamp 1632082664
transform 1 0 4048 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_31_29
timestamp 1632082664
transform 1 0 3772 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_48
timestamp 1632082664
transform 1 0 5520 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1258_
timestamp 1632082664
transform 1 0 6348 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1632082664
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1263_
timestamp 1632082664
transform 1 0 8188 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_73
timestamp 1632082664
transform 1 0 7820 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1632082664
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1632082664
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1309_
timestamp 1632082664
transform 1 0 11500 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1632082664
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1632082664
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1311_
timestamp 1632082664
transform 1 0 13340 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_129
timestamp 1632082664
transform 1 0 12972 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1632082664
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_149
timestamp 1632082664
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_169
timestamp 1632082664
transform 1 0 16652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1793_
timestamp 1632082664
transform 1 0 17296 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1632082664
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_175
timestamp 1632082664
transform 1 0 17204 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1632082664
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1438_
timestamp 1632082664
transform 1 0 19872 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_31_192
timestamp 1632082664
transform 1 0 18768 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1439_
timestamp 1632082664
transform 1 0 21804 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1632082664
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1632082664
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1441_
timestamp 1632082664
transform 1 0 23644 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_241
timestamp 1632082664
transform 1 0 23276 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_261
timestamp 1632082664
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1632082664
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0913_
timestamp 1632082664
transform 1 0 26956 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1632082664
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1632082664
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_309
timestamp 1632082664
transform 1 0 29532 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_297
timestamp 1632082664
transform 1 0 28428 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0880_
timestamp 1632082664
transform 1 0 30176 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_31_315
timestamp 1632082664
transform 1 0 30084 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1632082664
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0891_
timestamp 1632082664
transform 1 0 32108 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_31_353
timestamp 1632082664
transform 1 0 33580 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1632082664
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1661_
timestamp 1632082664
transform 1 0 35144 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_31_369
timestamp 1632082664
transform 1 0 35052 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_365
timestamp 1632082664
transform 1 0 34684 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_386
timestamp 1632082664
transform 1 0 36616 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1632082664
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1632082664
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1651_
timestamp 1632082664
transform 1 0 38640 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_31_405
timestamp 1632082664
transform 1 0 38364 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1648_
timestamp 1632082664
transform 1 0 40480 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_424
timestamp 1632082664
transform 1 0 40112 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1643_
timestamp 1632082664
transform 1 0 42412 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1632082664
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_444
timestamp 1632082664
transform 1 0 41952 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_477
timestamp 1632082664
transform 1 0 44988 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0264_
timestamp 1632082664
transform 1 0 45172 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_31_465
timestamp 1632082664
transform 1 0 43884 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_495
timestamp 1632082664
transform 1 0 46644 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0330_
timestamp 1632082664
transform 1 0 47564 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1632082664
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1632082664
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0363_
timestamp 1632082664
transform 1 0 49404 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_31_541
timestamp 1632082664
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_521
timestamp 1632082664
transform 1 0 49036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1632082664
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_561
timestamp 1632082664
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1632082664
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1632082664
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_86_clk
timestamp 1632082664
transform 1 0 54004 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_31_573
timestamp 1632082664
transform 1 0 53820 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_595
timestamp 1632082664
transform 1 0 55844 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_607
timestamp 1632082664
transform 1 0 56948 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_617
timestamp 1632082664
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1632082664
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1632082664
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_629
timestamp 1632082664
transform 1 0 58972 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1632082664
transform -1 0 59340 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1632082664
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1632082664
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1632082664
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp 1632082664
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1254_
timestamp 1632082664
transform 1 0 4324 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1632082664
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1632082664
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_clk
timestamp 1632082664
transform 1 0 6624 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_32_51
timestamp 1632082664
transform 1 0 5796 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_59
timestamp 1632082664
transform 1 0 6532 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1632082664
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1264_
timestamp 1632082664
transform 1 0 8924 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_32_101
timestamp 1632082664
transform 1 0 10396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1632082664
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1310_
timestamp 1632082664
transform 1 0 11500 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_32_141
timestamp 1632082664
transform 1 0 14076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_129
timestamp 1632082664
transform 1 0 12972 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1632082664
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_137
timestamp 1632082664
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_166
timestamp 1632082664
transform 1 0 16376 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1205_
timestamp 1632082664
transform 1 0 14904 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_32_149
timestamp 1632082664
transform 1 0 14812 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_174
timestamp 1632082664
transform 1 0 17112 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1794_
timestamp 1632082664
transform 1 0 17296 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1796_
timestamp 1632082664
transform 1 0 19228 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1632082664
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1632082664
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_109_clk
timestamp 1632082664
transform 1 0 21436 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_32_213
timestamp 1632082664
transform 1 0 20700 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_241
timestamp 1632082664
transform 1 0 23276 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_249
timestamp 1632082664
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1632082664
transform 1 0 24380 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_32_269
timestamp 1632082664
transform 1 0 25852 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1632082664
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_281
timestamp 1632082664
transform 1 0 26956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0924_
timestamp 1632082664
transform 1 0 27140 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_32_299
timestamp 1632082664
transform 1 0 28612 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1632082664
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1632082664
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1632082664
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0836_
timestamp 1632082664
transform 1 0 30728 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_32_321
timestamp 1632082664
transform 1 0 30636 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0858_
timestamp 1632082664
transform 1 0 32568 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_32_338
timestamp 1632082664
transform 1 0 32200 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_358
timestamp 1632082664
transform 1 0 34040 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1632082664
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0726_
timestamp 1632082664
transform 1 0 34868 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1632082664
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_383
timestamp 1632082664
transform 1 0 36340 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_395
timestamp 1632082664
transform 1 0 37444 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1655_
timestamp 1632082664
transform 1 0 37812 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_32_415
timestamp 1632082664
transform 1 0 39284 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_421
timestamp 1632082664
transform 1 0 39836 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1647_
timestamp 1632082664
transform 1 0 40480 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1632082664
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_427
timestamp 1632082664
transform 1 0 40388 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1632082664
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1644_
timestamp 1632082664
transform 1 0 42320 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_32_444
timestamp 1632082664
transform 1 0 41952 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_477
timestamp 1632082664
transform 1 0 44988 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0275_
timestamp 1632082664
transform 1 0 45172 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_32_464
timestamp 1632082664
transform 1 0 43792 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1632082664
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_495
timestamp 1632082664
transform 1 0 46644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0308_
timestamp 1632082664
transform 1 0 47196 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_32_517
timestamp 1632082664
transform 1 0 48668 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0352_
timestamp 1632082664
transform 1 0 50140 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1632082664
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_529
timestamp 1632082664
transform 1 0 49772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1911_
timestamp 1632082664
transform 1 0 51980 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_32_549
timestamp 1632082664
transform 1 0 51612 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1632082664
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_569
timestamp 1632082664
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1915_
timestamp 1632082664
transform 1 0 55292 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1632082664
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1632082664
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1918_
timestamp 1632082664
transform 1 0 57132 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_32_625
timestamp 1632082664
transform 1 0 58604 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_605
timestamp 1632082664
transform 1 0 56764 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_629
timestamp 1632082664
transform 1 0 58972 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1632082664
transform -1 0 59340 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1252_
timestamp 1632082664
transform 1 0 2484 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1632082664
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1632082664
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1632082664
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1632082664
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1632082664
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_clk
timestamp 1632082664
transform 1 0 4140 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1253_
timestamp 1632082664
transform 1 0 4324 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1632082664
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1632082664
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_29
timestamp 1632082664
transform 1 0 3772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_31
timestamp 1632082664
transform 1 0 3956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1257_
timestamp 1632082664
transform 1 0 6348 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1256_
timestamp 1632082664
transform 1 0 6348 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1632082664
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1632082664
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_53
timestamp 1632082664
transform 1 0 5980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1632082664
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_73
timestamp 1632082664
transform 1 0 7820 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1261_
timestamp 1632082664
transform 1 0 8188 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_33_73
timestamp 1632082664
transform 1 0 7820 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_81
timestamp 1632082664
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1266_
timestamp 1632082664
transform 1 0 8924 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_34_101
timestamp 1632082664
transform 1 0 10396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1632082664
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1632082664
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1632082664
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1209_
timestamp 1632082664
transform 1 0 11592 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1207_
timestamp 1632082664
transform 1 0 11868 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1632082664
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_113
timestamp 1632082664
transform 1 0 11500 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1632082664
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_113
timestamp 1632082664
transform 1 0 11500 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1632082664
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_142
timestamp 1632082664
transform 1 0 14168 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_141
timestamp 1632082664
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_130
timestamp 1632082664
transform 1 0 13064 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1632082664
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1632082664
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1204_
timestamp 1632082664
transform 1 0 14720 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1201_
timestamp 1632082664
transform 1 0 15088 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1632082664
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_149
timestamp 1632082664
transform 1 0 14812 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_clk
timestamp 1632082664
transform 1 0 16928 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_33_169
timestamp 1632082664
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1795_
timestamp 1632082664
transform 1 0 17664 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1632082664
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_168
timestamp 1632082664
transform 1 0 16560 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_177
timestamp 1632082664
transform 1 0 17388 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1799_
timestamp 1632082664
transform 1 0 19228 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1797_
timestamp 1632082664
transform 1 0 19504 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1632082664
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1632082664
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_196
timestamp 1632082664
transform 1 0 19136 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_216
timestamp 1632082664
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1804_
timestamp 1632082664
transform 1 0 21804 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1803_
timestamp 1632082664
transform 1 0 21068 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1632082664
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_213
timestamp 1632082664
transform 1 0 20700 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1632082664
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_233
timestamp 1632082664
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_241
timestamp 1632082664
transform 1 0 23276 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_270
timestamp 1632082664
transform 1 0 25944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 1632082664
transform 1 0 24380 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1632082664
transform 1 0 24472 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_34_269
timestamp 1632082664
transform 1 0 25852 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1632082664
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1632082664
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_253
timestamp 1632082664
transform 1 0 24380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1632082664
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0957_
timestamp 1632082664
transform 1 0 27416 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0935_
timestamp 1632082664
transform 1 0 27324 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1632082664
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_285
timestamp 1632082664
transform 1 0 27324 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_281
timestamp 1632082664
transform 1 0 26956 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_281
timestamp 1632082664
transform 1 0 26956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_302
timestamp 1632082664
transform 1 0 28888 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_301
timestamp 1632082664
transform 1 0 28796 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1632082664
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_309
timestamp 1632082664
transform 1 0 29532 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0847_
timestamp 1632082664
transform 1 0 30176 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0825_
timestamp 1632082664
transform 1 0 29992 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_34_313
timestamp 1632082664
transform 1 0 29900 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_330
timestamp 1632082664
transform 1 0 31464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_332
timestamp 1632082664
transform 1 0 31648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_313
timestamp 1632082664
transform 1 0 29900 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_104_clk
timestamp 1632082664
transform 1 0 31832 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_34_354
timestamp 1632082664
transform 1 0 33672 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0781_
timestamp 1632082664
transform 1 0 32476 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1632082664
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_337
timestamp 1632082664
transform 1 0 32108 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_103_clk
timestamp 1632082664
transform 1 0 34960 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_33_357
timestamp 1632082664
transform 1 0 33948 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1632082664
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1632082664
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1632082664
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_365
timestamp 1632082664
transform 1 0 34684 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1658_
timestamp 1632082664
transform 1 0 37260 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0693_
timestamp 1632082664
transform 1 0 36156 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1632082664
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_377
timestamp 1632082664
transform 1 0 35788 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_388
timestamp 1632082664
transform 1 0 36800 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_409
timestamp 1632082664
transform 1 0 38732 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_397
timestamp 1632082664
transform 1 0 37628 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_409
timestamp 1632082664
transform 1 0 38732 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_421
timestamp 1632082664
transform 1 0 39836 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1649_
timestamp 1632082664
transform 1 0 40480 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0605_
timestamp 1632082664
transform 1 0 39836 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_34_437
timestamp 1632082664
transform 1 0 41308 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1632082664
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_427
timestamp 1632082664
transform 1 0 40388 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_417
timestamp 1632082664
transform 1 0 39468 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1645_
timestamp 1632082664
transform 1 0 42412 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0550_
timestamp 1632082664
transform 1 0 42688 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1632082664
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_444
timestamp 1632082664
transform 1 0 41952 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_449
timestamp 1632082664
transform 1 0 42412 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_477
timestamp 1632082664
transform 1 0 44988 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_468
timestamp 1632082664
transform 1 0 44160 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_465
timestamp 1632082664
transform 1 0 43884 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1632082664
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_477
timestamp 1632082664
transform 1 0 44988 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1632082664
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0297_
timestamp 1632082664
transform 1 0 45632 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0286_
timestamp 1632082664
transform 1 0 45356 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_34_483
timestamp 1632082664
transform 1 0 45540 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_500
timestamp 1632082664
transform 1 0 47104 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_505
timestamp 1632082664
transform 1 0 47564 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0341_
timestamp 1632082664
transform 1 0 47748 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0319_
timestamp 1632082664
transform 1 0 47472 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_34_520
timestamp 1632082664
transform 1 0 48944 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1632082664
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1632082664
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_87_clk
timestamp 1632082664
transform 1 0 49956 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_33_523
timestamp 1632082664
transform 1 0 49220 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0374_
timestamp 1632082664
transform 1 0 50140 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1632082664
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_551
timestamp 1632082664
transform 1 0 51796 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1912_
timestamp 1632082664
transform 1 0 52716 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1909_
timestamp 1632082664
transform 1 0 51980 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1632082664
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1632082664
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_549
timestamp 1632082664
transform 1 0 51612 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1632082664
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1913_
timestamp 1632082664
transform 1 0 54556 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_34_569
timestamp 1632082664
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_577
timestamp 1632082664
transform 1 0 54188 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1916_
timestamp 1632082664
transform 1 0 55292 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_33_597
timestamp 1632082664
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1632082664
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1632082664
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1632082664
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1919_
timestamp 1632082664
transform 1 0 57132 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_33_617
timestamp 1632082664
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1632082664
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1632082664
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_625
timestamp 1632082664
transform 1 0 58604 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_605
timestamp 1632082664
transform 1 0 56764 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_629
timestamp 1632082664
transform 1 0 58972 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_629
timestamp 1632082664
transform 1 0 58972 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1632082664
transform -1 0 59340 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1632082664
transform -1 0 59340 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_3
timestamp 1632082664
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1249_
timestamp 1632082664
transform 1 0 2024 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_35_9
timestamp 1632082664
transform 1 0 1932 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1632082664
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1251_
timestamp 1632082664
transform 1 0 3864 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_35_26
timestamp 1632082664
transform 1 0 3496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_57
timestamp 1632082664
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_46
timestamp 1632082664
transform 1 0 5336 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1632082664
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1632082664
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1262_
timestamp 1632082664
transform 1 0 6992 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_35_80
timestamp 1632082664
transform 1 0 8464 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_63
timestamp 1632082664
transform 1 0 6900 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_104
timestamp 1632082664
transform 1 0 10672 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_92
timestamp 1632082664
transform 1 0 9568 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_113
timestamp 1632082664
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1206_
timestamp 1632082664
transform 1 0 12236 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1632082664
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_137
timestamp 1632082664
transform 1 0 13708 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_145
timestamp 1632082664
transform 1 0 14444 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1202_
timestamp 1632082664
transform 1 0 14720 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1632082664
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1203_
timestamp 1632082664
transform 1 0 16652 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1632082664
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_185
timestamp 1632082664
transform 1 0 18124 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1798_
timestamp 1632082664
transform 1 0 18492 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_35_205
timestamp 1632082664
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1632082664
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1807_
timestamp 1632082664
transform 1 0 21804 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1632082664
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1632082664
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1632082664
transform 1 0 23736 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_35_245
timestamp 1632082664
transform 1 0 23644 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_241
timestamp 1632082664
transform 1 0 23276 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_262
timestamp 1632082664
transform 1 0 25208 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_281
timestamp 1632082664
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_274
timestamp 1632082664
transform 1 0 26312 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0968_
timestamp 1632082664
transform 1 0 27600 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1632082664
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_287
timestamp 1632082664
transform 1 0 27508 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_304
timestamp 1632082664
transform 1 0 29072 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0814_
timestamp 1632082664
transform 1 0 30176 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1632082664
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0759_
timestamp 1632082664
transform 1 0 33488 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1632082664
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1632082664
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_349
timestamp 1632082664
transform 1 0 33212 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0704_
timestamp 1632082664
transform 1 0 35328 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_35_368
timestamp 1632082664
transform 1 0 34960 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1632082664
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1632082664
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_388
timestamp 1632082664
transform 1 0 36800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0627_
timestamp 1632082664
transform 1 0 38640 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_35_405
timestamp 1632082664
transform 1 0 38364 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0583_
timestamp 1632082664
transform 1 0 40480 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_35_424
timestamp 1632082664
transform 1 0 40112 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_79_clk
timestamp 1632082664
transform 1 0 42780 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1632082664
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_449
timestamp 1632082664
transform 1 0 42412 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_444
timestamp 1632082664
transform 1 0 41952 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1646_
timestamp 1632082664
transform 1 0 44988 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_35_473
timestamp 1632082664
transform 1 0 44620 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_493
timestamp 1632082664
transform 1 0 46460 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_505
timestamp 1632082664
transform 1 0 47564 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0396_
timestamp 1632082664
transform 1 0 48300 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1632082664
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_501
timestamp 1632082664
transform 1 0 47196 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0385_
timestamp 1632082664
transform 1 0 50140 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_35_529
timestamp 1632082664
transform 1 0 49772 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_549
timestamp 1632082664
transform 1 0 51612 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1632082664
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_561
timestamp 1632082664
transform 1 0 52716 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_557
timestamp 1632082664
transform 1 0 52348 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1908_
timestamp 1632082664
transform 1 0 53176 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_35_565
timestamp 1632082664
transform 1 0 53084 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_582
timestamp 1632082664
transform 1 0 54648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1917_
timestamp 1632082664
transform 1 0 55016 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_35_602
timestamp 1632082664
transform 1 0 56488 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_614
timestamp 1632082664
transform 1 0 57592 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_617
timestamp 1632082664
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1632082664
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_629
timestamp 1632082664
transform 1 0 58972 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1632082664
transform -1 0 59340 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1248_
timestamp 1632082664
transform 1 0 1840 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_36_7
timestamp 1632082664
transform 1 0 1748 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1632082664
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1632082664
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1250_
timestamp 1632082664
transform 1 0 3772 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1632082664
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1632082664
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_57
timestamp 1632082664
transform 1 0 6348 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_45
timestamp 1632082664
transform 1 0 5244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_69
timestamp 1632082664
transform 1 0 7452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_81
timestamp 1632082664
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1632082664
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1632082664
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1632082664
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1208_
timestamp 1632082664
transform 1 0 11592 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_36_113
timestamp 1632082664
transform 1 0 11500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_109
timestamp 1632082664
transform 1 0 11132 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_130
timestamp 1632082664
transform 1 0 13064 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1632082664
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1632082664
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1632082664
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_153
timestamp 1632082664
transform 1 0 15180 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1199_
timestamp 1632082664
transform 1 0 15732 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_36_187
timestamp 1632082664
transform 1 0 18308 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_175
timestamp 1632082664
transform 1 0 17204 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1801_
timestamp 1632082664
transform 1 0 19228 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1632082664
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1632082664
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1805_
timestamp 1632082664
transform 1 0 21068 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_36_213
timestamp 1632082664
transform 1 0 20700 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1632082664
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_233
timestamp 1632082664
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 1632082664
transform 1 0 24380 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_36_269
timestamp 1632082664
transform 1 0 25852 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1632082664
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1632082664
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_281
timestamp 1632082664
transform 1 0 26956 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0979_
timestamp 1632082664
transform 1 0 27600 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_36_287
timestamp 1632082664
transform 1 0 27508 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1632082664
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1632082664
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1632082664
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0792_
timestamp 1632082664
transform 1 0 30912 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_36_321
timestamp 1632082664
transform 1 0 30636 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0737_
timestamp 1632082664
transform 1 0 32752 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_36_340
timestamp 1632082664
transform 1 0 32384 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1632082664
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1632082664
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1632082664
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0671_
timestamp 1632082664
transform 1 0 36064 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_36_377
timestamp 1632082664
transform 1 0 35788 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0649_
timestamp 1632082664
transform 1 0 37904 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_36_416
timestamp 1632082664
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_396
timestamp 1632082664
transform 1 0 37536 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0561_
timestamp 1632082664
transform 1 0 41216 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1632082664
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1632082664
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_433
timestamp 1632082664
transform 1 0 40940 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0528_
timestamp 1632082664
transform 1 0 43056 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_36_452
timestamp 1632082664
transform 1 0 42688 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_477
timestamp 1632082664
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1632082664
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_472
timestamp 1632082664
transform 1 0 44528 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_80_clk
timestamp 1632082664
transform 1 0 46276 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_36_489
timestamp 1632082664
transform 1 0 46092 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_511
timestamp 1632082664
transform 1 0 48116 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_523
timestamp 1632082664
transform 1 0 49220 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1905_
timestamp 1632082664
transform 1 0 50600 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1632082664
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_537
timestamp 1632082664
transform 1 0 50508 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1632082664
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_533
timestamp 1632082664
transform 1 0 50140 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1907_
timestamp 1632082664
transform 1 0 52440 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_36_554
timestamp 1632082664
transform 1 0 52072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_574
timestamp 1632082664
transform 1 0 53912 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_85_clk
timestamp 1632082664
transform 1 0 56120 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_36_589
timestamp 1632082664
transform 1 0 55292 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_586
timestamp 1632082664
transform 1 0 55016 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1632082664
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_597
timestamp 1632082664
transform 1 0 56028 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_618
timestamp 1632082664
transform 1 0 57960 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1632082664
transform -1 0 59340 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_3
timestamp 1632082664
transform 1 0 1380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1247_
timestamp 1632082664
transform 1 0 2208 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_37_11
timestamp 1632082664
transform 1 0 2116 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1632082664
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_40
timestamp 1632082664
transform 1 0 4784 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_28
timestamp 1632082664
transform 1 0 3680 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1632082664
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1632082664
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1632082664
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_81
timestamp 1632082664
transform 1 0 8556 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1632082664
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_104
timestamp 1632082664
transform 1 0 10672 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1233_
timestamp 1632082664
transform 1 0 9200 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_37_87
timestamp 1632082664
transform 1 0 9108 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1632082664
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1210_
timestamp 1632082664
transform 1 0 11684 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1632082664
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_131
timestamp 1632082664
transform 1 0 13156 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_143
timestamp 1632082664
transform 1 0 14260 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1200_
timestamp 1632082664
transform 1 0 14720 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_37_147
timestamp 1632082664
transform 1 0 14628 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1632082664
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1802_
timestamp 1632082664
transform 1 0 18124 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1632082664
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1632082664
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_181
timestamp 1632082664
transform 1 0 17756 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_201
timestamp 1632082664
transform 1 0 19596 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_clk
timestamp 1632082664
transform 1 0 20884 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_218
timestamp 1632082664
transform 1 0 21160 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_213
timestamp 1632082664
transform 1 0 20700 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1809_
timestamp 1632082664
transform 1 0 21804 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1632082664
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1632082664
transform 1 0 23736 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_37_245
timestamp 1632082664
transform 1 0 23644 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_241
timestamp 1632082664
transform 1 0 23276 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_262
timestamp 1632082664
transform 1 0 25208 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_107_clk
timestamp 1632082664
transform 1 0 27324 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_37_274
timestamp 1632082664
transform 1 0 26312 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1632082664
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_281
timestamp 1632082664
transform 1 0 26956 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1632082664
transform 1 0 29532 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_37_305
timestamp 1632082664
transform 1 0 29164 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_325
timestamp 1632082664
transform 1 0 31004 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_333
timestamp 1632082664
transform 1 0 31740 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0748_
timestamp 1632082664
transform 1 0 33488 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1632082664
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1632082664
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_349
timestamp 1632082664
transform 1 0 33212 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0682_
timestamp 1632082664
transform 1 0 35328 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_37_368
timestamp 1632082664
transform 1 0 34960 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1632082664
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1632082664
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_388
timestamp 1632082664
transform 1 0 36800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0616_
timestamp 1632082664
transform 1 0 38456 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_37_405
timestamp 1632082664
transform 1 0 38364 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0594_
timestamp 1632082664
transform 1 0 40296 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_37_422
timestamp 1632082664
transform 1 0 39928 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_449
timestamp 1632082664
transform 1 0 42412 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_442
timestamp 1632082664
transform 1 0 41768 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0517_
timestamp 1632082664
transform 1 0 42964 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1632082664
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0495_
timestamp 1632082664
transform 1 0 44804 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_37_471
timestamp 1632082664
transform 1 0 44436 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_491
timestamp 1632082664
transform 1 0 46276 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_505
timestamp 1632082664
transform 1 0 47564 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0407_
timestamp 1632082664
transform 1 0 48208 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1632082664
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_511
timestamp 1632082664
transform 1 0 48116 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1632082664
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1904_
timestamp 1632082664
transform 1 0 50140 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_37_532
timestamp 1632082664
transform 1 0 50048 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_528
timestamp 1632082664
transform 1 0 49680 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_549
timestamp 1632082664
transform 1 0 51612 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1914_
timestamp 1632082664
transform 1 0 52716 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1632082664
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_557
timestamp 1632082664
transform 1 0 52348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_577
timestamp 1632082664
transform 1 0 54188 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_589
timestamp 1632082664
transform 1 0 55292 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1922_
timestamp 1632082664
transform 1 0 55844 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_37_617
timestamp 1632082664
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1632082664
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1632082664
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_611
timestamp 1632082664
transform 1 0 57316 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_629
timestamp 1632082664
transform 1 0 58972 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1632082664
transform -1 0 59340 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1246_
timestamp 1632082664
transform 1 0 1840 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_38_7
timestamp 1632082664
transform 1 0 1748 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_3
timestamp 1632082664
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1632082664
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1632082664
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1632082664
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1632082664
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_41
timestamp 1632082664
transform 1 0 4876 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1237_
timestamp 1632082664
transform 1 0 5152 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_60
timestamp 1632082664
transform 1 0 6624 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1235_
timestamp 1632082664
transform 1 0 6992 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1632082664
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1232_
timestamp 1632082664
transform 1 0 9292 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1632082664
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_85
timestamp 1632082664
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_clk
timestamp 1632082664
transform 1 0 11776 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_38_105
timestamp 1632082664
transform 1 0 10764 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_113
timestamp 1632082664
transform 1 0 11500 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1632082664
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1632082664
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1632082664
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1197_
timestamp 1632082664
transform 1 0 15456 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_38_153
timestamp 1632082664
transform 1 0 15180 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1194_
timestamp 1632082664
transform 1 0 17296 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_172
timestamp 1632082664
transform 1 0 16928 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1806_
timestamp 1632082664
transform 1 0 19228 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1632082664
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1632082664
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1808_
timestamp 1632082664
transform 1 0 21068 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_213
timestamp 1632082664
transform 1 0 20700 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1632082664
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_233
timestamp 1632082664
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1632082664
transform 1 0 24380 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1632082664
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1632082664
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_269
timestamp 1632082664
transform 1 0 25852 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1823_
timestamp 1632082664
transform 1 0 26220 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1632082664
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1632082664
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1632082664
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1632082664
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1632082664
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0803_
timestamp 1632082664
transform 1 0 30912 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_38_321
timestamp 1632082664
transform 1 0 30636 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0770_
timestamp 1632082664
transform 1 0 32752 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_340
timestamp 1632082664
transform 1 0 32384 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_365
timestamp 1632082664
transform 1 0 34684 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0715_
timestamp 1632082664
transform 1 0 35236 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1632082664
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1632082664
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_387
timestamp 1632082664
transform 1 0 36708 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_395
timestamp 1632082664
transform 1 0 37444 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1632082664
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0660_
timestamp 1632082664
transform 1 0 37628 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_clk
timestamp 1632082664
transform 1 0 40388 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_430
timestamp 1632082664
transform 1 0 40664 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_421
timestamp 1632082664
transform 1 0 39836 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0572_
timestamp 1632082664
transform 1 0 41216 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1632082664
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1632082664
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0539_
timestamp 1632082664
transform 1 0 43056 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_452
timestamp 1632082664
transform 1 0 42688 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_477
timestamp 1632082664
transform 1 0 44988 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1632082664
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_472
timestamp 1632082664
transform 1 0 44528 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_499
timestamp 1632082664
transform 1 0 47012 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0473_
timestamp 1632082664
transform 1 0 45540 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_38_507
timestamp 1632082664
transform 1 0 47748 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0418_
timestamp 1632082664
transform 1 0 47932 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1632082664
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1903_
timestamp 1632082664
transform 1 0 50140 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1632082664
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1632082664
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1906_
timestamp 1632082664
transform 1 0 51980 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_549
timestamp 1632082664
transform 1 0 51612 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1632082664
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_569
timestamp 1632082664
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_601
timestamp 1632082664
transform 1 0 56396 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_589
timestamp 1632082664
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1632082664
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1632082664
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1920_
timestamp 1632082664
transform 1 0 57132 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_625
timestamp 1632082664
transform 1 0 58604 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_629
timestamp 1632082664
transform 1 0 58972 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1632082664
transform -1 0 59340 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_3
timestamp 1632082664
transform 1 0 1380 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_11
timestamp 1632082664
transform 1 0 2116 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1245_
timestamp 1632082664
transform 1 0 2300 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1244_
timestamp 1632082664
transform 1 0 1840 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_40_7
timestamp 1632082664
transform 1 0 1748 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 1632082664
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1632082664
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1632082664
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_29
timestamp 1632082664
transform 1 0 3772 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1238_
timestamp 1632082664
transform 1 0 4416 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1632082664
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1632082664
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_35
timestamp 1632082664
transform 1 0 4324 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_41
timestamp 1632082664
transform 1 0 4876 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_24
timestamp 1632082664
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_clk
timestamp 1632082664
transform 1 0 5244 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1632082664
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1632082664
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1632082664
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1632082664
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1234_
timestamp 1632082664
transform 1 0 7544 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1632082664
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1632082664
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_69
timestamp 1632082664
transform 1 0 7452 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1231_
timestamp 1632082664
transform 1 0 9384 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1230_
timestamp 1632082664
transform 1 0 9292 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1632082664
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_85
timestamp 1632082664
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_86
timestamp 1632082664
transform 1 0 9016 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_clk
timestamp 1632082664
transform 1 0 11408 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_105
timestamp 1632082664
transform 1 0 10764 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_106
timestamp 1632082664
transform 1 0 10856 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1212_
timestamp 1632082664
transform 1 0 12052 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1211_
timestamp 1632082664
transform 1 0 11868 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1632082664
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_111
timestamp 1632082664
transform 1 0 11316 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_115
timestamp 1632082664
transform 1 0 11684 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 1632082664
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1632082664
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_133
timestamp 1632082664
transform 1 0 13340 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1632082664
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1632082664
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_135
timestamp 1632082664
transform 1 0 13524 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_145
timestamp 1632082664
transform 1 0 14444 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1198_
timestamp 1632082664
transform 1 0 14720 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1196_
timestamp 1632082664
transform 1 0 15456 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1632082664
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_153
timestamp 1632082664
transform 1 0 15180 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_169
timestamp 1632082664
transform 1 0 16652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1193_
timestamp 1632082664
transform 1 0 17388 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1192_
timestamp 1632082664
transform 1 0 17296 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1632082664
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_172
timestamp 1632082664
transform 1 0 16928 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1632082664
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1189_
timestamp 1632082664
transform 1 0 19228 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1188_
timestamp 1632082664
transform 1 0 19412 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1632082664
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1632082664
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_193
timestamp 1632082664
transform 1 0 18860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_213
timestamp 1632082664
transform 1 0 20700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1812_
timestamp 1632082664
transform 1 0 21804 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1810_
timestamp 1632082664
transform 1 0 21252 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1632082664
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_215
timestamp 1632082664
transform 1 0 20884 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1632082664
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_241
timestamp 1632082664
transform 1 0 23276 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 1632082664
transform 1 0 24104 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_40_235
timestamp 1632082664
transform 1 0 22724 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_249
timestamp 1632082664
transform 1 0 24012 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1632082664
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1816_
timestamp 1632082664
transform 1 0 24380 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_39_266
timestamp 1632082664
transform 1 0 25576 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1632082664
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1632082664
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_269
timestamp 1632082664
transform 1 0 25852 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1632082664
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1820_
timestamp 1632082664
transform 1 0 26956 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1819_
timestamp 1632082664
transform 1 0 26220 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_40_289
timestamp 1632082664
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1632082664
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1632082664
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1632082664
transform 1 0 29532 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1632082664
transform 1 0 28796 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1632082664
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1632082664
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_297
timestamp 1632082664
transform 1 0 28428 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1632082664
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1832_
timestamp 1632082664
transform 1 0 31372 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1632082664
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_325
timestamp 1632082664
transform 1 0 31004 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1850_
timestamp 1632082664
transform 1 0 32108 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1632082664
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1632082664
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1632082664
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_353
timestamp 1632082664
transform 1 0 33580 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1632082664
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1856_
timestamp 1632082664
transform 1 0 33948 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1854_
timestamp 1632082664
transform 1 0 34684 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1632082664
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1632082664
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1632082664
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1632082664
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1862_
timestamp 1632082664
transform 1 0 36524 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1632082664
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1632082664
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1632082664
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_381
timestamp 1632082664
transform 1 0 36156 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1632082664
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1632082664
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0638_
timestamp 1632082664
transform 1 0 38548 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1632082664
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1994_
timestamp 1632082664
transform 1 0 40480 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1868_
timestamp 1632082664
transform 1 0 39836 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1632082664
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1632082664
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_427
timestamp 1632082664
transform 1 0 40388 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_437
timestamp 1632082664
transform 1 0 41308 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_423
timestamp 1632082664
transform 1 0 40020 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1873_
timestamp 1632082664
transform 1 0 41676 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1632082664
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1632082664
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1632082664
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_444
timestamp 1632082664
transform 1 0 41952 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1632082664
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0506_
timestamp 1632082664
transform 1 0 43792 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0484_
timestamp 1632082664
transform 1 0 44988 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1632082664
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1632082664
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_461
timestamp 1632082664
transform 1 0 43516 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0462_
timestamp 1632082664
transform 1 0 45632 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_40_493
timestamp 1632082664
transform 1 0 46460 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_500
timestamp 1632082664
transform 1 0 47104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_480
timestamp 1632082664
transform 1 0 45264 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0440_
timestamp 1632082664
transform 1 0 47564 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0429_
timestamp 1632082664
transform 1 0 47564 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1632082664
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_clk
timestamp 1632082664
transform 1 0 49404 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1902_
timestamp 1632082664
transform 1 0 50140 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1901_
timestamp 1632082664
transform 1 0 49404 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_39_541
timestamp 1632082664
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1632082664
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_528
timestamp 1632082664
transform 1 0 49680 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_521
timestamp 1632082664
transform 1 0 49036 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_521
timestamp 1632082664
transform 1 0 49036 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_561
timestamp 1632082664
transform 1 0 52716 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1632082664
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_549
timestamp 1632082664
transform 1 0 51612 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1632082664
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1632082664
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_561
timestamp 1632082664
transform 1 0 52716 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1632082664
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1936_
timestamp 1632082664
transform 1 0 53360 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1935_
timestamp 1632082664
transform 1 0 53084 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_39_567
timestamp 1632082664
transform 1 0 53268 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1953_
timestamp 1632082664
transform 1 0 55292 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1924_
timestamp 1632082664
transform 1 0 55936 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_39_584
timestamp 1632082664
transform 1 0 54832 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1632082664
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1632082664
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1923_
timestamp 1632082664
transform 1 0 57132 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_39_617
timestamp 1632082664
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1632082664
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_625
timestamp 1632082664
transform 1 0 58604 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_605
timestamp 1632082664
transform 1 0 56764 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_612
timestamp 1632082664
transform 1 0 57408 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_629
timestamp 1632082664
transform 1 0 58972 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_629
timestamp 1632082664
transform 1 0 58972 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1632082664
transform -1 0 59340 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1632082664
transform -1 0 59340 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_3
timestamp 1632082664
transform 1 0 1380 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1243_
timestamp 1632082664
transform 1 0 1932 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1632082664
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1241_
timestamp 1632082664
transform 1 0 3772 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_25
timestamp 1632082664
transform 1 0 3404 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_45
timestamp 1632082664
transform 1 0 5244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1236_
timestamp 1632082664
transform 1 0 6348 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1632082664
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 1632082664
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_73
timestamp 1632082664
transform 1 0 7820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_102
timestamp 1632082664
transform 1 0 10488 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1229_
timestamp 1632082664
transform 1 0 9016 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_41_85
timestamp 1632082664
transform 1 0 8924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_113
timestamp 1632082664
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1632082664
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1213_
timestamp 1632082664
transform 1 0 12144 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1632082664
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_119
timestamp 1632082664
transform 1 0 12052 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_136
timestamp 1632082664
transform 1 0 13616 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1195_
timestamp 1632082664
transform 1 0 14720 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1632082664
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_169
timestamp 1632082664
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1191_
timestamp 1632082664
transform 1 0 17296 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1632082664
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_175
timestamp 1632082664
transform 1 0 17204 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_192
timestamp 1632082664
transform 1 0 18768 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1187_
timestamp 1632082664
transform 1 0 19780 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_41_200
timestamp 1632082664
transform 1 0 19504 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1813_
timestamp 1632082664
transform 1 0 21804 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1632082664
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1632082664
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_219
timestamp 1632082664
transform 1 0 21252 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_241
timestamp 1632082664
transform 1 0 23276 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 1632082664
transform 1 0 24104 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_41_249
timestamp 1632082664
transform 1 0 24012 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_266
timestamp 1632082664
transform 1 0 25576 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1632082664
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1821_
timestamp 1632082664
transform 1 0 26956 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1632082664
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1828_
timestamp 1632082664
transform 1 0 28796 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_297
timestamp 1632082664
transform 1 0 28428 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1632082664
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1632082664
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1848_
timestamp 1632082664
transform 1 0 32108 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1632082664
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1632082664
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_353
timestamp 1632082664
transform 1 0 33580 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1849_
timestamp 1632082664
transform 1 0 33948 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1632082664
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1632082664
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1859_
timestamp 1632082664
transform 1 0 37260 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1632082664
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1632082664
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1863_
timestamp 1632082664
transform 1 0 39100 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_409
timestamp 1632082664
transform 1 0 38732 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1632082664
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1632082664
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_449
timestamp 1632082664
transform 1 0 42412 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1874_
timestamp 1632082664
transform 1 0 43148 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1632082664
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1632082664
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1875_
timestamp 1632082664
transform 1 0 44988 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_473
timestamp 1632082664
transform 1 0 44620 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_493
timestamp 1632082664
transform 1 0 46460 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0451_
timestamp 1632082664
transform 1 0 47564 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1632082664
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_501
timestamp 1632082664
transform 1 0 47196 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1900_
timestamp 1632082664
transform 1 0 49404 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_41_541
timestamp 1632082664
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_521
timestamp 1632082664
transform 1 0 49036 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1632082664
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_561
timestamp 1632082664
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1632082664
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1632082664
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1933_
timestamp 1632082664
transform 1 0 54096 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_41_573
timestamp 1632082664
transform 1 0 53820 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1925_
timestamp 1632082664
transform 1 0 55936 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_592
timestamp 1632082664
transform 1 0 55568 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_617
timestamp 1632082664
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1632082664
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_612
timestamp 1632082664
transform 1 0 57408 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_629
timestamp 1632082664
transform 1 0 58972 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1632082664
transform -1 0 59340 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1632082664
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1632082664
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1632082664
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_29
timestamp 1632082664
transform 1 0 3772 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1240_
timestamp 1632082664
transform 1 0 4508 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1632082664
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1632082664
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1239_
timestamp 1632082664
transform 1 0 6348 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_42_53
timestamp 1632082664
transform 1 0 5980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_73
timestamp 1632082664
transform 1 0 7820 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_81
timestamp 1632082664
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1228_
timestamp 1632082664
transform 1 0 8924 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_42_101
timestamp 1632082664
transform 1 0 10396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1632082664
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_113
timestamp 1632082664
transform 1 0 11500 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1214_
timestamp 1632082664
transform 1 0 12144 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_42_119
timestamp 1632082664
transform 1 0 12052 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_141
timestamp 1632082664
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1632082664
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1632082664
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1217_
timestamp 1632082664
transform 1 0 15088 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_42_149
timestamp 1632082664
transform 1 0 14812 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_168
timestamp 1632082664
transform 1 0 16560 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1190_
timestamp 1632082664
transform 1 0 17296 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_42_197
timestamp 1632082664
transform 1 0 19228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1186_
timestamp 1632082664
transform 1 0 19872 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1632082664
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_203
timestamp 1632082664
transform 1 0 19780 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1632082664
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1814_
timestamp 1632082664
transform 1 0 21712 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_42_220
timestamp 1632082664
transform 1 0 21344 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_240
timestamp 1632082664
transform 1 0 23184 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1817_
timestamp 1632082664
transform 1 0 24380 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1632082664
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_269
timestamp 1632082664
transform 1 0 25852 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1818_
timestamp 1632082664
transform 1 0 26220 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1632082664
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1632082664
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1632082664
transform 1 0 29532 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1632082664
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1632082664
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1845_
timestamp 1632082664
transform 1 0 31372 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_42_325
timestamp 1632082664
transform 1 0 31004 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1632082664
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1632082664
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1853_
timestamp 1632082664
transform 1 0 34684 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1632082664
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1632082664
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1858_
timestamp 1632082664
transform 1 0 36524 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_42_381
timestamp 1632082664
transform 1 0 36156 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1632082664
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1632082664
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1867_
timestamp 1632082664
transform 1 0 39836 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1632082664
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1632082664
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_437
timestamp 1632082664
transform 1 0 41308 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1871_
timestamp 1632082664
transform 1 0 41676 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1632082664
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1632082664
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1879_
timestamp 1632082664
transform 1 0 44988 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1632082664
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1632082664
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1883_
timestamp 1632082664
transform 1 0 46828 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_42_493
timestamp 1632082664
transform 1 0 46460 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_513
timestamp 1632082664
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1632082664
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1898_
timestamp 1632082664
transform 1 0 50140 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1632082664
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1632082664
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_561
timestamp 1632082664
transform 1 0 52716 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_549
timestamp 1632082664
transform 1 0 51612 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1937_
timestamp 1632082664
transform 1 0 53360 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_42_567
timestamp 1632082664
transform 1 0 53268 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_589
timestamp 1632082664
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1632082664
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_601
timestamp 1632082664
transform 1 0 56396 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_584
timestamp 1632082664
transform 1 0 54832 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_621
timestamp 1632082664
transform 1 0 58236 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1926_
timestamp 1632082664
transform 1 0 56764 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_42_629
timestamp 1632082664
transform 1 0 58972 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1632082664
transform -1 0 59340 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1632082664
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1632082664
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1632082664
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_27
timestamp 1632082664
transform 1 0 3588 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1242_
timestamp 1632082664
transform 1 0 4416 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_43_35
timestamp 1632082664
transform 1 0 4324 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_57
timestamp 1632082664
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1632082664
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1632082664
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1225_
timestamp 1632082664
transform 1 0 7084 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_43_81
timestamp 1632082664
transform 1 0 8556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_101
timestamp 1632082664
transform 1 0 10396 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1227_
timestamp 1632082664
transform 1 0 8924 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1632082664
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1215_
timestamp 1632082664
transform 1 0 12144 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1632082664
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_119
timestamp 1632082664
transform 1 0 12052 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_109
timestamp 1632082664
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1216_
timestamp 1632082664
transform 1 0 13984 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_43_136
timestamp 1632082664
transform 1 0 13616 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_156
timestamp 1632082664
transform 1 0 15456 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1219_
timestamp 1632082664
transform 1 0 16652 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1632082664
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_185
timestamp 1632082664
transform 1 0 18124 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_clk
timestamp 1632082664
transform 1 0 18584 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_43_189
timestamp 1632082664
transform 1 0 18492 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1632082664
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1815_
timestamp 1632082664
transform 1 0 21804 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_43_210
timestamp 1632082664
transform 1 0 20424 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1632082664
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_241
timestamp 1632082664
transform 1 0 23276 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp 1632082664
transform 1 0 24104 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_43_249
timestamp 1632082664
transform 1 0 24012 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_266
timestamp 1632082664
transform 1 0 25576 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1632082664
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1632082664
transform 1 0 26956 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1632082664
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_297
timestamp 1632082664
transform 1 0 28428 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_309
timestamp 1632082664
transform 1 0 29532 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_330
timestamp 1632082664
transform 1 0 31464 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1632082664
transform 1 0 29992 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_43_313
timestamp 1632082664
transform 1 0 29900 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_105_clk
timestamp 1632082664
transform 1 0 32936 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_43_337
timestamp 1632082664
transform 1 0 32108 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1632082664
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_345
timestamp 1632082664
transform 1 0 32844 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1852_
timestamp 1632082664
transform 1 0 35144 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_43_366
timestamp 1632082664
transform 1 0 34776 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_386
timestamp 1632082664
transform 1 0 36616 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1860_
timestamp 1632082664
transform 1 0 37260 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1632082664
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1865_
timestamp 1632082664
transform 1 0 39100 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_43_409
timestamp 1632082664
transform 1 0 38732 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1632082664
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1632082664
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1872_
timestamp 1632082664
transform 1 0 42412 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1632082664
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1632082664
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1878_
timestamp 1632082664
transform 1 0 44252 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_43_465
timestamp 1632082664
transform 1 0 43884 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1632082664
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1632082664
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_81_clk
timestamp 1632082664
transform 1 0 47932 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1632082664
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1632082664
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_505
timestamp 1632082664
transform 1 0 47564 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1897_
timestamp 1632082664
transform 1 0 50140 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_43_529
timestamp 1632082664
transform 1 0 49772 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_549
timestamp 1632082664
transform 1 0 51612 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_561
timestamp 1632082664
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1632082664
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_557
timestamp 1632082664
transform 1 0 52348 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1931_
timestamp 1632082664
transform 1 0 54096 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_43_573
timestamp 1632082664
transform 1 0 53820 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1927_
timestamp 1632082664
transform 1 0 55936 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_43_592
timestamp 1632082664
transform 1 0 55568 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_617
timestamp 1632082664
transform 1 0 57868 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1632082664
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_612
timestamp 1632082664
transform 1 0 57408 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_629
timestamp 1632082664
transform 1 0 58972 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1632082664
transform -1 0 59340 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1632082664
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1632082664
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1632082664
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1632082664
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1632082664
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1632082664
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1632082664
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_53
timestamp 1632082664
transform 1 0 5980 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1224_
timestamp 1632082664
transform 1 0 6624 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_44_59
timestamp 1632082664
transform 1 0 6532 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_76
timestamp 1632082664
transform 1 0 8096 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1222_
timestamp 1632082664
transform 1 0 10304 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1632082664
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1632082664
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_97
timestamp 1632082664
transform 1 0 10028 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1218_
timestamp 1632082664
transform 1 0 12144 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_44_116
timestamp 1632082664
transform 1 0 11776 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0078_
timestamp 1632082664
transform 1 0 14076 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1632082664
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1632082664
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1220_
timestamp 1632082664
transform 1 0 15916 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_44_157
timestamp 1632082664
transform 1 0 15548 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1632082664
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_197
timestamp 1632082664
transform 1 0 19228 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1632082664
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1185_
timestamp 1632082664
transform 1 0 19872 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1632082664
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_203
timestamp 1632082664
transform 1 0 19780 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1632082664
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1177_
timestamp 1632082664
transform 1 0 21712 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_44_220
timestamp 1632082664
transform 1 0 21344 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_240
timestamp 1632082664
transform 1 0 23184 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1100_
timestamp 1632082664
transform 1 0 24380 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_44_269
timestamp 1632082664
transform 1 0 25852 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1632082664
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_281
timestamp 1632082664
transform 1 0 26956 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1835_
timestamp 1632082664
transform 1 0 27600 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_44_287
timestamp 1632082664
transform 1 0 27508 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1831_
timestamp 1632082664
transform 1 0 29532 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1632082664
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_304
timestamp 1632082664
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1843_
timestamp 1632082664
transform 1 0 31372 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_44_325
timestamp 1632082664
transform 1 0 31004 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1632082664
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1632082664
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1851_
timestamp 1632082664
transform 1 0 34684 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1632082664
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1632082664
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1857_
timestamp 1632082664
transform 1 0 36524 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_44_381
timestamp 1632082664
transform 1 0 36156 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1632082664
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1632082664
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_437
timestamp 1632082664
transform 1 0 41308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1869_
timestamp 1632082664
transform 1 0 39836 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1632082664
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1632082664
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_78_clk
timestamp 1632082664
transform 1 0 42044 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_44_465
timestamp 1632082664
transform 1 0 43884 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1880_
timestamp 1632082664
transform 1 0 44988 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1632082664
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_473
timestamp 1632082664
transform 1 0 44620 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1884_
timestamp 1632082664
transform 1 0 46828 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_44_493
timestamp 1632082664
transform 1 0 46460 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_513
timestamp 1632082664
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1632082664
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1895_
timestamp 1632082664
transform 1 0 50140 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1632082664
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1632082664
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_561
timestamp 1632082664
transform 1 0 52716 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_549
timestamp 1632082664
transform 1 0 51612 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1938_
timestamp 1632082664
transform 1 0 53360 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_44_567
timestamp 1632082664
transform 1 0 53268 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_84_clk
timestamp 1632082664
transform 1 0 56488 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_44_589
timestamp 1632082664
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1632082664
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_601
timestamp 1632082664
transform 1 0 56396 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_584
timestamp 1632082664
transform 1 0 54832 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_622
timestamp 1632082664
transform 1 0 58328 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1632082664
transform -1 0 59340 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1632082664
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1632082664
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1632082664
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1632082664
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1632082664
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1632082664
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1632082664
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1632082664
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1632082664
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_69
timestamp 1632082664
transform 1 0 7452 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1226_
timestamp 1632082664
transform 1 0 7636 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_45_99
timestamp 1632082664
transform 1 0 10212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_87
timestamp 1632082664
transform 1 0 9108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1223_
timestamp 1632082664
transform 1 0 11500 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1632082664
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1632082664
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_clk
timestamp 1632082664
transform 1 0 13524 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_45_129
timestamp 1632082664
transform 1 0 12972 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_155
timestamp 1632082664
transform 1 0 15364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0071_
timestamp 1632082664
transform 1 0 16652 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_45_185
timestamp 1632082664
transform 1 0 18124 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1632082664
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1632082664
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_197
timestamp 1632082664
transform 1 0 19228 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1184_
timestamp 1632082664
transform 1 0 19872 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_45_203
timestamp 1632082664
transform 1 0 19780 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1155_
timestamp 1632082664
transform 1 0 22080 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1632082664
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1632082664
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_225
timestamp 1632082664
transform 1 0 21804 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1111_
timestamp 1632082664
transform 1 0 23920 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_45_244
timestamp 1632082664
transform 1 0 23552 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_264
timestamp 1632082664
transform 1 0 25392 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1632082664
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1632082664
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1632082664
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_106_clk
timestamp 1632082664
transform 1 0 28704 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_45_293
timestamp 1632082664
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_299
timestamp 1632082664
transform 1 0 28612 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_320
timestamp 1632082664
transform 1 0 30544 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1632082664
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1847_
timestamp 1632082664
transform 1 0 32476 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1632082664
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_337
timestamp 1632082664
transform 1 0 32108 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_357
timestamp 1632082664
transform 1 0 33948 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0025_
timestamp 1632082664
transform 1 0 34684 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_45_381
timestamp 1632082664
transform 1 0 36156 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1632082664
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_393
timestamp 1632082664
transform 1 0 37260 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_389
timestamp 1632082664
transform 1 0 36892 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1861_
timestamp 1632082664
transform 1 0 37628 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_45_413
timestamp 1632082664
transform 1 0 39100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1870_
timestamp 1632082664
transform 1 0 39468 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_45_433
timestamp 1632082664
transform 1 0 40940 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1876_
timestamp 1632082664
transform 1 0 42412 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1632082664
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_445
timestamp 1632082664
transform 1 0 42044 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1881_
timestamp 1632082664
transform 1 0 44252 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_45_465
timestamp 1632082664
transform 1 0 43884 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1632082664
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1632082664
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1886_
timestamp 1632082664
transform 1 0 47564 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1632082664
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1632082664
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1893_
timestamp 1632082664
transform 1 0 49404 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_45_541
timestamp 1632082664
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_521
timestamp 1632082664
transform 1 0 49036 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_561
timestamp 1632082664
transform 1 0 52716 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1632082664
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1632082664
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1632082664
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1939_
timestamp 1632082664
transform 1 0 53360 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_45_567
timestamp 1632082664
transform 1 0 53268 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1929_
timestamp 1632082664
transform 1 0 55936 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_45_584
timestamp 1632082664
transform 1 0 54832 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_617
timestamp 1632082664
transform 1 0 57868 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1632082664
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_612
timestamp 1632082664
transform 1 0 57408 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_629
timestamp 1632082664
transform 1 0 58972 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1632082664
transform -1 0 59340 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1632082664
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1632082664
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1632082664
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1632082664
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1632082664
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1632082664
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1632082664
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1632082664
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1632082664
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1632082664
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1632082664
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1632082664
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_53
timestamp 1632082664
transform 1 0 5980 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0094_
timestamp 1632082664
transform 1 0 6808 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1632082664
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1632082664
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1632082664
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_61
timestamp 1632082664
transform 1 0 6716 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1632082664
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_78
timestamp 1632082664
transform 1 0 8280 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0090_
timestamp 1632082664
transform 1 0 7728 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_47_69
timestamp 1632082664
transform 1 0 7452 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0084_
timestamp 1632082664
transform 1 0 9568 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1632082664
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1632082664
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1632082664
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_88
timestamp 1632082664
transform 1 0 9200 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_109
timestamp 1632082664
transform 1 0 11132 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0081_
timestamp 1632082664
transform 1 0 12144 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1632082664
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1632082664
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_125
timestamp 1632082664
transform 1 0 12604 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1632082664
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_117
timestamp 1632082664
transform 1 0 11868 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_142
timestamp 1632082664
transform 1 0 14168 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_141
timestamp 1632082664
transform 1 0 14076 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0080_
timestamp 1632082664
transform 1 0 12696 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1632082664
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1632082664
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_149
timestamp 1632082664
transform 1 0 14812 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0074_
timestamp 1632082664
transform 1 0 14996 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0073_
timestamp 1632082664
transform 1 0 14720 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1632082664
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_187
timestamp 1632082664
transform 1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0070_
timestamp 1632082664
transform 1 0 16836 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0069_
timestamp 1632082664
transform 1 0 17020 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1632082664
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_169
timestamp 1632082664
transform 1 0 16652 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_167
timestamp 1632082664
transform 1 0 16468 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_189
timestamp 1632082664
transform 1 0 18492 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0065_
timestamp 1632082664
transform 1 0 19228 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0064_
timestamp 1632082664
transform 1 0 19228 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1632082664
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1632082664
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_225
timestamp 1632082664
transform 1 0 21804 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_225
timestamp 1632082664
transform 1 0 21804 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_213
timestamp 1632082664
transform 1 0 20700 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_213
timestamp 1632082664
transform 1 0 20700 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1632082664
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 1632082664
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_233
timestamp 1632082664
transform 1 0 22540 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1144_
timestamp 1632082664
transform 1 0 22448 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1133_
timestamp 1632082664
transform 1 0 22724 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_46_231
timestamp 1632082664
transform 1 0 22356 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1632082664
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_13_clk
timestamp 1632082664
transform 1 0 24564 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1122_
timestamp 1632082664
transform 1 0 24380 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_46_269
timestamp 1632082664
transform 1 0 25852 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1632082664
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_251
timestamp 1632082664
transform 1 0 24196 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1837_
timestamp 1632082664
transform 1 0 26956 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1836_
timestamp 1632082664
transform 1 0 26956 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1632082664
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1632082664
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_275
timestamp 1632082664
transform 1 0 26404 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_297
timestamp 1632082664
transform 1 0 28428 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1839_
timestamp 1632082664
transform 1 0 28796 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1834_
timestamp 1632082664
transform 1 0 29532 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1632082664
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_297
timestamp 1632082664
transform 1 0 28428 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_305
timestamp 1632082664
transform 1 0 29164 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1632082664
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1842_
timestamp 1632082664
transform 1 0 31372 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1632082664
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_325
timestamp 1632082664
transform 1 0 31004 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1846_
timestamp 1632082664
transform 1 0 32108 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_47_353
timestamp 1632082664
transform 1 0 33580 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1632082664
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1632082664
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1632082664
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1632082664
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0024_
timestamp 1632082664
transform 1 0 34684 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0023_
timestamp 1632082664
transform 1 0 34776 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1632082664
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_365
timestamp 1632082664
transform 1 0 34684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1632082664
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_382
timestamp 1632082664
transform 1 0 36248 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_390
timestamp 1632082664
transform 1 0 36984 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1864_
timestamp 1632082664
transform 1 0 37260 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1632082664
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_381
timestamp 1632082664
transform 1 0 36156 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1632082664
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_77_clk
timestamp 1632082664
transform 1 0 38640 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_46_409
timestamp 1632082664
transform 1 0 38732 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_405
timestamp 1632082664
transform 1 0 38364 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_421
timestamp 1632082664
transform 1 0 39836 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0003_
timestamp 1632082664
transform 1 0 40480 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_47_428
timestamp 1632082664
transform 1 0 40480 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1632082664
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_427
timestamp 1632082664
transform 1 0 40388 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_417
timestamp 1632082664
transform 1 0 39468 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_440
timestamp 1632082664
transform 1 0 41584 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1990_
timestamp 1632082664
transform 1 0 43056 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1632082664
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_444
timestamp 1632082664
transform 1 0 41952 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1632082664
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1985_
timestamp 1632082664
transform 1 0 43792 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1882_
timestamp 1632082664
transform 1 0 44988 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1632082664
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_472
timestamp 1632082664
transform 1 0 44528 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_461
timestamp 1632082664
transform 1 0 43516 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1983_
timestamp 1632082664
transform 1 0 45632 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1885_
timestamp 1632082664
transform 1 0 46828 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_47_500
timestamp 1632082664
transform 1 0 47104 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_480
timestamp 1632082664
transform 1 0 45264 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_493
timestamp 1632082664
transform 1 0 46460 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1887_
timestamp 1632082664
transform 1 0 47656 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_46_513
timestamp 1632082664
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1632082664
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_505
timestamp 1632082664
transform 1 0 47564 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1632082664
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1894_
timestamp 1632082664
transform 1 0 50140 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1891_
timestamp 1632082664
transform 1 0 49496 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1632082664
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1632082664
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_522
timestamp 1632082664
transform 1 0 49128 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_561
timestamp 1632082664
transform 1 0 52716 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_554
timestamp 1632082664
transform 1 0 52072 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_46_561
timestamp 1632082664
transform 1 0 52716 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_542
timestamp 1632082664
transform 1 0 50968 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_549
timestamp 1632082664
transform 1 0 51612 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1632082664
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1941_
timestamp 1632082664
transform 1 0 53360 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1940_
timestamp 1632082664
transform 1 0 53360 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_47_567
timestamp 1632082664
transform 1 0 53268 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_567
timestamp 1632082664
transform 1 0 53268 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1930_
timestamp 1632082664
transform 1 0 55936 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1928_
timestamp 1632082664
transform 1 0 56488 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_47_584
timestamp 1632082664
transform 1 0 54832 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_589
timestamp 1632082664
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1632082664
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_601
timestamp 1632082664
transform 1 0 56396 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_584
timestamp 1632082664
transform 1 0 54832 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_617
timestamp 1632082664
transform 1 0 57868 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_618
timestamp 1632082664
transform 1 0 57960 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1632082664
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_612
timestamp 1632082664
transform 1 0 57408 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_629
timestamp 1632082664
transform 1 0 58972 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1632082664
transform -1 0 59340 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1632082664
transform -1 0 59340 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1632082664
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1632082664
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1632082664
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1632082664
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1632082664
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_41
timestamp 1632082664
transform 1 0 4876 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1632082664
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_58
timestamp 1632082664
transform 1 0 6440 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0097_
timestamp 1632082664
transform 1 0 4968 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0091_
timestamp 1632082664
transform 1 0 6992 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1632082664
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_clk
timestamp 1632082664
transform 1 0 10672 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_48_97
timestamp 1632082664
transform 1 0 10028 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1632082664
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1632082664
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_103
timestamp 1632082664
transform 1 0 10580 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_124
timestamp 1632082664
transform 1 0 12512 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1632082664
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1632082664
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1632082664
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0072_
timestamp 1632082664
transform 1 0 15456 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_48_153
timestamp 1632082664
transform 1 0 15180 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0067_
timestamp 1632082664
transform 1 0 17296 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_48_172
timestamp 1632082664
transform 1 0 16928 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0061_
timestamp 1632082664
transform 1 0 19228 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1632082664
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1632082664
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1166_
timestamp 1632082664
transform 1 0 21804 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_48_213
timestamp 1632082664
transform 1 0 20700 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_241
timestamp 1632082664
transform 1 0 23276 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_249
timestamp 1632082664
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_253
timestamp 1632082664
transform 1 0 24380 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1840_
timestamp 1632082664
transform 1 0 25116 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1632082664
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1838_
timestamp 1632082664
transform 1 0 26956 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_48_277
timestamp 1632082664
transform 1 0 26588 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_297
timestamp 1632082664
transform 1 0 28428 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1841_
timestamp 1632082664
transform 1 0 29532 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1632082664
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_305
timestamp 1632082664
transform 1 0 29164 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_325
timestamp 1632082664
transform 1 0 31004 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0027_
timestamp 1632082664
transform 1 0 32384 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_48_337
timestamp 1632082664
transform 1 0 32108 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_356
timestamp 1632082664
transform 1 0 33856 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0021_
timestamp 1632082664
transform 1 0 34776 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1632082664
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_365
timestamp 1632082664
transform 1 0 34684 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0005_
timestamp 1632082664
transform 1 0 37352 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_48_382
timestamp 1632082664
transform 1 0 36248 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_410
timestamp 1632082664
transform 1 0 38824 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_418
timestamp 1632082664
transform 1 0 39560 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0001_
timestamp 1632082664
transform 1 0 40112 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1632082664
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_421
timestamp 1632082664
transform 1 0 39836 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1988_
timestamp 1632082664
transform 1 0 43056 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_48_440
timestamp 1632082664
transform 1 0 41584 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_452
timestamp 1632082664
transform 1 0 42688 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_477
timestamp 1632082664
transform 1 0 44988 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1632082664
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_472
timestamp 1632082664
transform 1 0 44528 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1982_
timestamp 1632082664
transform 1 0 45724 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1889_
timestamp 1632082664
transform 1 0 47564 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_48_501
timestamp 1632082664
transform 1 0 47196 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_521
timestamp 1632082664
transform 1 0 49036 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1896_
timestamp 1632082664
transform 1 0 50140 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1632082664
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_529
timestamp 1632082664
transform 1 0 49772 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_549
timestamp 1632082664
transform 1 0 51612 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_561
timestamp 1632082664
transform 1 0 52716 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_582
timestamp 1632082664
transform 1 0 54648 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1942_
timestamp 1632082664
transform 1 0 53176 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_48_565
timestamp 1632082664
transform 1 0 53084 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_601
timestamp 1632082664
transform 1 0 56396 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_589
timestamp 1632082664
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1632082664
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_624
timestamp 1632082664
transform 1 0 58512 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1934_
timestamp 1632082664
transform 1 0 57040 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_48_607
timestamp 1632082664
transform 1 0 56948 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1632082664
transform -1 0 59340 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0102_
timestamp 1632082664
transform 1 0 2576 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1632082664
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_15
timestamp 1632082664
transform 1 0 2484 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1632082664
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0098_
timestamp 1632082664
transform 1 0 4416 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_49_32
timestamp 1632082664
transform 1 0 4048 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_clk
timestamp 1632082664
transform 1 0 6716 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1632082664
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_57
timestamp 1632082664
transform 1 0 6348 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_52
timestamp 1632082664
transform 1 0 5888 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_81
timestamp 1632082664
transform 1 0 8556 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0086_
timestamp 1632082664
transform 1 0 9568 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_49_89
timestamp 1632082664
transform 1 0 9292 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1632082664
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1632082664
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_108
timestamp 1632082664
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_125
timestamp 1632082664
transform 1 0 12604 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0079_
timestamp 1632082664
transform 1 0 12880 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_49_144
timestamp 1632082664
transform 1 0 14352 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0075_
timestamp 1632082664
transform 1 0 14720 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1632082664
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_169
timestamp 1632082664
transform 1 0 16652 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0068_
timestamp 1632082664
transform 1 0 17388 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1632082664
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_12_clk
timestamp 1632082664
transform 1 0 19504 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_49_193
timestamp 1632082664
transform 1 0 18860 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_199
timestamp 1632082664
transform 1 0 19412 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_225
timestamp 1632082664
transform 1 0 21804 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1632082664
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1632082664
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_248
timestamp 1632082664
transform 1 0 23920 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0053_
timestamp 1632082664
transform 1 0 22448 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_49_231
timestamp 1632082664
transform 1 0 22356 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_270
timestamp 1632082664
transform 1 0 25944 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0049_
timestamp 1632082664
transform 1 0 24472 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1632082664
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0042_
timestamp 1632082664
transform 1 0 27232 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1632082664
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_281
timestamp 1632082664
transform 1 0 26956 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_300
timestamp 1632082664
transform 1 0 28704 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_312
timestamp 1632082664
transform 1 0 29808 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0029_
timestamp 1632082664
transform 1 0 30176 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1632082664
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_337
timestamp 1632082664
transform 1 0 32108 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0026_
timestamp 1632082664
transform 1 0 32844 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1632082664
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0020_
timestamp 1632082664
transform 1 0 34684 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_49_361
timestamp 1632082664
transform 1 0 34316 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_381
timestamp 1632082664
transform 1 0 36156 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1632082664
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_393
timestamp 1632082664
transform 1 0 37260 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_389
timestamp 1632082664
transform 1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_412
timestamp 1632082664
transform 1 0 39008 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0004_
timestamp 1632082664
transform 1 0 37536 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0002_
timestamp 1632082664
transform 1 0 39652 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_49_435
timestamp 1632082664
transform 1 0 41124 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_418
timestamp 1632082664
transform 1 0 39560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1632082664
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1632082664
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1632082664
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1984_
timestamp 1632082664
transform 1 0 43792 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_49_461
timestamp 1632082664
transform 1 0 43516 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1979_
timestamp 1632082664
transform 1 0 45632 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_49_500
timestamp 1632082664
transform 1 0 47104 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_480
timestamp 1632082664
transform 1 0 45264 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1890_
timestamp 1632082664
transform 1 0 47564 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1632082664
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1892_
timestamp 1632082664
transform 1 0 49404 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_49_541
timestamp 1632082664
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_521
timestamp 1632082664
transform 1 0 49036 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1632082664
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1632082664
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1632082664
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_561
timestamp 1632082664
transform 1 0 52716 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_83_clk
timestamp 1632082664
transform 1 0 53084 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1946_
timestamp 1632082664
transform 1 0 55292 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_49_585
timestamp 1632082664
transform 1 0 54924 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_605
timestamp 1632082664
transform 1 0 56764 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_617
timestamp 1632082664
transform 1 0 57868 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1632082664
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_613
timestamp 1632082664
transform 1 0 57500 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_49_629
timestamp 1632082664
transform 1 0 58972 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1632082664
transform -1 0 59340 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1632082664
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1632082664
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1632082664
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1632082664
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1632082664
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1632082664
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_41
timestamp 1632082664
transform 1 0 4876 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0096_
timestamp 1632082664
transform 1 0 5152 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_50_60
timestamp 1632082664
transform 1 0 6624 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0093_
timestamp 1632082664
transform 1 0 6992 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_50_80
timestamp 1632082664
transform 1 0 8464 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0085_
timestamp 1632082664
transform 1 0 10028 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1632082664
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1632082664
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0082_
timestamp 1632082664
transform 1 0 11868 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_50_113
timestamp 1632082664
transform 1 0 11500 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1632082664
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1632082664
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1632082664
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1632082664
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_163
timestamp 1632082664
transform 1 0 16100 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0076_
timestamp 1632082664
transform 1 0 14628 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_50_171
timestamp 1632082664
transform 1 0 16836 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1221_
timestamp 1632082664
transform 1 0 17020 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1632082664
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1632082664
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1632082664
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1632082664
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0057_
timestamp 1632082664
transform 1 0 20608 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_50_228
timestamp 1632082664
transform 1 0 22080 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_209
timestamp 1632082664
transform 1 0 20332 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0052_
timestamp 1632082664
transform 1 0 22448 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1632082664
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0045_
timestamp 1632082664
transform 1 0 25760 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1632082664
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1632082664
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_265
timestamp 1632082664
transform 1 0 25484 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0039_
timestamp 1632082664
transform 1 0 27600 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_50_284
timestamp 1632082664
transform 1 0 27232 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1632082664
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_309
timestamp 1632082664
transform 1 0 29532 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1632082664
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0032_
timestamp 1632082664
transform 1 0 29992 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_50_313
timestamp 1632082664
transform 1 0 29900 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_330
timestamp 1632082664
transform 1 0 31464 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0028_
timestamp 1632082664
transform 1 0 31832 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_50_350
timestamp 1632082664
transform 1 0 33304 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_362
timestamp 1632082664
transform 1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0019_
timestamp 1632082664
transform 1 0 34684 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1632082664
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_393
timestamp 1632082664
transform 1 0 37260 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0006_
timestamp 1632082664
transform 1 0 37444 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_50_381
timestamp 1632082664
transform 1 0 36156 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_411
timestamp 1632082664
transform 1 0 38916 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1992_
timestamp 1632082664
transform 1 0 41216 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1632082664
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1632082664
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1632082664
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_433
timestamp 1632082664
transform 1 0 40940 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1986_
timestamp 1632082664
transform 1 0 43056 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_50_452
timestamp 1632082664
transform 1 0 42688 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_477
timestamp 1632082664
transform 1 0 44988 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1632082664
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_472
timestamp 1632082664
transform 1 0 44528 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1975_
timestamp 1632082664
transform 1 0 45724 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_82_clk
timestamp 1632082664
transform 1 0 47564 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_50_501
timestamp 1632082664
transform 1 0 47196 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1632082664
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_533
timestamp 1632082664
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1632082664
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1632082664
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1944_
timestamp 1632082664
transform 1 0 51704 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_50_549
timestamp 1632082664
transform 1 0 51612 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_545
timestamp 1632082664
transform 1 0 51244 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_578
timestamp 1632082664
transform 1 0 54280 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_566
timestamp 1632082664
transform 1 0 53176 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_586
timestamp 1632082664
transform 1 0 55016 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1948_
timestamp 1632082664
transform 1 0 55292 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1632082664
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1952_
timestamp 1632082664
transform 1 0 57132 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_50_625
timestamp 1632082664
transform 1 0 58604 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_605
timestamp 1632082664
transform 1 0 56764 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_629
timestamp 1632082664
transform 1 0 58972 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1632082664
transform -1 0 59340 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0103_
timestamp 1632082664
transform 1 0 2576 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1632082664
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_15
timestamp 1632082664
transform 1 0 2484 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1632082664
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0100_
timestamp 1632082664
transform 1 0 4416 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_51_32
timestamp 1632082664
transform 1 0 4048 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1632082664
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1632082664
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_52
timestamp 1632082664
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0092_
timestamp 1632082664
transform 1 0 7728 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_51_69
timestamp 1632082664
transform 1 0 7452 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0087_
timestamp 1632082664
transform 1 0 9568 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_51_88
timestamp 1632082664
transform 1 0 9200 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0083_
timestamp 1632082664
transform 1 0 11500 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1632082664
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_108
timestamp 1632082664
transform 1 0 11040 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1142_
timestamp 1632082664
transform 1 0 14076 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_51_129
timestamp 1632082664
transform 1 0 12972 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_157
timestamp 1632082664
transform 1 0 15548 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_165
timestamp 1632082664
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0062_
timestamp 1632082664
transform 1 0 18032 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1632082664
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1632082664
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_181
timestamp 1632082664
transform 1 0 17756 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0058_
timestamp 1632082664
transform 1 0 19872 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_51_200
timestamp 1632082664
transform 1 0 19504 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1632082664
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1632082664
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1632082664
transform 1 0 21344 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0050_
timestamp 1632082664
transform 1 0 23184 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_51_237
timestamp 1632082664
transform 1 0 22908 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0047_
timestamp 1632082664
transform 1 0 25024 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_51_256
timestamp 1632082664
transform 1 0 24656 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1632082664
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1632082664
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_276
timestamp 1632082664
transform 1 0 26496 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0036_
timestamp 1632082664
transform 1 0 28336 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_51_312
timestamp 1632082664
transform 1 0 29808 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_293
timestamp 1632082664
transform 1 0 28060 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0034_
timestamp 1632082664
transform 1 0 30176 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1632082664
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_353
timestamp 1632082664
transform 1 0 33580 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0030_
timestamp 1632082664
transform 1 0 32108 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1632082664
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_76_clk
timestamp 1632082664
transform 1 0 34224 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_51_359
timestamp 1632082664
transform 1 0 34132 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_380
timestamp 1632082664
transform 1 0 36064 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1632082664
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_393
timestamp 1632082664
transform 1 0 37260 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0007_
timestamp 1632082664
transform 1 0 37720 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_51_397
timestamp 1632082664
transform 1 0 37628 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_414
timestamp 1632082664
transform 1 0 39192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0008_
timestamp 1632082664
transform 1 0 39560 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_51_434
timestamp 1632082664
transform 1 0 41032 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_446
timestamp 1632082664
transform 1 0 42136 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1632082664
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1632082664
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1981_
timestamp 1632082664
transform 1 0 43792 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_51_461
timestamp 1632082664
transform 1 0 43516 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1978_
timestamp 1632082664
transform 1 0 45632 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_51_500
timestamp 1632082664
transform 1 0 47104 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_480
timestamp 1632082664
transform 1 0 45264 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1972_
timestamp 1632082664
transform 1 0 48944 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_51_505
timestamp 1632082664
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1632082664
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_517
timestamp 1632082664
transform 1 0 48668 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1968_
timestamp 1632082664
transform 1 0 50784 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_51_536
timestamp 1632082664
transform 1 0 50416 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1945_
timestamp 1632082664
transform 1 0 52716 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1632082664
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_556
timestamp 1632082664
transform 1 0 52256 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_577
timestamp 1632082664
transform 1 0 54188 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1949_
timestamp 1632082664
transform 1 0 55292 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_51_605
timestamp 1632082664
transform 1 0 56764 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_617
timestamp 1632082664
transform 1 0 57868 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1632082664
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_613
timestamp 1632082664
transform 1 0 57500 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_629
timestamp 1632082664
transform 1 0 58972 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1632082664
transform -1 0 59340 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0104_
timestamp 1632082664
transform 1 0 2852 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1632082664
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1632082664
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1632082664
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_15
timestamp 1632082664
transform 1 0 2484 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1632082664
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1632082664
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0101_
timestamp 1632082664
transform 1 0 3864 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_53_35
timestamp 1632082664
transform 1 0 4324 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1632082664
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_29
timestamp 1632082664
transform 1 0 3772 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1632082664
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_47
timestamp 1632082664
transform 1 0 5428 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0095_
timestamp 1632082664
transform 1 0 6440 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1632082664
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_46
timestamp 1632082664
transform 1 0 5336 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1632082664
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1632082664
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_74
timestamp 1632082664
transform 1 0 7912 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1632082664
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1632082664
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1632082664
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0089_
timestamp 1632082664
transform 1 0 9292 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1632082664
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1632082664
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_85
timestamp 1632082664
transform 1 0 8924 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1632082664
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_117
timestamp 1632082664
transform 1 0 11868 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0128_
timestamp 1632082664
transform 1 0 12052 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0127_
timestamp 1632082664
transform 1 0 11500 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_52_105
timestamp 1632082664
transform 1 0 10764 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1632082664
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1632082664
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0134_
timestamp 1632082664
transform 1 0 14076 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0130_
timestamp 1632082664
transform 1 0 13340 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1632082664
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1632082664
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_129
timestamp 1632082664
transform 1 0 12972 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_135
timestamp 1632082664
transform 1 0 13524 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1632082664
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0137_
timestamp 1632082664
transform 1 0 15916 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1632082664
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_157
timestamp 1632082664
transform 1 0 15548 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0063_
timestamp 1632082664
transform 1 0 18032 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1632082664
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1632082664
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1632082664
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1632082664
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_181
timestamp 1632082664
transform 1 0 17756 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1632082664
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0059_
timestamp 1632082664
transform 1 0 19872 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1632082664
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1632082664
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1632082664
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_200
timestamp 1632082664
transform 1 0 19504 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0056_
timestamp 1632082664
transform 1 0 20608 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1632082664
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1632082664
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1632082664
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_228
timestamp 1632082664
transform 1 0 22080 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_209
timestamp 1632082664
transform 1 0 20332 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0051_
timestamp 1632082664
transform 1 0 22448 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0048_
timestamp 1632082664
transform 1 0 23184 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1632082664
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_237
timestamp 1632082664
transform 1 0 22908 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0046_
timestamp 1632082664
transform 1 0 25024 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0041_
timestamp 1632082664
transform 1 0 25760 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1632082664
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1632082664
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_256
timestamp 1632082664
transform 1 0 24656 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_265
timestamp 1632082664
transform 1 0 25484 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_281
timestamp 1632082664
transform 1 0 26956 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0038_
timestamp 1632082664
transform 1 0 27600 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1632082664
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1632082664
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_284
timestamp 1632082664
transform 1 0 27232 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_289
timestamp 1632082664
transform 1 0 27692 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1632082664
transform 1 0 29808 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _0037_
timestamp 1632082664
transform 1 0 27968 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1632082664
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1632082664
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_308
timestamp 1632082664
transform 1 0 29440 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1632082664
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0031_
timestamp 1632082664
transform 1 0 31096 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_52_325
timestamp 1632082664
transform 1 0 31004 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1632082664
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_321
timestamp 1632082664
transform 1 0 30636 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_354
timestamp 1632082664
transform 1 0 33672 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1995_
timestamp 1632082664
transform 1 0 33212 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1632082664
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_342
timestamp 1632082664
transform 1 0 32568 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1632082664
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_362
timestamp 1632082664
transform 1 0 34408 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0018_
timestamp 1632082664
transform 1 0 34684 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0016_
timestamp 1632082664
transform 1 0 35052 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1632082664
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_365
timestamp 1632082664
transform 1 0 34684 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1632082664
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_393
timestamp 1632082664
transform 1 0 37260 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_393
timestamp 1632082664
transform 1 0 37260 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_381
timestamp 1632082664
transform 1 0 36156 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1632082664
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1632082664
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0010_
timestamp 1632082664
transform 1 0 37904 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0009_
timestamp 1632082664
transform 1 0 38272 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_52_399
timestamp 1632082664
transform 1 0 37812 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_416
timestamp 1632082664
transform 1 0 39376 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_401
timestamp 1632082664
transform 1 0 37996 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_420
timestamp 1632082664
transform 1 0 39744 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1993_
timestamp 1632082664
transform 1 0 40480 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1991_
timestamp 1632082664
transform 1 0 41216 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1632082664
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1632082664
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_433
timestamp 1632082664
transform 1 0 40940 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_449
timestamp 1632082664
transform 1 0 42412 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1989_
timestamp 1632082664
transform 1 0 43056 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0298_
timestamp 1632082664
transform 1 0 42596 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1632082664
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_444
timestamp 1632082664
transform 1 0 41952 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_452
timestamp 1632082664
transform 1 0 42688 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_467
timestamp 1632082664
transform 1 0 44068 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1632082664
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1632082664
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_479
timestamp 1632082664
transform 1 0 45172 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_472
timestamp 1632082664
transform 1 0 44528 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1980_
timestamp 1632082664
transform 1 0 45632 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1977_
timestamp 1632082664
transform 1 0 46368 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_53_483
timestamp 1632082664
transform 1 0 45540 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_500
timestamp 1632082664
transform 1 0 47104 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_489
timestamp 1632082664
transform 1 0 46092 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1974_
timestamp 1632082664
transform 1 0 48208 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1970_
timestamp 1632082664
transform 1 0 48944 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_53_505
timestamp 1632082664
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1632082664
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_508
timestamp 1632082664
transform 1 0 47840 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_517
timestamp 1632082664
transform 1 0 48668 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_533
timestamp 1632082664
transform 1 0 50140 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1969_
timestamp 1632082664
transform 1 0 50784 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1966_
timestamp 1632082664
transform 1 0 50876 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1632082664
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_536
timestamp 1632082664
transform 1 0 50416 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_528
timestamp 1632082664
transform 1 0 49680 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1947_
timestamp 1632082664
transform 1 0 52716 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_53_561
timestamp 1632082664
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1632082664
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_556
timestamp 1632082664
transform 1 0 52256 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_557
timestamp 1632082664
transform 1 0 52348 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_577
timestamp 1632082664
transform 1 0 54188 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1950_
timestamp 1632082664
transform 1 0 54188 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_53_573
timestamp 1632082664
transform 1 0 53820 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1951_
timestamp 1632082664
transform 1 0 55292 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_53_593
timestamp 1632082664
transform 1 0 55660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1632082664
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_585
timestamp 1632082664
transform 1 0 54924 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_605
timestamp 1632082664
transform 1 0 56764 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1955_
timestamp 1632082664
transform 1 0 57132 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_53_617
timestamp 1632082664
transform 1 0 57868 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1632082664
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_625
timestamp 1632082664
transform 1 0 58604 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_605
timestamp 1632082664
transform 1 0 56764 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_613
timestamp 1632082664
transform 1 0 57500 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_629
timestamp 1632082664
transform 1 0 58972 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_629
timestamp 1632082664
transform 1 0 58972 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1632082664
transform -1 0 59340 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1632082664
transform -1 0 59340 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1632082664
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1632082664
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1632082664
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0105_
timestamp 1632082664
transform 1 0 3772 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1632082664
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1632082664
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_57
timestamp 1632082664
transform 1 0 6348 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_45
timestamp 1632082664
transform 1 0 5244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_69
timestamp 1632082664
transform 1 0 7452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_81
timestamp 1632082664
transform 1 0 8556 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_97
timestamp 1632082664
transform 1 0 10028 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0125_
timestamp 1632082664
transform 1 0 10212 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1632082664
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1632082664
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0126_
timestamp 1632082664
transform 1 0 12052 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_54_115
timestamp 1632082664
transform 1 0 11684 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0133_
timestamp 1632082664
transform 1 0 14076 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1632082664
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1632082664
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_135
timestamp 1632082664
transform 1 0 13524 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0135_
timestamp 1632082664
transform 1 0 15916 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_54_157
timestamp 1632082664
transform 1 0 15548 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1632082664
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1632082664
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0060_
timestamp 1632082664
transform 1 0 19596 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1632082664
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1632082664
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_197
timestamp 1632082664
transform 1 0 19228 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_229
timestamp 1632082664
transform 1 0 22172 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_217
timestamp 1632082664
transform 1 0 21068 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0054_
timestamp 1632082664
transform 1 0 22356 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_54_247
timestamp 1632082664
transform 1 0 23828 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_265
timestamp 1632082664
transform 1 0 25484 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1632082664
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1632082664
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1632082664
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_14_clk
timestamp 1632082664
transform 1 0 26036 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_54_291
timestamp 1632082664
transform 1 0 27876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_309
timestamp 1632082664
transform 1 0 29532 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1632082664
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1632082664
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_303
timestamp 1632082664
transform 1 0 28980 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0035_
timestamp 1632082664
transform 1 0 30176 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_54_315
timestamp 1632082664
transform 1 0 30084 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_332
timestamp 1632082664
transform 1 0 31648 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_353
timestamp 1632082664
transform 1 0 33580 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0188_
timestamp 1632082664
transform 1 0 32108 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_54_336
timestamp 1632082664
transform 1 0 32016 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1632082664
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1632082664
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_361
timestamp 1632082664
transform 1 0 34316 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_394
timestamp 1632082664
transform 1 0 37352 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0015_
timestamp 1632082664
transform 1 0 35880 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_54_377
timestamp 1632082664
transform 1 0 35788 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0012_
timestamp 1632082664
transform 1 0 37904 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_54_416
timestamp 1632082664
transform 1 0 39376 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_421
timestamp 1632082664
transform 1 0 39836 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0228_
timestamp 1632082664
transform 1 0 40388 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1632082664
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0230_
timestamp 1632082664
transform 1 0 42228 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_54_443
timestamp 1632082664
transform 1 0 41860 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0240_
timestamp 1632082664
transform 1 0 44988 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_54_463
timestamp 1632082664
transform 1 0 43700 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1632082664
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1632082664
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_493
timestamp 1632082664
transform 1 0 46460 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_505
timestamp 1632082664
transform 1 0 47564 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1973_
timestamp 1632082664
transform 1 0 48208 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_54_511
timestamp 1632082664
transform 1 0 48116 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_533
timestamp 1632082664
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1632082664
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_528
timestamp 1632082664
transform 1 0 49680 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1964_
timestamp 1632082664
transform 1 0 51520 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_54_545
timestamp 1632082664
transform 1 0 51244 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1961_
timestamp 1632082664
transform 1 0 53360 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_54_564
timestamp 1632082664
transform 1 0 52992 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1956_
timestamp 1632082664
transform 1 0 56488 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_54_589
timestamp 1632082664
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1632082664
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_601
timestamp 1632082664
transform 1 0 56396 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_584
timestamp 1632082664
transform 1 0 54832 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_618
timestamp 1632082664
transform 1 0 57960 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1632082664
transform -1 0 59340 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_15
timestamp 1632082664
transform 1 0 2484 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1632082664
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1632082664
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0106_
timestamp 1632082664
transform 1 0 3312 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_55_40
timestamp 1632082664
transform 1 0 4784 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_23
timestamp 1632082664
transform 1 0 3220 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0114_
timestamp 1632082664
transform 1 0 6348 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1632082664
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1632082664
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0117_
timestamp 1632082664
transform 1 0 8188 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_55_73
timestamp 1632082664
transform 1 0 7820 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1632082664
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1632082664
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_113
timestamp 1632082664
transform 1 0 11500 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0124_
timestamp 1632082664
transform 1 0 12236 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1632082664
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1632082664
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0129_
timestamp 1632082664
transform 1 0 14076 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_55_137
timestamp 1632082664
transform 1 0 13708 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_157
timestamp 1632082664
transform 1 0 15548 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_165
timestamp 1632082664
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0138_
timestamp 1632082664
transform 1 0 16652 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1632082664
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_185
timestamp 1632082664
transform 1 0 18124 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0140_
timestamp 1632082664
transform 1 0 18492 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1632082664
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1632082664
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_225
timestamp 1632082664
transform 1 0 21804 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1632082664
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1632082664
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0158_
timestamp 1632082664
transform 1 0 22540 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_55_249
timestamp 1632082664
transform 1 0 24012 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_269
timestamp 1632082664
transform 1 0 25852 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0160_
timestamp 1632082664
transform 1 0 24380 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_55_281
timestamp 1632082664
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_289
timestamp 1632082664
transform 1 0 27692 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0040_
timestamp 1632082664
transform 1 0 27876 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1632082664
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_277
timestamp 1632082664
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_307
timestamp 1632082664
transform 1 0 29348 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0182_
timestamp 1632082664
transform 1 0 30084 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_55_331
timestamp 1632082664
transform 1 0 31556 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_353
timestamp 1632082664
transform 1 0 33580 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0186_
timestamp 1632082664
transform 1 0 32108 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1632082664
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1632082664
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0017_
timestamp 1632082664
transform 1 0 34592 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_55_361
timestamp 1632082664
transform 1 0 34316 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0013_
timestamp 1632082664
transform 1 0 37260 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_55_380
timestamp 1632082664
transform 1 0 36064 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1632082664
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_409
timestamp 1632082664
transform 1 0 38732 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_437
timestamp 1632082664
transform 1 0 41308 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0227_
timestamp 1632082664
transform 1 0 39836 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0232_
timestamp 1632082664
transform 1 0 42412 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1632082664
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_445
timestamp 1632082664
transform 1 0 42044 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0238_
timestamp 1632082664
transform 1 0 44252 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_55_465
timestamp 1632082664
transform 1 0 43884 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1632082664
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1632082664
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0243_
timestamp 1632082664
transform 1 0 47564 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1632082664
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1632082664
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_533
timestamp 1632082664
transform 1 0 50140 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1967_
timestamp 1632082664
transform 1 0 50784 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_55_521
timestamp 1632082664
transform 1 0 49036 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_539
timestamp 1632082664
transform 1 0 50692 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_561
timestamp 1632082664
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1632082664
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_556
timestamp 1632082664
transform 1 0 52256 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1960_
timestamp 1632082664
transform 1 0 54096 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_55_573
timestamp 1632082664
transform 1 0 53820 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1957_
timestamp 1632082664
transform 1 0 55936 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_55_592
timestamp 1632082664
transform 1 0 55568 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_617
timestamp 1632082664
transform 1 0 57868 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1632082664
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_612
timestamp 1632082664
transform 1 0 57408 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_629
timestamp 1632082664
transform 1 0 58972 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1632082664
transform -1 0 59340 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1632082664
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1632082664
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1632082664
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0107_
timestamp 1632082664
transform 1 0 3772 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1632082664
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1632082664
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0109_
timestamp 1632082664
transform 1 0 5612 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_56_45
timestamp 1632082664
transform 1 0 5244 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1632082664
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1632082664
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1632082664
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0118_
timestamp 1632082664
transform 1 0 8924 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1632082664
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_101
timestamp 1632082664
transform 1 0 10396 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0122_
timestamp 1632082664
transform 1 0 10764 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1632082664
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1632082664
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_56_141
timestamp 1632082664
transform 1 0 14076 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1632082664
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1632082664
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0136_
timestamp 1632082664
transform 1 0 14812 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_56_165
timestamp 1632082664
transform 1 0 16284 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_185
timestamp 1632082664
transform 1 0 18124 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0139_
timestamp 1632082664
transform 1 0 16652 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0153_
timestamp 1632082664
transform 1 0 19596 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1632082664
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_197
timestamp 1632082664
transform 1 0 19228 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_193
timestamp 1632082664
transform 1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0156_
timestamp 1632082664
transform 1 0 21436 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_56_217
timestamp 1632082664
transform 1 0 21068 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_237
timestamp 1632082664
transform 1 0 22908 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_249
timestamp 1632082664
transform 1 0 24012 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0164_
timestamp 1632082664
transform 1 0 24380 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_56_269
timestamp 1632082664
transform 1 0 25852 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1632082664
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0043_
timestamp 1632082664
transform 1 0 26956 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_56_297
timestamp 1632082664
transform 1 0 28428 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1632082664
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_309
timestamp 1632082664
transform 1 0 29532 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_305
timestamp 1632082664
transform 1 0 29164 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_329
timestamp 1632082664
transform 1 0 31372 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0181_
timestamp 1632082664
transform 1 0 29900 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0185_
timestamp 1632082664
transform 1 0 31924 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_56_351
timestamp 1632082664
transform 1 0 33396 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1996_
timestamp 1632082664
transform 1 0 34776 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1632082664
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_365
timestamp 1632082664
transform 1 0 34684 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1632082664
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0014_
timestamp 1632082664
transform 1 0 36616 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_56_382
timestamp 1632082664
transform 1 0 36248 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_414
timestamp 1632082664
transform 1 0 39192 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_402
timestamp 1632082664
transform 1 0 38088 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0226_
timestamp 1632082664
transform 1 0 40296 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1632082664
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_425
timestamp 1632082664
transform 1 0 40204 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_421
timestamp 1632082664
transform 1 0 39836 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0229_
timestamp 1632082664
transform 1 0 42136 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_56_442
timestamp 1632082664
transform 1 0 41768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_474
timestamp 1632082664
transform 1 0 44712 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0236_
timestamp 1632082664
transform 1 0 44988 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_56_462
timestamp 1632082664
transform 1 0 43608 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1632082664
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0241_
timestamp 1632082664
transform 1 0 46828 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_56_493
timestamp 1632082664
transform 1 0 46460 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_513
timestamp 1632082664
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1632082664
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_56_533
timestamp 1632082664
transform 1 0 50140 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0251_
timestamp 1632082664
transform 1 0 50876 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1632082664
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1632082664
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_557
timestamp 1632082664
transform 1 0 52348 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1963_
timestamp 1632082664
transform 1 0 53360 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_56_565
timestamp 1632082664
transform 1 0 53084 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0260_
timestamp 1632082664
transform 1 0 55292 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1632082664
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_584
timestamp 1632082664
transform 1 0 54832 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1958_
timestamp 1632082664
transform 1 0 57132 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_56_625
timestamp 1632082664
transform 1 0 58604 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_605
timestamp 1632082664
transform 1 0 56764 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_629
timestamp 1632082664
transform 1 0 58972 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1632082664
transform -1 0 59340 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1632082664
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1632082664
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1632082664
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0108_
timestamp 1632082664
transform 1 0 4048 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_57_31
timestamp 1632082664
transform 1 0 3956 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_27
timestamp 1632082664
transform 1 0 3588 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_48
timestamp 1632082664
transform 1 0 5520 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0112_
timestamp 1632082664
transform 1 0 6348 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1632082664
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0115_
timestamp 1632082664
transform 1 0 8188 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_57_73
timestamp 1632082664
transform 1 0 7820 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1632082664
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_20_clk
timestamp 1632082664
transform 1 0 11868 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1632082664
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1632082664
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1632082664
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_113
timestamp 1632082664
transform 1 0 11500 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0131_
timestamp 1632082664
transform 1 0 14076 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_57_137
timestamp 1632082664
transform 1 0 13708 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_157
timestamp 1632082664
transform 1 0 15548 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_165
timestamp 1632082664
transform 1 0 16284 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0141_
timestamp 1632082664
transform 1 0 17020 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1632082664
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_169
timestamp 1632082664
transform 1 0 16652 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_189
timestamp 1632082664
transform 1 0 18492 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0151_
timestamp 1632082664
transform 1 0 19228 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_57_213
timestamp 1632082664
transform 1 0 20700 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0155_
timestamp 1632082664
transform 1 0 21804 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1632082664
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_221
timestamp 1632082664
transform 1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0162_
timestamp 1632082664
transform 1 0 23644 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_57_241
timestamp 1632082664
transform 1 0 23276 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_261
timestamp 1632082664
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1632082664
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0168_
timestamp 1632082664
transform 1 0 26956 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1632082664
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1632082664
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0180_
timestamp 1632082664
transform 1 0 29808 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_57_297
timestamp 1632082664
transform 1 0 28428 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_309
timestamp 1632082664
transform 1 0 29532 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_328
timestamp 1632082664
transform 1 0 31280 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0183_
timestamp 1632082664
transform 1 0 32108 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1632082664
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_353
timestamp 1632082664
transform 1 0 33580 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0189_
timestamp 1632082664
transform 1 0 33948 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1632082664
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1632082664
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_393
timestamp 1632082664
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1632082664
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1632082664
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0224_
timestamp 1632082664
transform 1 0 38272 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_57_401
timestamp 1632082664
transform 1 0 37996 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_74_clk
timestamp 1632082664
transform 1 0 40112 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_57_420
timestamp 1632082664
transform 1 0 39744 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0233_
timestamp 1632082664
transform 1 0 42412 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1632082664
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_444
timestamp 1632082664
transform 1 0 41952 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0235_
timestamp 1632082664
transform 1 0 44252 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_57_465
timestamp 1632082664
transform 1 0 43884 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1632082664
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1632082664
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0245_
timestamp 1632082664
transform 1 0 47564 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1632082664
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1632082664
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0248_
timestamp 1632082664
transform 1 0 49404 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_57_541
timestamp 1632082664
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_521
timestamp 1632082664
transform 1 0 49036 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1632082664
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0257_
timestamp 1632082664
transform 1 0 52716 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1632082664
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1632082664
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_68_clk
timestamp 1632082664
transform 1 0 54740 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_57_577
timestamp 1632082664
transform 1 0 54188 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_603
timestamp 1632082664
transform 1 0 56580 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_617
timestamp 1632082664
transform 1 0 57868 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1632082664
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1632082664
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_629
timestamp 1632082664
transform 1 0 58972 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1632082664
transform -1 0 59340 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1632082664
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1632082664
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1632082664
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0111_
timestamp 1632082664
transform 1 0 4876 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1632082664
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1632082664
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1632082664
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0113_
timestamp 1632082664
transform 1 0 6716 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_58_57
timestamp 1632082664
transform 1 0 6348 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1632082664
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1632082664
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0119_
timestamp 1632082664
transform 1 0 8924 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1632082664
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_101
timestamp 1632082664
transform 1 0 10396 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0123_
timestamp 1632082664
transform 1 0 10764 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1632082664
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1632082664
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1140_
timestamp 1632082664
transform 1 0 14076 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1632082664
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1632082664
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_157
timestamp 1632082664
transform 1 0 15548 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0142_
timestamp 1632082664
transform 1 0 17112 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_58_173
timestamp 1632082664
transform 1 0 17020 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_169
timestamp 1632082664
transform 1 0 16652 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_190
timestamp 1632082664
transform 1 0 18584 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0150_
timestamp 1632082664
transform 1 0 19228 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1632082664
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_15_clk
timestamp 1632082664
transform 1 0 21068 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_58_213
timestamp 1632082664
transform 1 0 20700 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_237
timestamp 1632082664
transform 1 0 22908 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_249
timestamp 1632082664
transform 1 0 24012 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0161_
timestamp 1632082664
transform 1 0 24380 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1632082664
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_269
timestamp 1632082664
transform 1 0 25852 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0166_
timestamp 1632082664
transform 1 0 26220 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1632082664
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1632082664
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0178_
timestamp 1632082664
transform 1 0 29532 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1632082664
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1632082664
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_325
timestamp 1632082664
transform 1 0 31004 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0184_
timestamp 1632082664
transform 1 0 31648 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_58_331
timestamp 1632082664
transform 1 0 31556 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_348
timestamp 1632082664
transform 1 0 33120 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0191_
timestamp 1632082664
transform 1 0 34684 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1632082664
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 1632082664
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_393
timestamp 1632082664
transform 1 0 37260 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_381
timestamp 1632082664
transform 1 0 36156 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0223_
timestamp 1632082664
transform 1 0 37904 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_58_399
timestamp 1632082664
transform 1 0 37812 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_416
timestamp 1632082664
transform 1 0 39376 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0225_
timestamp 1632082664
transform 1 0 39836 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_58_437
timestamp 1632082664
transform 1 0 41308 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1632082664
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0234_
timestamp 1632082664
transform 1 0 42504 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_58_449
timestamp 1632082664
transform 1 0 42412 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_466
timestamp 1632082664
transform 1 0 43976 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_474
timestamp 1632082664
transform 1 0 44712 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0239_
timestamp 1632082664
transform 1 0 44988 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1632082664
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0244_
timestamp 1632082664
transform 1 0 46828 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_58_493
timestamp 1632082664
transform 1 0 46460 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_513
timestamp 1632082664
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1632082664
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0249_
timestamp 1632082664
transform 1 0 50140 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1632082664
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1632082664
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0254_
timestamp 1632082664
transform 1 0 51980 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_58_549
timestamp 1632082664
transform 1 0 51612 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1632082664
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_569
timestamp 1632082664
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0263_
timestamp 1632082664
transform 1 0 55292 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1632082664
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1632082664
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1959_
timestamp 1632082664
transform 1 0 57132 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_58_625
timestamp 1632082664
transform 1 0 58604 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_605
timestamp 1632082664
transform 1 0 56764 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_629
timestamp 1632082664
transform 1 0 58972 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1632082664
transform -1 0 59340 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1632082664
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1632082664
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1632082664
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1632082664
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1632082664
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1632082664
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1632082664
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1632082664
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1632082664
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1632082664
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1632082664
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1632082664
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_21_clk
timestamp 1632082664
transform 1 0 6716 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_60_53
timestamp 1632082664
transform 1 0 5980 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_61
timestamp 1632082664
transform 1 0 6716 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1632082664
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1632082664
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_57
timestamp 1632082664
transform 1 0 6348 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1632082664
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0116_
timestamp 1632082664
transform 1 0 6900 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1632082664
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_79
timestamp 1632082664
transform 1 0 8372 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_81
timestamp 1632082664
transform 1 0 8556 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_101
timestamp 1632082664
transform 1 0 10396 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0120_
timestamp 1632082664
transform 1 0 8924 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1632082664
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1632082664
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1632082664
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1136_
timestamp 1632082664
transform 1 0 11500 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1134_
timestamp 1632082664
transform 1 0 11500 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1632082664
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_109
timestamp 1632082664
transform 1 0 11132 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_109
timestamp 1632082664
transform 1 0 11132 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_129
timestamp 1632082664
transform 1 0 12972 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1139_
timestamp 1632082664
transform 1 0 14076 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1138_
timestamp 1632082664
transform 1 0 13340 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1632082664
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_129
timestamp 1632082664
transform 1 0 12972 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_137
timestamp 1632082664
transform 1 0 13708 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1632082664
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_157
timestamp 1632082664
transform 1 0 15548 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0145_
timestamp 1632082664
transform 1 0 16376 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1632082664
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_165
timestamp 1632082664
transform 1 0 16284 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_187
timestamp 1632082664
transform 1 0 18308 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_169
timestamp 1632082664
transform 1 0 16652 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0144_
timestamp 1632082664
transform 1 0 16836 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_60_182
timestamp 1632082664
transform 1 0 17848 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1632082664
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1632082664
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1632082664
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_195
timestamp 1632082664
transform 1 0 19044 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0149_
timestamp 1632082664
transform 1 0 19228 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0148_
timestamp 1632082664
transform 1 0 19228 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1632082664
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_213
timestamp 1632082664
transform 1 0 20700 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0159_
timestamp 1632082664
transform 1 0 21804 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0157_
timestamp 1632082664
transform 1 0 21068 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1632082664
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_213
timestamp 1632082664
transform 1 0 20700 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_221
timestamp 1632082664
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1632082664
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0163_
timestamp 1632082664
transform 1 0 23736 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1632082664
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_245
timestamp 1632082664
transform 1 0 23644 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_241
timestamp 1632082664
transform 1 0 23276 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_253
timestamp 1632082664
transform 1 0 24380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0167_
timestamp 1632082664
transform 1 0 25208 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_59_262
timestamp 1632082664
transform 1 0 25208 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1632082664
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_261
timestamp 1632082664
transform 1 0 25116 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1632082664
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_274
timestamp 1632082664
transform 1 0 26312 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0170_
timestamp 1632082664
transform 1 0 27048 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0169_
timestamp 1632082664
transform 1 0 26956 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1632082664
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_278
timestamp 1632082664
transform 1 0 26680 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_298
timestamp 1632082664
transform 1 0 28520 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_306
timestamp 1632082664
transform 1 0 29256 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0174_
timestamp 1632082664
transform 1 0 29624 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0172_
timestamp 1632082664
transform 1 0 28796 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1632082664
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_309
timestamp 1632082664
transform 1 0 29532 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_297
timestamp 1632082664
transform 1 0 28428 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1632082664
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0179_
timestamp 1632082664
transform 1 0 31464 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1632082664
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_326
timestamp 1632082664
transform 1 0 31096 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_337
timestamp 1632082664
transform 1 0 32108 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0190_
timestamp 1632082664
transform 1 0 33120 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_60_346
timestamp 1632082664
transform 1 0 32936 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1632082664
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1632082664
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_345
timestamp 1632082664
transform 1 0 32844 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_358
timestamp 1632082664
transform 1 0 34040 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0192_
timestamp 1632082664
transform 1 0 34960 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1632082664
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1632082664
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_364
timestamp 1632082664
transform 1 0 34592 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_75_clk
timestamp 1632082664
transform 1 0 35972 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_59_384
timestamp 1632082664
transform 1 0 36432 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_377
timestamp 1632082664
transform 1 0 35788 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0195_
timestamp 1632082664
transform 1 0 37260 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1632082664
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_411
timestamp 1632082664
transform 1 0 38916 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0222_
timestamp 1632082664
transform 1 0 39100 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_60_399
timestamp 1632082664
transform 1 0 37812 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_409
timestamp 1632082664
transform 1 0 38732 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_421
timestamp 1632082664
transform 1 0 39836 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0221_
timestamp 1632082664
transform 1 0 40388 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1632082664
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1632082664
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1632082664
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1632082664
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0294_
timestamp 1632082664
transform 1 0 43056 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_60_443
timestamp 1632082664
transform 1 0 41860 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1632082664
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1632082664
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_455
timestamp 1632082664
transform 1 0 42964 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1632082664
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_477
timestamp 1632082664
transform 1 0 44988 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0237_
timestamp 1632082664
transform 1 0 43608 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1632082664
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_461
timestamp 1632082664
transform 1 0 43516 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_472
timestamp 1632082664
transform 1 0 44528 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_478
timestamp 1632082664
transform 1 0 45080 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_500
timestamp 1632082664
transform 1 0 47104 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_498
timestamp 1632082664
transform 1 0 46920 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0293_
timestamp 1632082664
transform 1 0 45448 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0290_
timestamp 1632082664
transform 1 0 45632 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_60_483
timestamp 1632082664
transform 1 0 45540 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0247_
timestamp 1632082664
transform 1 0 47656 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0246_
timestamp 1632082664
transform 1 0 47564 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1632082664
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_69_clk
timestamp 1632082664
transform 1 0 49496 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_60_522
timestamp 1632082664
transform 1 0 49128 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_530
timestamp 1632082664
transform 1 0 49864 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0252_
timestamp 1632082664
transform 1 0 50140 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1632082664
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_525
timestamp 1632082664
transform 1 0 49404 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_521
timestamp 1632082664
transform 1 0 49036 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_558
timestamp 1632082664
transform 1 0 52440 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0256_
timestamp 1632082664
transform 1 0 51980 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0255_
timestamp 1632082664
transform 1 0 52716 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_59_546
timestamp 1632082664
transform 1 0 51336 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1632082664
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_549
timestamp 1632082664
transform 1 0 51612 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1632082664
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0259_
timestamp 1632082664
transform 1 0 54556 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_60_569
timestamp 1632082664
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_577
timestamp 1632082664
transform 1 0 54188 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0262_
timestamp 1632082664
transform 1 0 55292 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_59_597
timestamp 1632082664
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1632082664
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1632082664
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1632082664
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1962_
timestamp 1632082664
transform 1 0 57132 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_59_617
timestamp 1632082664
transform 1 0 57868 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1632082664
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1632082664
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_625
timestamp 1632082664
transform 1 0 58604 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_605
timestamp 1632082664
transform 1 0 56764 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_629
timestamp 1632082664
transform 1 0 58972 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_629
timestamp 1632082664
transform 1 0 58972 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1632082664
transform -1 0 59340 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1632082664
transform -1 0 59340 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1632082664
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1632082664
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1632082664
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_22_clk
timestamp 1632082664
transform 1 0 3956 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_61_27
timestamp 1632082664
transform 1 0 3588 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0743_
timestamp 1632082664
transform 1 0 6348 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1632082664
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1632082664
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1632082664
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_73
timestamp 1632082664
transform 1 0 7820 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_97
timestamp 1632082664
transform 1 0 10028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_85
timestamp 1632082664
transform 1 0 8924 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1132_
timestamp 1632082664
transform 1 0 11500 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1632082664
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_109
timestamp 1632082664
transform 1 0 11132 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1137_
timestamp 1632082664
transform 1 0 13340 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_61_129
timestamp 1632082664
transform 1 0 12972 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1632082664
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1632082664
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_16_clk
timestamp 1632082664
transform 1 0 18216 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1632082664
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1632082664
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_185
timestamp 1632082664
transform 1 0 18124 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1632082664
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_181
timestamp 1632082664
transform 1 0 17756 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_206
timestamp 1632082664
transform 1 0 20056 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_218
timestamp 1632082664
transform 1 0 21160 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1164_
timestamp 1632082664
transform 1 0 21804 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1632082664
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1165_
timestamp 1632082664
transform 1 0 23644 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_61_241
timestamp 1632082664
transform 1 0 23276 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1632082664
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1632082664
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0171_
timestamp 1632082664
transform 1 0 27048 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1632082664
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_281
timestamp 1632082664
transform 1 0 26956 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1632082664
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0173_
timestamp 1632082664
transform 1 0 28888 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_61_298
timestamp 1632082664
transform 1 0 28520 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_330
timestamp 1632082664
transform 1 0 31464 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_318
timestamp 1632082664
transform 1 0 30360 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0197_
timestamp 1632082664
transform 1 0 32108 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_61_353
timestamp 1632082664
transform 1 0 33580 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1632082664
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0193_
timestamp 1632082664
transform 1 0 34684 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 1632082664
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_381
timestamp 1632082664
transform 1 0 36156 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1632082664
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_389
timestamp 1632082664
transform 1 0 36892 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0214_
timestamp 1632082664
transform 1 0 37996 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0218_
timestamp 1632082664
transform 1 0 39928 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_61_421
timestamp 1632082664
transform 1 0 39836 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_417
timestamp 1632082664
transform 1 0 39468 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_438
timestamp 1632082664
transform 1 0 41400 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_446
timestamp 1632082664
transform 1 0 42136 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0219_
timestamp 1632082664
transform 1 0 42412 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1632082664
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_477
timestamp 1632082664
transform 1 0 44988 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_465
timestamp 1632082664
transform 1 0 43884 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0289_
timestamp 1632082664
transform 1 0 45632 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_61_483
timestamp 1632082664
transform 1 0 45540 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_500
timestamp 1632082664
transform 1 0 47104 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_505
timestamp 1632082664
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1632082664
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_517
timestamp 1632082664
transform 1 0 48668 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0250_
timestamp 1632082664
transform 1 0 49036 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_61_537
timestamp 1632082664
transform 1 0 50508 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_549
timestamp 1632082664
transform 1 0 51612 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0258_
timestamp 1632082664
transform 1 0 52716 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1632082664
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_557
timestamp 1632082664
transform 1 0 52348 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0261_
timestamp 1632082664
transform 1 0 54556 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_61_577
timestamp 1632082664
transform 1 0 54188 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_597
timestamp 1632082664
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1632082664
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_617
timestamp 1632082664
transform 1 0 57868 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1632082664
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1632082664
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_629
timestamp 1632082664
transform 1 0 58972 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1632082664
transform -1 0 59340 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1632082664
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1632082664
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1632082664
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1632082664
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1632082664
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1632082664
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1632082664
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_53
timestamp 1632082664
transform 1 0 5980 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0742_
timestamp 1632082664
transform 1 0 6532 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_62_75
timestamp 1632082664
transform 1 0 8004 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1632082664
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0740_
timestamp 1632082664
transform 1 0 8924 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_62_101
timestamp 1632082664
transform 1 0 10396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1632082664
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1131_
timestamp 1632082664
transform 1 0 11500 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_62_129
timestamp 1632082664
transform 1 0 12972 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1135_
timestamp 1632082664
transform 1 0 14076 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1632082664
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_137
timestamp 1632082664
transform 1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_157
timestamp 1632082664
transform 1 0 15548 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_185
timestamp 1632082664
transform 1 0 18124 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0146_
timestamp 1632082664
transform 1 0 16652 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0152_
timestamp 1632082664
transform 1 0 19228 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1632082664
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_193
timestamp 1632082664
transform 1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1161_
timestamp 1632082664
transform 1 0 21068 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_62_213
timestamp 1632082664
transform 1 0 20700 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1632082664
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1632082664
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1170_
timestamp 1632082664
transform 1 0 24380 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1632082664
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1632082664
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_269
timestamp 1632082664
transform 1 0 25852 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1171_
timestamp 1632082664
transform 1 0 26220 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1632082664
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1632082664
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0175_
timestamp 1632082664
transform 1 0 29532 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1632082664
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1632082664
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_325
timestamp 1632082664
transform 1 0 31004 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_45_clk
timestamp 1632082664
transform 1 0 32292 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_62_337
timestamp 1632082664
transform 1 0 32108 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_365
timestamp 1632082664
transform 1 0 34684 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0194_
timestamp 1632082664
transform 1 0 34868 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1632082664
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1632082664
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_359
timestamp 1632082664
transform 1 0 34132 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_383
timestamp 1632082664
transform 1 0 36340 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_391
timestamp 1632082664
transform 1 0 37076 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0212_
timestamp 1632082664
transform 1 0 37260 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_62_409
timestamp 1632082664
transform 1 0 38732 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0216_
timestamp 1632082664
transform 1 0 39836 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1632082664
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_437
timestamp 1632082664
transform 1 0 41308 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_417
timestamp 1632082664
transform 1 0 39468 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0217_
timestamp 1632082664
transform 1 0 41676 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1632082664
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1632082664
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1632082664
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1632082664
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1632082664
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_70_clk
timestamp 1632082664
transform 1 0 46460 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_62_489
timestamp 1632082664
transform 1 0 46092 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_513
timestamp 1632082664
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1632082664
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0284_
timestamp 1632082664
transform 1 0 50140 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1632082664
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1632082664
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1971_
timestamp 1632082664
transform 1 0 51980 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_62_549
timestamp 1632082664
transform 1 0 51612 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1632082664
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_569
timestamp 1632082664
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0265_
timestamp 1632082664
transform 1 0 55292 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1632082664
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1632082664
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_617
timestamp 1632082664
transform 1 0 57868 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_605
timestamp 1632082664
transform 1 0 56764 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_629
timestamp 1632082664
transform 1 0 58972 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1632082664
transform -1 0 59340 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1632082664
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1632082664
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1632082664
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_27
timestamp 1632082664
transform 1 0 3588 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0745_
timestamp 1632082664
transform 1 0 4416 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_63_35
timestamp 1632082664
transform 1 0 4324 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_57
timestamp 1632082664
transform 1 0 6348 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0741_
timestamp 1632082664
transform 1 0 6532 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1632082664
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1632082664
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0738_
timestamp 1632082664
transform 1 0 8372 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_63_75
timestamp 1632082664
transform 1 0 8004 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_95
timestamp 1632082664
transform 1 0 9844 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1130_
timestamp 1632082664
transform 1 0 11500 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1632082664
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1632082664
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_107
timestamp 1632082664
transform 1 0 10948 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_19_clk
timestamp 1632082664
transform 1 0 13524 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_63_129
timestamp 1632082664
transform 1 0 12972 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_155
timestamp 1632082664
transform 1 0 15364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_185
timestamp 1632082664
transform 1 0 18124 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0147_
timestamp 1632082664
transform 1 0 16652 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1632082664
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1632082664
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1158_
timestamp 1632082664
transform 1 0 18860 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1162_
timestamp 1632082664
transform 1 0 21804 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_209
timestamp 1632082664
transform 1 0 20332 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1632082664
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_221
timestamp 1632082664
transform 1 0 21436 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1167_
timestamp 1632082664
transform 1 0 23644 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_63_241
timestamp 1632082664
transform 1 0 23276 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_261
timestamp 1632082664
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_44_clk
timestamp 1632082664
transform 1 0 27324 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1632082664
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1632082664
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1632082664
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_281
timestamp 1632082664
transform 1 0 26956 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0177_
timestamp 1632082664
transform 1 0 29532 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_63_305
timestamp 1632082664
transform 1 0 29164 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_325
timestamp 1632082664
transform 1 0 31004 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_333
timestamp 1632082664
transform 1 0 31740 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0199_
timestamp 1632082664
transform 1 0 32108 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_353
timestamp 1632082664
transform 1 0 33580 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1632082664
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_365
timestamp 1632082664
transform 1 0 34684 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0196_
timestamp 1632082664
transform 1 0 35328 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_63_371
timestamp 1632082664
transform 1 0 35236 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0210_
timestamp 1632082664
transform 1 0 37260 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1632082664
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_388
timestamp 1632082664
transform 1 0 36800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0213_
timestamp 1632082664
transform 1 0 39100 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_63_409
timestamp 1632082664
transform 1 0 38732 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1632082664
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1632082664
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1632082664
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1632082664
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1632082664
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0292_
timestamp 1632082664
transform 1 0 43792 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_63_461
timestamp 1632082664
transform 1 0 43516 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0288_
timestamp 1632082664
transform 1 0 45632 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_63_500
timestamp 1632082664
transform 1 0 47104 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_480
timestamp 1632082664
transform 1 0 45264 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0282_
timestamp 1632082664
transform 1 0 48944 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_505
timestamp 1632082664
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1632082664
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_517
timestamp 1632082664
transform 1 0 48668 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0279_
timestamp 1632082664
transform 1 0 50784 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_63_536
timestamp 1632082664
transform 1 0 50416 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_561
timestamp 1632082664
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1632082664
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_556
timestamp 1632082664
transform 1 0 52256 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_573
timestamp 1632082664
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0266_
timestamp 1632082664
transform 1 0 55016 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_602
timestamp 1632082664
transform 1 0 56488 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_585
timestamp 1632082664
transform 1 0 54924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_614
timestamp 1632082664
transform 1 0 57592 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_617
timestamp 1632082664
transform 1 0 57868 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1632082664
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_629
timestamp 1632082664
transform 1 0 58972 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1632082664
transform -1 0 59340 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1632082664
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1632082664
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1632082664
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1632082664
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1632082664
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1632082664
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_41
timestamp 1632082664
transform 1 0 4876 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0744_
timestamp 1632082664
transform 1 0 5152 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_64_60
timestamp 1632082664
transform 1 0 6624 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0739_
timestamp 1632082664
transform 1 0 6992 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_64_80
timestamp 1632082664
transform 1 0 8464 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0736_
timestamp 1632082664
transform 1 0 8924 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_64_101
timestamp 1632082664
transform 1 0 10396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1632082664
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1129_
timestamp 1632082664
transform 1 0 11500 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_64_141
timestamp 1632082664
transform 1 0 14076 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_129
timestamp 1632082664
transform 1 0 12972 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1632082664
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1632082664
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1141_
timestamp 1632082664
transform 1 0 14812 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_64_165
timestamp 1632082664
transform 1 0 16284 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_185
timestamp 1632082664
transform 1 0 18124 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1146_
timestamp 1632082664
transform 1 0 16652 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1157_
timestamp 1632082664
transform 1 0 19228 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1632082664
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 1632082664
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1159_
timestamp 1632082664
transform 1 0 21068 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_64_213
timestamp 1632082664
transform 1 0 20700 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1632082664
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1632082664
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1169_
timestamp 1632082664
transform 1 0 24380 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1632082664
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1632082664
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_269
timestamp 1632082664
transform 1 0 25852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1173_
timestamp 1632082664
transform 1 0 26220 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_64_289
timestamp 1632082664
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1632082664
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1176_
timestamp 1632082664
transform 1 0 29532 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1632082664
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1632082664
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_325
timestamp 1632082664
transform 1 0 31004 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0200_
timestamp 1632082664
transform 1 0 31740 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_64_349
timestamp 1632082664
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0203_
timestamp 1632082664
transform 1 0 34684 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1632082664
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 1632082664
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0207_
timestamp 1632082664
transform 1 0 36524 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_64_381
timestamp 1632082664
transform 1 0 36156 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1632082664
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1632082664
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_73_clk
timestamp 1632082664
transform 1 0 41216 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1632082664
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1632082664
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1632082664
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_433
timestamp 1632082664
transform 1 0 40940 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_456
timestamp 1632082664
transform 1 0 43056 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_468
timestamp 1632082664
transform 1 0 44160 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1632082664
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1632082664
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0287_
timestamp 1632082664
transform 1 0 46368 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_64_489
timestamp 1632082664
transform 1 0 46092 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0283_
timestamp 1632082664
transform 1 0 48208 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_64_508
timestamp 1632082664
transform 1 0 47840 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_533
timestamp 1632082664
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1632082664
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_528
timestamp 1632082664
transform 1 0 49680 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0276_
timestamp 1632082664
transform 1 0 51520 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_64_545
timestamp 1632082664
transform 1 0 51244 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0272_
timestamp 1632082664
transform 1 0 53360 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_64_564
timestamp 1632082664
transform 1 0 52992 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0267_
timestamp 1632082664
transform 1 0 55292 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1632082664
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_584
timestamp 1632082664
transform 1 0 54832 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_617
timestamp 1632082664
transform 1 0 57868 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_605
timestamp 1632082664
transform 1 0 56764 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_629
timestamp 1632082664
transform 1 0 58972 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1632082664
transform -1 0 59340 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0750_
timestamp 1632082664
transform 1 0 2576 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1632082664
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_15
timestamp 1632082664
transform 1 0 2484 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1632082664
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0747_
timestamp 1632082664
transform 1 0 4416 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_65_32
timestamp 1632082664
transform 1 0 4048 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1632082664
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1632082664
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_52
timestamp 1632082664
transform 1 0 5888 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_69
timestamp 1632082664
transform 1 0 7452 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_77
timestamp 1632082664
transform 1 0 8188 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0735_
timestamp 1632082664
transform 1 0 8372 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_95
timestamp 1632082664
transform 1 0 9844 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1128_
timestamp 1632082664
transform 1 0 11776 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1632082664
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1632082664
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_107
timestamp 1632082664
transform 1 0 10948 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_65_113
timestamp 1632082664
transform 1 0 11500 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1143_
timestamp 1632082664
transform 1 0 14444 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_132
timestamp 1632082664
transform 1 0 13248 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_144
timestamp 1632082664
transform 1 0 14352 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1632082664
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1148_
timestamp 1632082664
transform 1 0 16652 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1632082664
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1632082664
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_185
timestamp 1632082664
transform 1 0 18124 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1156_
timestamp 1632082664
transform 1 0 18492 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_205
timestamp 1632082664
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1632082664
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1163_
timestamp 1632082664
transform 1 0 21804 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1632082664
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1632082664
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1168_
timestamp 1632082664
transform 1 0 23644 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_65_241
timestamp 1632082664
transform 1 0 23276 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_261
timestamp 1632082664
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _1180_ sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632082664
transform 1 0 27140 0 -1 38080
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1632082664
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_281
timestamp 1632082664
transform 1 0 26956 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1632082664
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1632082664
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1178_
timestamp 1632082664
transform 1 0 29072 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_65_300
timestamp 1632082664
transform 1 0 28704 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_320
timestamp 1632082664
transform 1 0 30544 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_332
timestamp 1632082664
transform 1 0 31648 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0201_
timestamp 1632082664
transform 1 0 32108 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1632082664
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_353
timestamp 1632082664
transform 1 0 33580 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0204_
timestamp 1632082664
transform 1 0 33948 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1632082664
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1632082664
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0211_
timestamp 1632082664
transform 1 0 37260 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1632082664
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1632082664
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0215_
timestamp 1632082664
transform 1 0 39100 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_65_409
timestamp 1632082664
transform 1 0 38732 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1632082664
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_449
timestamp 1632082664
transform 1 0 42412 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1632082664
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0295_
timestamp 1632082664
transform 1 0 43056 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1632082664
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_455
timestamp 1632082664
transform 1 0 42964 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1632082664
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_472
timestamp 1632082664
transform 1 0 44528 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0291_
timestamp 1632082664
transform 1 0 45540 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_65_499
timestamp 1632082664
transform 1 0 47012 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_65_480
timestamp 1632082664
transform 1 0 45264 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0281_
timestamp 1632082664
transform 1 0 48944 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_505
timestamp 1632082664
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1632082664
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1632082664
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_517
timestamp 1632082664
transform 1 0 48668 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0278_
timestamp 1632082664
transform 1 0 50784 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_65_536
timestamp 1632082664
transform 1 0 50416 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_561
timestamp 1632082664
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1632082664
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_556
timestamp 1632082664
transform 1 0 52256 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_67_clk
timestamp 1632082664
transform 1 0 54740 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_65_573
timestamp 1632082664
transform 1 0 53820 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_581
timestamp 1632082664
transform 1 0 54556 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_603
timestamp 1632082664
transform 1 0 56580 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_617
timestamp 1632082664
transform 1 0 57868 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1632082664
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1632082664
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_629
timestamp 1632082664
transform 1 0 58972 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1632082664
transform -1 0 59340 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1632082664
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1632082664
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1632082664
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1632082664
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1632082664
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1632082664
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_27
timestamp 1632082664
transform 1 0 3588 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0749_
timestamp 1632082664
transform 1 0 3772 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1632082664
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1632082664
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_41
timestamp 1632082664
transform 1 0 4876 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1632082664
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_57
timestamp 1632082664
transform 1 0 6348 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_67_45
timestamp 1632082664
transform 1 0 5244 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0746_
timestamp 1632082664
transform 1 0 4968 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_58
timestamp 1632082664
transform 1 0 6440 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1632082664
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp 1632082664
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_82
timestamp 1632082664
transform 1 0 8648 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0731_
timestamp 1632082664
transform 1 0 7084 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_70
timestamp 1632082664
transform 1 0 7544 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_81
timestamp 1632082664
transform 1 0 8556 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_101
timestamp 1632082664
transform 1 0 10396 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0734_
timestamp 1632082664
transform 1 0 8924 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0733_
timestamp 1632082664
transform 1 0 8924 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_101
timestamp 1632082664
transform 1 0 10396 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1632082664
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_113
timestamp 1632082664
transform 1 0 11500 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_66_113
timestamp 1632082664
transform 1 0 11500 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1127_
timestamp 1632082664
transform 1 0 12052 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1126_
timestamp 1632082664
transform 1 0 12144 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1632082664
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_119
timestamp 1632082664
transform 1 0 12052 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_109
timestamp 1632082664
transform 1 0 11132 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_66_141
timestamp 1632082664
transform 1 0 14076 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_136
timestamp 1632082664
transform 1 0 13616 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1632082664
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1632082664
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_135
timestamp 1632082664
transform 1 0 13524 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_160
timestamp 1632082664
transform 1 0 15824 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1145_
timestamp 1632082664
transform 1 0 14628 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_67_148
timestamp 1632082664
transform 1 0 14720 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_163
timestamp 1632082664
transform 1 0 16100 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1149_
timestamp 1632082664
transform 1 0 16928 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1147_
timestamp 1632082664
transform 1 0 16468 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_183
timestamp 1632082664
transform 1 0 17940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1632082664
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_169
timestamp 1632082664
transform 1 0 16652 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1154_
timestamp 1632082664
transform 1 0 19228 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1153_
timestamp 1632082664
transform 1 0 18768 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1632082664
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1632082664
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_208
timestamp 1632082664
transform 1 0 20240 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_188
timestamp 1632082664
transform 1 0 18400 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_clk
timestamp 1632082664
transform 1 0 20608 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_225
timestamp 1632082664
transform 1 0 21804 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_67_215
timestamp 1632082664
transform 1 0 20884 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1160_
timestamp 1632082664
transform 1 0 21068 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1632082664
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1632082664
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_213
timestamp 1632082664
transform 1 0 20700 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1632082664
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0357_
timestamp 1632082664
transform 1 0 22816 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1632082664
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_233
timestamp 1632082664
transform 1 0 22540 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1172_
timestamp 1632082664
transform 1 0 24380 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_67_264
timestamp 1632082664
transform 1 0 25392 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_252
timestamp 1632082664
transform 1 0 24288 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1632082664
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1632082664
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_269
timestamp 1632082664
transform 1 0 25852 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1181_
timestamp 1632082664
transform 1 0 26956 0 -1 39168
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1174_
timestamp 1632082664
transform 1 0 26220 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1632082664
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1632082664
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1632082664
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_310
timestamp 1632082664
transform 1 0 29624 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1632082664
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_309
timestamp 1632082664
transform 1 0 29532 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0337_
timestamp 1632082664
transform 1 0 29716 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_67_298
timestamp 1632082664
transform 1 0 28520 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1632082664
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1632082664
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0334_
timestamp 1632082664
transform 1 0 30176 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_327
timestamp 1632082664
transform 1 0 31188 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_332
timestamp 1632082664
transform 1 0 31648 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_337
timestamp 1632082664
transform 1 0 32108 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_339
timestamp 1632082664
transform 1 0 32292 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0325_
timestamp 1632082664
transform 1 0 32844 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0202_
timestamp 1632082664
transform 1 0 32476 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1632082664
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1632082664
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0206_
timestamp 1632082664
transform 1 0 34684 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0205_
timestamp 1632082664
transform 1 0 34684 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1632082664
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1632082664
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_361
timestamp 1632082664
transform 1 0 34316 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_381
timestamp 1632082664
transform 1 0 36156 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0208_
timestamp 1632082664
transform 1 0 36524 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1632082664
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1632082664
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_381
timestamp 1632082664
transform 1 0 36156 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_389
timestamp 1632082664
transform 1 0 36892 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1632082664
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0314_
timestamp 1632082664
transform 1 0 38824 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1632082664
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_409
timestamp 1632082664
transform 1 0 38732 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_405
timestamp 1632082664
transform 1 0 38364 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_426
timestamp 1632082664
transform 1 0 40296 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1632082664
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1632082664
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1632082664
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1632082664
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_438
timestamp 1632082664
transform 1 0 41400 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_66_445
timestamp 1632082664
transform 1 0 42044 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_446
timestamp 1632082664
transform 1 0 42136 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0299_
timestamp 1632082664
transform 1 0 42412 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0296_
timestamp 1632082664
transform 1 0 42872 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1632082664
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_453
timestamp 1632082664
transform 1 0 42780 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_470
timestamp 1632082664
transform 1 0 44344 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_465
timestamp 1632082664
transform 1 0 43884 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1632082664
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_477
timestamp 1632082664
transform 1 0 44988 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_477
timestamp 1632082664
transform 1 0 44988 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1632082664
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_66_498
timestamp 1632082664
transform 1 0 46920 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1632082664
transform 1 0 45448 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1632082664
transform 1 0 45356 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_66_481
timestamp 1632082664
transform 1 0 45356 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1632082664
transform 1 0 47932 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0285_
timestamp 1632082664
transform 1 0 47472 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_520
timestamp 1632082664
transform 1 0 48944 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1632082664
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1632082664
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_505
timestamp 1632082664
transform 1 0 47564 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_clk
timestamp 1632082664
transform 1 0 49772 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0280_
timestamp 1632082664
transform 1 0 50508 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_533
timestamp 1632082664
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1632082664
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_536
timestamp 1632082664
transform 1 0 50416 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_532
timestamp 1632082664
transform 1 0 50048 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_525
timestamp 1632082664
transform 1 0 49404 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1632082664
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_561
timestamp 1632082664
transform 1 0 52716 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0273_
timestamp 1632082664
transform 1 0 51520 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1632082664
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1632082664
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_545
timestamp 1632082664
transform 1 0 51244 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0271_
timestamp 1632082664
transform 1 0 53360 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0270_
timestamp 1632082664
transform 1 0 53452 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_66_564
timestamp 1632082664
transform 1 0 52992 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0269_
timestamp 1632082664
transform 1 0 55292 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0268_
timestamp 1632082664
transform 1 0 55292 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1632082664
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_585
timestamp 1632082664
transform 1 0 54924 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_584
timestamp 1632082664
transform 1 0 54832 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_605
timestamp 1632082664
transform 1 0 56764 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_617
timestamp 1632082664
transform 1 0 57868 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_617
timestamp 1632082664
transform 1 0 57868 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_605
timestamp 1632082664
transform 1 0 56764 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1632082664
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_613
timestamp 1632082664
transform 1 0 57500 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_67_629
timestamp 1632082664
transform 1 0 58972 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_629
timestamp 1632082664
transform 1 0 58972 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1632082664
transform -1 0 59340 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1632082664
transform -1 0 59340 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0753_
timestamp 1632082664
transform 1 0 1840 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_68_7
timestamp 1632082664
transform 1 0 1748 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_3
timestamp 1632082664
transform 1 0 1380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1632082664
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0751_
timestamp 1632082664
transform 1 0 3772 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1632082664
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_24
timestamp 1632082664
transform 1 0 3312 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0729_
timestamp 1632082664
transform 1 0 6348 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_68_45
timestamp 1632082664
transform 1 0 5244 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_73
timestamp 1632082664
transform 1 0 7820 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_81
timestamp 1632082664
transform 1 0 8556 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0732_
timestamp 1632082664
transform 1 0 8924 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_68_101
timestamp 1632082664
transform 1 0 10396 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1632082664
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_clk
timestamp 1632082664
transform 1 0 11500 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1125_
timestamp 1632082664
transform 1 0 12144 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_68_116
timestamp 1632082664
transform 1 0 11776 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1121_
timestamp 1632082664
transform 1 0 14168 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1632082664
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_141
timestamp 1632082664
transform 1 0 14076 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_136
timestamp 1632082664
transform 1 0 13616 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_158
timestamp 1632082664
transform 1 0 15640 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_166
timestamp 1632082664
transform 1 0 16376 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_185
timestamp 1632082664
transform 1 0 18124 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1150_
timestamp 1632082664
transform 1 0 16652 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1152_
timestamp 1632082664
transform 1 0 19228 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1632082664
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_193
timestamp 1632082664
transform 1 0 18860 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_68_225
timestamp 1632082664
transform 1 0 21804 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_213
timestamp 1632082664
transform 1 0 20700 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0356_
timestamp 1632082664
transform 1 0 22448 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_68_231
timestamp 1632082664
transform 1 0 22356 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_248
timestamp 1632082664
transform 1 0 23920 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1175_
timestamp 1632082664
transform 1 0 25760 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1632082664
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1632082664
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_265
timestamp 1632082664
transform 1 0 25484 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1179_
timestamp 1632082664
transform 1 0 27600 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_68_284
timestamp 1632082664
transform 1 0 27232 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1632082664
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1632082664
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_304
timestamp 1632082664
transform 1 0 29072 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0331_
timestamp 1632082664
transform 1 0 30912 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_68_321
timestamp 1632082664
transform 1 0 30636 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0328_
timestamp 1632082664
transform 1 0 32752 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_68_340
timestamp 1632082664
transform 1 0 32384 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1632082664
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1632082664
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_360
timestamp 1632082664
transform 1 0 34224 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0321_
timestamp 1632082664
transform 1 0 36064 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_68_377
timestamp 1632082664
transform 1 0 35788 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0317_
timestamp 1632082664
transform 1 0 37904 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_68_416
timestamp 1632082664
transform 1 0 39376 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_396
timestamp 1632082664
transform 1 0 37536 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_clk
timestamp 1632082664
transform 1 0 40296 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_429
timestamp 1632082664
transform 1 0 40572 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1632082664
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_425
timestamp 1632082664
transform 1 0 40204 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_421
timestamp 1632082664
transform 1 0 39836 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_441
timestamp 1632082664
transform 1 0 41676 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0300_
timestamp 1632082664
transform 1 0 42412 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_68_465
timestamp 1632082664
transform 1 0 43884 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1632082664
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1632082664
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_473
timestamp 1632082664
transform 1 0 44620 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1632082664
transform 1 0 46368 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_68_489
timestamp 1632082664
transform 1 0 46092 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1632082664
transform 1 0 48208 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_68_508
timestamp 1632082664
transform 1 0 47840 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_533
timestamp 1632082664
transform 1 0 50140 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0277_
timestamp 1632082664
transform 1 0 50876 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1632082664
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_528
timestamp 1632082664
transform 1 0 49680 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0274_
timestamp 1632082664
transform 1 0 52716 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_68_557
timestamp 1632082664
transform 1 0 52348 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_577
timestamp 1632082664
transform 1 0 54188 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_601
timestamp 1632082664
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_589
timestamp 1632082664
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1632082664
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_585
timestamp 1632082664
transform 1 0 54924 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_613
timestamp 1632082664
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_625
timestamp 1632082664
transform 1 0 58604 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_629
timestamp 1632082664
transform 1 0 58972 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1632082664
transform -1 0 59340 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_3
timestamp 1632082664
transform 1 0 1380 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0752_
timestamp 1632082664
transform 1 0 2208 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_69_11
timestamp 1632082664
transform 1 0 2116 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1632082664
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_23_clk
timestamp 1632082664
transform 1 0 4048 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_69_28
timestamp 1632082664
transform 1 0 3680 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0728_
timestamp 1632082664
transform 1 0 6348 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1632082664
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_52
timestamp 1632082664
transform 1 0 5888 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0730_
timestamp 1632082664
transform 1 0 8188 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_69_73
timestamp 1632082664
transform 1 0 7820 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1632082664
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_113
timestamp 1632082664
transform 1 0 11500 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1632082664
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1124_
timestamp 1632082664
transform 1 0 12144 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1632082664
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_119
timestamp 1632082664
transform 1 0 12052 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1632082664
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_136
timestamp 1632082664
transform 1 0 13616 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1120_
timestamp 1632082664
transform 1 0 14720 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_69_164
timestamp 1632082664
transform 1 0 16192 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1151_
timestamp 1632082664
transform 1 0 16652 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_69_185
timestamp 1632082664
transform 1 0 18124 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1632082664
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_197
timestamp 1632082664
transform 1 0 19228 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0358_
timestamp 1632082664
transform 1 0 19872 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_69_203
timestamp 1632082664
transform 1 0 19780 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1632082664
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1632082664
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_220
timestamp 1632082664
transform 1 0 21344 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0355_
timestamp 1632082664
transform 1 0 22908 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0349_
timestamp 1632082664
transform 1 0 24748 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_69_253
timestamp 1632082664
transform 1 0 24380 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1632082664
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1632082664
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1632082664
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1632082664
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0339_
timestamp 1632082664
transform 1 0 28336 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_69_312
timestamp 1632082664
transform 1 0 29808 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_69_293
timestamp 1632082664
transform 1 0 28060 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0335_
timestamp 1632082664
transform 1 0 30176 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_69_332
timestamp 1632082664
transform 1 0 31648 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_337
timestamp 1632082664
transform 1 0 32108 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0327_
timestamp 1632082664
transform 1 0 32752 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1632082664
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_343
timestamp 1632082664
transform 1 0 32660 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0322_
timestamp 1632082664
transform 1 0 35328 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_69_360
timestamp 1632082664
transform 1 0 34224 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1632082664
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_388
timestamp 1632082664
transform 1 0 36800 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_69_393
timestamp 1632082664
transform 1 0 37260 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0316_
timestamp 1632082664
transform 1 0 37536 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0311_
timestamp 1632082664
transform 1 0 39376 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_69_412
timestamp 1632082664
transform 1 0 39008 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_432
timestamp 1632082664
transform 1 0 40848 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0301_
timestamp 1632082664
transform 1 0 42412 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1632082664
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_444
timestamp 1632082664
transform 1 0 41952 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_477
timestamp 1632082664
transform 1 0 44988 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_465
timestamp 1632082664
transform 1 0 43884 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1632082664
transform 1 0 45632 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_69_483
timestamp 1632082664
transform 1 0 45540 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_500
timestamp 1632082664
transform 1 0 47104 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_71_clk
timestamp 1632082664
transform 1 0 47932 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1632082664
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_505
timestamp 1632082664
transform 1 0 47564 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1632082664
transform 1 0 50140 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_69_529
timestamp 1632082664
transform 1 0 49772 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_549
timestamp 1632082664
transform 1 0 51612 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_561
timestamp 1632082664
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1632082664
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_557
timestamp 1632082664
transform 1 0 52348 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_573
timestamp 1632082664
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_597
timestamp 1632082664
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_585
timestamp 1632082664
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1632082664
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_617
timestamp 1632082664
transform 1 0 57868 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1632082664
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1632082664
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_629
timestamp 1632082664
transform 1 0 58972 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1632082664
transform -1 0 59340 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0754_
timestamp 1632082664
transform 1 0 1840 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_70_7
timestamp 1632082664
transform 1 0 1748 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1632082664
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1632082664
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1632082664
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1632082664
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1632082664
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_24
timestamp 1632082664
transform 1 0 3312 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_53
timestamp 1632082664
transform 1 0 5980 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0727_
timestamp 1632082664
transform 1 0 6164 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_70_71
timestamp 1632082664
transform 1 0 7636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1632082664
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_85
timestamp 1632082664
transform 1 0 8924 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0719_
timestamp 1632082664
transform 1 0 9568 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1632082664
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_91
timestamp 1632082664
transform 1 0 9476 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0721_
timestamp 1632082664
transform 1 0 11408 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_70_108
timestamp 1632082664
transform 1 0 11040 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1632082664
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_128
timestamp 1632082664
transform 1 0 12880 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1632082664
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1119_
timestamp 1632082664
transform 1 0 15272 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_70_153
timestamp 1632082664
transform 1 0 15180 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_170
timestamp 1632082664
transform 1 0 16744 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1115_
timestamp 1632082664
transform 1 0 17296 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_17_clk
timestamp 1632082664
transform 1 0 19596 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1632082664
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_197
timestamp 1632082664
transform 1 0 19228 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_192
timestamp 1632082664
transform 1 0 18768 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_221
timestamp 1632082664
transform 1 0 21436 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_229
timestamp 1632082664
transform 1 0 22172 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0353_
timestamp 1632082664
transform 1 0 22448 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_70_248
timestamp 1632082664
transform 1 0 23920 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0347_
timestamp 1632082664
transform 1 0 25760 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1632082664
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1632082664
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_265
timestamp 1632082664
transform 1 0 25484 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0340_
timestamp 1632082664
transform 1 0 27600 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_70_284
timestamp 1632082664
transform 1 0 27232 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_309
timestamp 1632082664
transform 1 0 29532 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1632082664
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_304
timestamp 1632082664
transform 1 0 29072 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0333_
timestamp 1632082664
transform 1 0 30544 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_70_317
timestamp 1632082664
transform 1 0 30268 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_46_clk
timestamp 1632082664
transform 1 0 32384 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_70_336
timestamp 1632082664
transform 1 0 32016 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1632082664
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1632082664
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_360
timestamp 1632082664
transform 1 0 34224 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0320_
timestamp 1632082664
transform 1 0 36064 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_70_377
timestamp 1632082664
transform 1 0 35788 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0313_
timestamp 1632082664
transform 1 0 37904 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_70_416
timestamp 1632082664
transform 1 0 39376 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_396
timestamp 1632082664
transform 1 0 37536 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_421
timestamp 1632082664
transform 1 0 39836 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0309_
timestamp 1632082664
transform 1 0 40388 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1632082664
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_443
timestamp 1632082664
transform 1 0 41860 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0302_
timestamp 1632082664
transform 1 0 42412 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_70_465
timestamp 1632082664
transform 1 0 43884 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0306_
timestamp 1632082664
transform 1 0 44988 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1632082664
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_473
timestamp 1632082664
transform 1 0 44620 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_493
timestamp 1632082664
transform 1 0 46460 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_505
timestamp 1632082664
transform 1 0 47564 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1632082664
transform 1 0 48208 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_70_511
timestamp 1632082664
transform 1 0 48116 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1632082664
transform 1 0 50416 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1632082664
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_528
timestamp 1632082664
transform 1 0 49680 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_70_533
timestamp 1632082664
transform 1 0 50140 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 1632082664
transform 1 0 52256 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_70_552
timestamp 1632082664
transform 1 0 51888 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_572
timestamp 1632082664
transform 1 0 53728 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1632082664
transform 1 0 55292 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1632082664
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_584
timestamp 1632082664
transform 1 0 54832 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_617
timestamp 1632082664
transform 1 0 57868 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_605
timestamp 1632082664
transform 1 0 56764 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_629
timestamp 1632082664
transform 1 0 58972 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1632082664
transform -1 0 59340 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_3
timestamp 1632082664
transform 1 0 1380 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0755_
timestamp 1632082664
transform 1 0 2208 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_71_11
timestamp 1632082664
transform 1 0 2116 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1632082664
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0756_
timestamp 1632082664
transform 1 0 4048 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_71_28
timestamp 1632082664
transform 1 0 3680 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_48
timestamp 1632082664
transform 1 0 5520 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0725_
timestamp 1632082664
transform 1 0 6440 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1632082664
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_57
timestamp 1632082664
transform 1 0 6348 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_74
timestamp 1632082664
transform 1 0 7912 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_104
timestamp 1632082664
transform 1 0 10672 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_86
timestamp 1632082664
transform 1 0 9016 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0718_
timestamp 1632082664
transform 1 0 9200 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1632082664
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1632082664
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_125
timestamp 1632082664
transform 1 0 12604 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1123_
timestamp 1632082664
transform 1 0 12880 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_71_144
timestamp 1632082664
transform 1 0 14352 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1117_
timestamp 1632082664
transform 1 0 14720 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_71_164
timestamp 1632082664
transform 1 0 16192 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_169
timestamp 1632082664
transform 1 0 16652 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1114_
timestamp 1632082664
transform 1 0 17664 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1632082664
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_177
timestamp 1632082664
transform 1 0 17388 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_196
timestamp 1632082664
transform 1 0 19136 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0359_
timestamp 1632082664
transform 1 0 19872 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1632082664
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1632082664
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_220
timestamp 1632082664
transform 1 0 21344 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0351_
timestamp 1632082664
transform 1 0 23184 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_71_237
timestamp 1632082664
transform 1 0 22908 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0348_
timestamp 1632082664
transform 1 0 25024 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_71_256
timestamp 1632082664
transform 1 0 24656 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1632082664
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1632082664
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_276
timestamp 1632082664
transform 1 0 26496 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_293
timestamp 1632082664
transform 1 0 28060 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0342_
timestamp 1632082664
transform 1 0 28244 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_71_311
timestamp 1632082664
transform 1 0 29716 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0336_
timestamp 1632082664
transform 1 0 30176 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_71_315
timestamp 1632082664
transform 1 0 30084 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_332
timestamp 1632082664
transform 1 0 31648 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0329_
timestamp 1632082664
transform 1 0 32476 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1632082664
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_337
timestamp 1632082664
transform 1 0 32108 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0323_
timestamp 1632082664
transform 1 0 35328 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_71_357
timestamp 1632082664
transform 1 0 33948 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_369
timestamp 1632082664
transform 1 0 35052 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1632082664
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1632082664
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_388
timestamp 1632082664
transform 1 0 36800 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0312_
timestamp 1632082664
transform 1 0 38640 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_71_405
timestamp 1632082664
transform 1 0 38364 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0310_
timestamp 1632082664
transform 1 0 40480 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_71_424
timestamp 1632082664
transform 1 0 40112 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0303_
timestamp 1632082664
transform 1 0 42412 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1632082664
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_444
timestamp 1632082664
transform 1 0 41952 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_477
timestamp 1632082664
transform 1 0 44988 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 1632082664
transform 1 0 45172 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_71_465
timestamp 1632082664
transform 1 0 43884 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_495
timestamp 1632082664
transform 1 0 46644 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1632082664
transform 1 0 48944 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_71_505
timestamp 1632082664
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1632082664
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1632082664
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_517
timestamp 1632082664
transform 1 0 48668 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1632082664
transform 1 0 50784 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_71_536
timestamp 1632082664
transform 1 0 50416 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1632082664
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_556
timestamp 1632082664
transform 1 0 52256 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_71_561
timestamp 1632082664
transform 1 0 52716 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 1632082664
transform 1 0 52992 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_71_580
timestamp 1632082664
transform 1 0 54464 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1632082664
transform 1 0 55660 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_71_592
timestamp 1632082664
transform 1 0 55568 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1632082664
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_617
timestamp 1632082664
transform 1 0 57868 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1632082664
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1632082664
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_629
timestamp 1632082664
transform 1 0 58972 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1632082664
transform -1 0 59340 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0757_
timestamp 1632082664
transform 1 0 2852 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1632082664
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1632082664
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1632082664
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_15
timestamp 1632082664
transform 1 0 2484 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1632082664
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1632082664
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0758_
timestamp 1632082664
transform 1 0 3772 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_73_35
timestamp 1632082664
transform 1 0 4324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1632082664
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1632082664
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_57
timestamp 1632082664
transform 1 0 6348 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_73_57
timestamp 1632082664
transform 1 0 6348 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_47
timestamp 1632082664
transform 1 0 5428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_45
timestamp 1632082664
transform 1 0 5244 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1632082664
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1632082664
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_82
timestamp 1632082664
transform 1 0 8648 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0723_
timestamp 1632082664
transform 1 0 6992 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0722_
timestamp 1632082664
transform 1 0 7176 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_73_65
timestamp 1632082664
transform 1 0 7084 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_63
timestamp 1632082664
transform 1 0 6900 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_80
timestamp 1632082664
transform 1 0 8464 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_90
timestamp 1632082664
transform 1 0 9384 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_97
timestamp 1632082664
transform 1 0 10028 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0716_
timestamp 1632082664
transform 1 0 9568 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0714_
timestamp 1632082664
transform 1 0 10212 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1632082664
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1632082664
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0713_
timestamp 1632082664
transform 1 0 12052 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1632082664
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1632082664
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_108
timestamp 1632082664
transform 1 0 11040 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_115
timestamp 1632082664
transform 1 0 11684 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_73_125
timestamp 1632082664
transform 1 0 12604 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_18_clk
timestamp 1632082664
transform 1 0 14444 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _0711_
timestamp 1632082664
transform 1 0 12880 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1632082664
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1632082664
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_144
timestamp 1632082664
transform 1 0 14352 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_141
timestamp 1632082664
transform 1 0 14076 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_135
timestamp 1632082664
transform 1 0 13524 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_165
timestamp 1632082664
transform 1 0 16284 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1116_
timestamp 1632082664
transform 1 0 14720 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_73_164
timestamp 1632082664
transform 1 0 16192 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_169
timestamp 1632082664
transform 1 0 16652 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1113_
timestamp 1632082664
transform 1 0 17296 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1110_
timestamp 1632082664
transform 1 0 17388 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1632082664
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_72_173
timestamp 1632082664
transform 1 0 17020 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_193
timestamp 1632082664
transform 1 0 18860 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_72_197
timestamp 1632082664
transform 1 0 19228 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_205
timestamp 1632082664
transform 1 0 19964 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0361_
timestamp 1632082664
transform 1 0 19872 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0360_
timestamp 1632082664
transform 1 0 20148 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1632082664
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_192
timestamp 1632082664
transform 1 0 18768 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_73_201
timestamp 1632082664
transform 1 0 19596 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_225
timestamp 1632082664
transform 1 0 21804 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_72_223
timestamp 1632082664
transform 1 0 21620 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1632082664
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_220
timestamp 1632082664
transform 1 0 21344 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 1632082664
transform 1 0 22632 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0354_
timestamp 1632082664
transform 1 0 22448 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_73_233
timestamp 1632082664
transform 1 0 22540 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_231
timestamp 1632082664
transform 1 0 22356 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_250
timestamp 1632082664
transform 1 0 24104 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_248
timestamp 1632082664
transform 1 0 23920 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_270
timestamp 1632082664
transform 1 0 25944 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0350_
timestamp 1632082664
transform 1 0 24472 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0346_
timestamp 1632082664
transform 1 0 25760 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1632082664
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1632082664
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_72_265
timestamp 1632082664
transform 1 0 25484 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_281
timestamp 1632082664
transform 1 0 26956 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_278
timestamp 1632082664
transform 1 0 26680 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0344_
timestamp 1632082664
transform 1 0 27692 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0343_
timestamp 1632082664
transform 1 0 27600 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1632082664
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_284
timestamp 1632082664
transform 1 0 27232 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0338_
timestamp 1632082664
transform 1 0 29532 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1632082664
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1632082664
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_304
timestamp 1632082664
transform 1 0 29072 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1632082664
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1632082664
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_325
timestamp 1632082664
transform 1 0 31004 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_353
timestamp 1632082664
transform 1 0 33580 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0332_
timestamp 1632082664
transform 1 0 32108 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1632082664
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1632082664
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1632082664
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1632082664
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_365
timestamp 1632082664
transform 1 0 34684 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0326_
timestamp 1632082664
transform 1 0 34684 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0324_
timestamp 1632082664
transform 1 0 35328 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1632082664
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_371
timestamp 1632082664
transform 1 0 35236 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_361
timestamp 1632082664
transform 1 0 34316 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_72_361
timestamp 1632082664
transform 1 0 34316 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_381
timestamp 1632082664
transform 1 0 36156 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_72_388
timestamp 1632082664
transform 1 0 36800 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1632082664
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1632082664
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_73_389
timestamp 1632082664
transform 1 0 36892 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0318_
timestamp 1632082664
transform 1 0 37812 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0315_
timestamp 1632082664
transform 1 0 38732 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_73_405
timestamp 1632082664
transform 1 0 38364 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_415
timestamp 1632082664
transform 1 0 39284 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_72_396
timestamp 1632082664
transform 1 0 37536 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_72_421
timestamp 1632082664
transform 1 0 39836 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_73_437
timestamp 1632082664
transform 1 0 41308 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1632082664
transform 1 0 40480 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_73_425
timestamp 1632082664
transform 1 0 40204 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1632082664
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_427
timestamp 1632082664
transform 1 0 40388 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1632082664
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_72_clk
timestamp 1632082664
transform 1 0 43148 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_73_449
timestamp 1632082664
transform 1 0 42412 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0304_
timestamp 1632082664
transform 1 0 42412 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1632082664
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_448
timestamp 1632082664
transform 1 0 42320 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_444
timestamp 1632082664
transform 1 0 41952 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_73_445
timestamp 1632082664
transform 1 0 42044 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_72_465
timestamp 1632082664
transform 1 0 43884 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1632082664
transform 1 0 44988 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1632082664
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_477
timestamp 1632082664
transform 1 0 44988 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_72_473
timestamp 1632082664
transform 1 0 44620 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1632082664
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1632082664
transform 1 0 45356 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_72_493
timestamp 1632082664
transform 1 0 46460 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1632082664
transform 1 0 47656 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1632082664
transform 1 0 48944 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_73_505
timestamp 1632082664
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1632082664
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1632082664
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_505
timestamp 1632082664
transform 1 0 47564 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_73_517
timestamp 1632082664
transform 1 0 48668 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_72_522
timestamp 1632082664
transform 1 0 49128 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_530
timestamp 1632082664
transform 1 0 49864 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1632082664
transform 1 0 50784 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_72_533
timestamp 1632082664
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1632082664
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_536
timestamp 1632082664
transform 1 0 50416 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_561
timestamp 1632082664
transform 1 0 52716 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1632082664
transform 1 0 51520 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1632082664
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_556
timestamp 1632082664
transform 1 0 52256 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_72_545
timestamp 1632082664
transform 1 0 51244 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 1632082664
transform 1 0 53360 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1632082664
transform 1 0 53728 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_72_564
timestamp 1632082664
transform 1 0 52992 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_73_569
timestamp 1632082664
transform 1 0 53452 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_66_clk
timestamp 1632082664
transform 1 0 55568 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_72_589
timestamp 1632082664
transform 1 0 55292 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1632082664
transform 1 0 55936 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1632082664
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_595
timestamp 1632082664
transform 1 0 55844 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_588
timestamp 1632082664
transform 1 0 55200 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_584
timestamp 1632082664
transform 1 0 54832 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_624
timestamp 1632082664
transform 1 0 58512 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_617
timestamp 1632082664
transform 1 0 57868 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_612
timestamp 1632082664
transform 1 0 57408 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1632082664
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_612
timestamp 1632082664
transform 1 0 57408 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_629
timestamp 1632082664
transform 1 0 58972 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1632082664
transform -1 0 59340 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1632082664
transform -1 0 59340 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1632082664
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1632082664
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1632082664
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0760_
timestamp 1632082664
transform 1 0 3772 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1632082664
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1632082664
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_57
timestamp 1632082664
transform 1 0 6348 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_74_45
timestamp 1632082664
transform 1 0 5244 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0724_
timestamp 1632082664
transform 1 0 6992 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_74_63
timestamp 1632082664
transform 1 0 6900 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_80
timestamp 1632082664
transform 1 0 8464 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_25_clk
timestamp 1632082664
transform 1 0 10212 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_74_97
timestamp 1632082664
transform 1 0 10028 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1632082664
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1632082664
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_119
timestamp 1632082664
transform 1 0 12052 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_131
timestamp 1632082664
transform 1 0 13156 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1632082664
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1632082664
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1632082664
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1118_
timestamp 1632082664
transform 1 0 15456 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_74_153
timestamp 1632082664
transform 1 0 15180 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1109_
timestamp 1632082664
transform 1 0 17296 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_74_172
timestamp 1632082664
transform 1 0 16928 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1632082664
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1632082664
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_192
timestamp 1632082664
transform 1 0 18768 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0362_
timestamp 1632082664
transform 1 0 20424 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_74_209
timestamp 1632082664
transform 1 0 20332 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_226
timestamp 1632082664
transform 1 0 21896 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_246
timestamp 1632082664
transform 1 0 23736 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0364_
timestamp 1632082664
transform 1 0 22264 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1632082664
transform 1 0 24380 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_74_269
timestamp 1632082664
transform 1 0 25852 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1632082664
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_43_clk
timestamp 1632082664
transform 1 0 27232 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_74_281
timestamp 1632082664
transform 1 0 26956 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1632082664
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1632082664
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_304
timestamp 1632082664
transform 1 0 29072 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_321
timestamp 1632082664
transform 1 0 30636 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 1632082664
transform 1 0 30820 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1632082664
transform 1 0 32660 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_74_339
timestamp 1632082664
transform 1 0 32292 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_365
timestamp 1632082664
transform 1 0 34684 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1632082664
transform 1 0 35328 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1632082664
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_371
timestamp 1632082664
transform 1 0 35236 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1632082664
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_359
timestamp 1632082664
transform 1 0 34132 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_388
timestamp 1632082664
transform 1 0 36800 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1632082664
transform 1 0 37904 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_74_416
timestamp 1632082664
transform 1 0 39376 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_421
timestamp 1632082664
transform 1 0 39836 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1044_
timestamp 1632082664
transform 1 0 40480 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1632082664
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_427
timestamp 1632082664
transform 1 0 40388 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0305_
timestamp 1632082664
transform 1 0 42320 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_74_444
timestamp 1632082664
transform 1 0 41952 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 1632082664
transform 1 0 44988 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_74_464
timestamp 1632082664
transform 1 0 43792 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1632082664
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_493
timestamp 1632082664
transform 1 0 46460 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1037_
timestamp 1632082664
transform 1 0 47564 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_74_521
timestamp 1632082664
transform 1 0 49036 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1632082664
transform 1 0 50140 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1632082664
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_529
timestamp 1632082664
transform 1 0 49772 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_74_561
timestamp 1632082664
transform 1 0 52716 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_74_549
timestamp 1632082664
transform 1 0 51612 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 1632082664
transform 1 0 53360 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_74_567
timestamp 1632082664
transform 1 0 53268 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_589
timestamp 1632082664
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1632082664
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_601
timestamp 1632082664
transform 1 0 56396 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_584
timestamp 1632082664
transform 1 0 54832 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_621
timestamp 1632082664
transform 1 0 58236 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1632082664
transform 1 0 56764 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_74_629
timestamp 1632082664
transform 1 0 58972 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1632082664
transform -1 0 59340 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0767_
timestamp 1632082664
transform 1 0 1656 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1632082664
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_75_3
timestamp 1632082664
transform 1 0 1380 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_22
timestamp 1632082664
transform 1 0 3128 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0761_
timestamp 1632082664
transform 1 0 3956 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_75_30
timestamp 1632082664
transform 1 0 3864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_47
timestamp 1632082664
transform 1 0 5428 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0763_
timestamp 1632082664
transform 1 0 6348 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1632082664
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1632082664
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_73
timestamp 1632082664
transform 1 0 7820 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_85
timestamp 1632082664
transform 1 0 8924 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0717_
timestamp 1632082664
transform 1 0 9568 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_75_91
timestamp 1632082664
transform 1 0 9476 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0712_
timestamp 1632082664
transform 1 0 11592 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1632082664
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_113
timestamp 1632082664
transform 1 0 11500 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_108
timestamp 1632082664
transform 1 0 11040 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0709_
timestamp 1632082664
transform 1 0 13432 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_75_130
timestamp 1632082664
transform 1 0 13064 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_162
timestamp 1632082664
transform 1 0 16008 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_150
timestamp 1632082664
transform 1 0 14904 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_169
timestamp 1632082664
transform 1 0 16652 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1108_
timestamp 1632082664
transform 1 0 17204 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1632082664
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_191
timestamp 1632082664
transform 1 0 18676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1112_
timestamp 1632082664
transform 1 0 19228 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_75_213
timestamp 1632082664
transform 1 0 20700 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0365_
timestamp 1632082664
transform 1 0 21804 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1632082664
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_75_221
timestamp 1632082664
transform 1 0 21436 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_241
timestamp 1632082664
transform 1 0 23276 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_42_clk
timestamp 1632082664
transform 1 0 24472 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_75_253
timestamp 1632082664
transform 1 0 24380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_274
timestamp 1632082664
transform 1 0 26312 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0345_
timestamp 1632082664
transform 1 0 27232 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1632082664
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_75_281
timestamp 1632082664
transform 1 0 26956 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1632082664
transform 1 0 29072 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_75_300
timestamp 1632082664
transform 1 0 28704 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_320
timestamp 1632082664
transform 1 0 30544 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_332
timestamp 1632082664
transform 1 0 31648 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1632082664
transform 1 0 33488 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1632082664
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1632082664
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_75_349
timestamp 1632082664
transform 1 0 33212 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1632082664
transform 1 0 35328 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_75_368
timestamp 1632082664
transform 1 0 34960 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1632082664
transform 1 0 37352 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1632082664
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_393
timestamp 1632082664
transform 1 0 37260 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_388
timestamp 1632082664
transform 1 0 36800 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_48_clk
timestamp 1632082664
transform 1 0 39192 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_75_410
timestamp 1632082664
transform 1 0 38824 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_434
timestamp 1632082664
transform 1 0 41032 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_446
timestamp 1632082664
transform 1 0 42136 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0307_
timestamp 1632082664
transform 1 0 42412 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1632082664
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1033_
timestamp 1632082664
transform 1 0 45080 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_75_465
timestamp 1632082664
transform 1 0 43884 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_477
timestamp 1632082664
transform 1 0 44988 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_494
timestamp 1632082664
transform 1 0 46552 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_75_505
timestamp 1632082664
transform 1 0 47564 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_75_502
timestamp 1632082664
transform 1 0 47288 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0981_
timestamp 1632082664
transform 1 0 48208 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1632082664
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_511
timestamp 1632082664
transform 1 0 48116 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1632082664
transform 1 0 50048 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_75_528
timestamp 1632082664
transform 1 0 49680 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_548
timestamp 1632082664
transform 1 0 51520 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1632082664
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_561
timestamp 1632082664
transform 1 0 52716 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_65_clk
timestamp 1632082664
transform 1 0 53084 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_75_585
timestamp 1632082664
transform 1 0 54924 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1632082664
transform 1 0 55936 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_75_593
timestamp 1632082664
transform 1 0 55660 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_617
timestamp 1632082664
transform 1 0 57868 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1632082664
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_612
timestamp 1632082664
transform 1 0 57408 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_629
timestamp 1632082664
transform 1 0 58972 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1632082664
transform -1 0 59340 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0766_
timestamp 1632082664
transform 1 0 1840 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_76_7
timestamp 1632082664
transform 1 0 1748 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_3
timestamp 1632082664
transform 1 0 1380 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1632082664
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_76_41
timestamp 1632082664
transform 1 0 4876 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1632082664
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1632082664
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_24
timestamp 1632082664
transform 1 0 3312 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_24_clk
timestamp 1632082664
transform 1 0 5612 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_76_69
timestamp 1632082664
transform 1 0 7452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_81
timestamp 1632082664
transform 1 0 8556 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_76_85
timestamp 1632082664
transform 1 0 8924 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0720_
timestamp 1632082664
transform 1 0 9568 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1632082664
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_91
timestamp 1632082664
transform 1 0 9476 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0710_
timestamp 1632082664
transform 1 0 12144 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_76_108
timestamp 1632082664
transform 1 0 11040 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0708_
timestamp 1632082664
transform 1 0 14076 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1632082664
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_136
timestamp 1632082664
transform 1 0 13616 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_157
timestamp 1632082664
transform 1 0 15548 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1107_
timestamp 1632082664
transform 1 0 17112 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_76_173
timestamp 1632082664
transform 1 0 17020 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_169
timestamp 1632082664
transform 1 0 16652 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_41_clk
timestamp 1632082664
transform 1 0 20240 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_76_190
timestamp 1632082664
transform 1 0 18584 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_76_197
timestamp 1632082664
transform 1 0 19228 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1632082664
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_76_205
timestamp 1632082664
transform 1 0 19964 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_228
timestamp 1632082664
transform 1 0 22080 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0366_
timestamp 1632082664
transform 1 0 22448 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_76_248
timestamp 1632082664
transform 1 0 23920 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_265
timestamp 1632082664
transform 1 0 25484 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1632082664
transform 1 0 25668 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1632082664
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1632082664
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1632082664
transform 1 0 27508 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_76_283
timestamp 1632082664
transform 1 0 27140 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1632082664
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1632082664
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1632082664
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_303
timestamp 1632082664
transform 1 0 28980 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_321
timestamp 1632082664
transform 1 0 30636 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1632082664
transform 1 0 30820 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1632082664
transform 1 0 32752 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_76_343
timestamp 1632082664
transform 1 0 32660 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_339
timestamp 1632082664
transform 1 0 32292 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_47_clk
timestamp 1632082664
transform 1 0 35052 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1632082664
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_365
timestamp 1632082664
transform 1 0 34684 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_360
timestamp 1632082664
transform 1 0 34224 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_389
timestamp 1632082664
transform 1 0 36892 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1632082664
transform 1 0 37904 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_76_416
timestamp 1632082664
transform 1 0 39376 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_76_397
timestamp 1632082664
transform 1 0 37628 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1632082664
transform 1 0 41216 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1632082664
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1632082664
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_76_433
timestamp 1632082664
transform 1 0 40940 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1039_
timestamp 1632082664
transform 1 0 43056 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_76_452
timestamp 1632082664
transform 1 0 42688 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1632082664
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_472
timestamp 1632082664
transform 1 0 44528 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_76_477
timestamp 1632082664
transform 1 0 44988 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 1632082664
transform 1 0 45264 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_76_496
timestamp 1632082664
transform 1 0 46736 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_64_clk
timestamp 1632082664
transform 1 0 47840 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1632082664
transform 1 0 50140 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1632082664
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_528
timestamp 1632082664
transform 1 0 49680 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1632082664
transform 1 0 51980 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_76_549
timestamp 1632082664
transform 1 0 51612 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1632082664
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_569
timestamp 1632082664
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 1632082664
transform 1 0 56488 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_76_589
timestamp 1632082664
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1632082664
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_601
timestamp 1632082664
transform 1 0 56396 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1632082664
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_618
timestamp 1632082664
transform 1 0 57960 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1632082664
transform -1 0 59340 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0768_
timestamp 1632082664
transform 1 0 1656 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1632082664
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_77_3
timestamp 1632082664
transform 1 0 1380 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0762_
timestamp 1632082664
transform 1 0 4324 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_77_22
timestamp 1632082664
transform 1 0 3128 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_34
timestamp 1632082664
transform 1 0 4232 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0764_
timestamp 1632082664
transform 1 0 6348 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1632082664
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1632082664
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1632082664
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0789_
timestamp 1632082664
transform 1 0 8188 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_77_73
timestamp 1632082664
transform 1 0 7820 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1632082664
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1632082664
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0793_
timestamp 1632082664
transform 1 0 11500 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1632082664
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1632082664
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_129
timestamp 1632082664
transform 1 0 12972 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0707_
timestamp 1632082664
transform 1 0 13616 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_77_135
timestamp 1632082664
transform 1 0 13524 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_152
timestamp 1632082664
transform 1 0 15088 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_164
timestamp 1632082664
transform 1 0 16192 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1106_
timestamp 1632082664
transform 1 0 16928 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1632082664
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_169
timestamp 1632082664
transform 1 0 16652 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_200
timestamp 1632082664
transform 1 0 19504 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_188
timestamp 1632082664
transform 1 0 18400 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0367_
timestamp 1632082664
transform 1 0 21804 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_77_212
timestamp 1632082664
transform 1 0 20608 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1632082664
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_241
timestamp 1632082664
transform 1 0 23276 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_253
timestamp 1632082664
transform 1 0 24380 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1632082664
transform 1 0 25024 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_77_259
timestamp 1632082664
transform 1 0 24932 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1632082664
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1632082664
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_276
timestamp 1632082664
transform 1 0 26496 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1632082664
transform 1 0 28336 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_77_312
timestamp 1632082664
transform 1 0 29808 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_77_293
timestamp 1632082664
transform 1 0 28060 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1632082664
transform 1 0 30176 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_77_332
timestamp 1632082664
transform 1 0 31648 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1632082664
transform 1 0 33488 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1632082664
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1632082664
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_349
timestamp 1632082664
transform 1 0 33212 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1632082664
transform 1 0 35328 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_77_368
timestamp 1632082664
transform 1 0 34960 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1632082664
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1632082664
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_388
timestamp 1632082664
transform 1 0 36800 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1632082664
transform 1 0 38640 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_77_405
timestamp 1632082664
transform 1 0 38364 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1043_
timestamp 1632082664
transform 1 0 40480 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_77_424
timestamp 1632082664
transform 1 0 40112 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_449
timestamp 1632082664
transform 1 0 42412 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1040_
timestamp 1632082664
transform 1 0 43056 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1632082664
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_455
timestamp 1632082664
transform 1 0 42964 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_444
timestamp 1632082664
transform 1 0 41952 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_472
timestamp 1632082664
transform 1 0 44528 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1632082664
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1036_
timestamp 1632082664
transform 1 0 45356 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_77_480
timestamp 1632082664
transform 1 0 45264 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0978_
timestamp 1632082664
transform 1 0 47564 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1632082664
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1632082664
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0980_
timestamp 1632082664
transform 1 0 49404 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_77_541
timestamp 1632082664
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_521
timestamp 1632082664
transform 1 0 49036 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1632082664
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1632082664
transform 1 0 52716 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1632082664
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1632082664
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1632082664
transform 1 0 54556 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_77_577
timestamp 1632082664
transform 1 0 54188 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_597
timestamp 1632082664
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1632082664
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_617
timestamp 1632082664
transform 1 0 57868 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1632082664
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1632082664
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_629
timestamp 1632082664
transform 1 0 58972 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1632082664
transform -1 0 59340 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0769_
timestamp 1632082664
transform 1 0 1748 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_78_3
timestamp 1632082664
transform 1 0 1380 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1632082664
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1632082664
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1632082664
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1632082664
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1632082664
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_23
timestamp 1632082664
transform 1 0 3220 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0765_
timestamp 1632082664
transform 1 0 6348 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_78_53
timestamp 1632082664
transform 1 0 5980 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_73
timestamp 1632082664
transform 1 0 7820 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_81
timestamp 1632082664
transform 1 0 8556 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0790_
timestamp 1632082664
transform 1 0 8924 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1632082664
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_101
timestamp 1632082664
transform 1 0 10396 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0791_
timestamp 1632082664
transform 1 0 10764 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1632082664
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1632082664
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0706_
timestamp 1632082664
transform 1 0 14076 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1632082664
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1632082664
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_157
timestamp 1632082664
transform 1 0 15548 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_187
timestamp 1632082664
transform 1 0 18308 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_169
timestamp 1632082664
transform 1 0 16652 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1105_
timestamp 1632082664
transform 1 0 16836 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_78_197
timestamp 1632082664
transform 1 0 19228 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0370_
timestamp 1632082664
transform 1 0 19964 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1632082664
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1632082664
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0368_
timestamp 1632082664
transform 1 0 21804 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_78_221
timestamp 1632082664
transform 1 0 21436 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_241
timestamp 1632082664
transform 1 0 23276 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_249
timestamp 1632082664
transform 1 0 24012 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1632082664
transform 1 0 25760 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1632082664
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1632082664
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_78_265
timestamp 1632082664
transform 1 0 25484 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp 1632082664
transform 1 0 27600 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_78_284
timestamp 1632082664
transform 1 0 27232 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_309
timestamp 1632082664
transform 1 0 29532 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1632082664
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_304
timestamp 1632082664
transform 1 0 29072 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp 1632082664
transform 1 0 30268 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_78_333
timestamp 1632082664
transform 1 0 31740 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_353
timestamp 1632082664
transform 1 0 33580 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1632082664
transform 1 0 32108 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1632082664
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1632082664
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_78_361
timestamp 1632082664
transform 1 0 34316 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1632082664
transform 1 0 36064 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_78_377
timestamp 1632082664
transform 1 0 35788 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1632082664
transform 1 0 37904 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_78_416
timestamp 1632082664
transform 1 0 39376 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_396
timestamp 1632082664
transform 1 0 37536 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_421
timestamp 1632082664
transform 1 0 39836 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1632082664
transform 1 0 40572 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1632082664
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 1632082664
transform 1 0 42412 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_78_445
timestamp 1632082664
transform 1 0 42044 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_477
timestamp 1632082664
transform 1 0 44988 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_465
timestamp 1632082664
transform 1 0 43884 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1632082664
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_78_473
timestamp 1632082664
transform 1 0 44620 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1038_
timestamp 1632082664
transform 1 0 45724 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0977_
timestamp 1632082664
transform 1 0 47564 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_78_501
timestamp 1632082664
transform 1 0 47196 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_521
timestamp 1632082664
transform 1 0 49036 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1632082664
transform 1 0 50140 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1632082664
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_78_529
timestamp 1632082664
transform 1 0 49772 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1632082664
transform 1 0 51980 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_78_549
timestamp 1632082664
transform 1 0 51612 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1632082664
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_78_569
timestamp 1632082664
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 1632082664
transform 1 0 55292 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1632082664
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1632082664
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1632082664
transform 1 0 57132 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_78_625
timestamp 1632082664
transform 1 0 58604 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_605
timestamp 1632082664
transform 1 0 56764 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_629
timestamp 1632082664
transform 1 0 58972 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1632082664
transform -1 0 59340 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0773_
timestamp 1632082664
transform 1 0 1840 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0771_
timestamp 1632082664
transform 1 0 1840 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_80_7
timestamp 1632082664
transform 1 0 1748 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_7
timestamp 1632082664
transform 1 0 1748 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_3
timestamp 1632082664
transform 1 0 1380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_3
timestamp 1632082664
transform 1 0 1380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1632082664
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1632082664
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_29
timestamp 1632082664
transform 1 0 3772 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0779_
timestamp 1632082664
transform 1 0 4508 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0772_
timestamp 1632082664
transform 1 0 3680 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1632082664
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_24
timestamp 1632082664
transform 1 0 3312 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_24
timestamp 1632082664
transform 1 0 3312 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_57
timestamp 1632082664
transform 1 0 6348 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0784_
timestamp 1632082664
transform 1 0 6440 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_79_44
timestamp 1632082664
transform 1 0 5152 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1632082664
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_57
timestamp 1632082664
transform 1 0 6348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_53
timestamp 1632082664
transform 1 0 5980 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_74
timestamp 1632082664
transform 1 0 7912 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_82
timestamp 1632082664
transform 1 0 8648 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0786_
timestamp 1632082664
transform 1 0 7176 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_79_65
timestamp 1632082664
transform 1 0 7084 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_82
timestamp 1632082664
transform 1 0 8648 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_102
timestamp 1632082664
transform 1 0 10488 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0788_
timestamp 1632082664
transform 1 0 9016 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0787_
timestamp 1632082664
transform 1 0 8924 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1632082664
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_101
timestamp 1632082664
transform 1 0 10396 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_110
timestamp 1632082664
transform 1 0 11224 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0795_
timestamp 1632082664
transform 1 0 10764 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0794_
timestamp 1632082664
transform 1 0 11500 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_80_121
timestamp 1632082664
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1632082664
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1632082664
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0705_
timestamp 1632082664
transform 1 0 14076 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0703_
timestamp 1632082664
transform 1 0 14352 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_79_129
timestamp 1632082664
transform 1 0 12972 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1632082664
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1632082664
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_80_141
timestamp 1632082664
transform 1 0 14076 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_160
timestamp 1632082664
transform 1 0 15824 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_157
timestamp 1632082664
transform 1 0 15548 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_165
timestamp 1632082664
transform 1 0 16284 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_185
timestamp 1632082664
transform 1 0 18124 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0700_
timestamp 1632082664
transform 1 0 16652 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0699_
timestamp 1632082664
transform 1 0 16652 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_79_185
timestamp 1632082664
transform 1 0 18124 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1632082664
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_168
timestamp 1632082664
transform 1 0 16560 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_197
timestamp 1632082664
transform 1 0 19228 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0372_
timestamp 1632082664
transform 1 0 19688 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0371_
timestamp 1632082664
transform 1 0 19872 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1632082664
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_201
timestamp 1632082664
transform 1 0 19596 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_203
timestamp 1632082664
transform 1 0 19780 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_197
timestamp 1632082664
transform 1 0 19228 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_80_193
timestamp 1632082664
transform 1 0 18860 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0369_
timestamp 1632082664
transform 1 0 21804 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_80_218
timestamp 1632082664
transform 1 0 21160 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1632082664
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_220
timestamp 1632082664
transform 1 0 21344 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_241
timestamp 1632082664
transform 1 0 23276 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_230
timestamp 1632082664
transform 1 0 22264 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1103_
timestamp 1632082664
transform 1 0 22448 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_80_248
timestamp 1632082664
transform 1 0 23920 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_79_249
timestamp 1632082664
transform 1 0 24012 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp 1632082664
transform 1 0 24840 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1632082664
transform 1 0 24288 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_79_268
timestamp 1632082664
transform 1 0 25760 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1632082664
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_257
timestamp 1632082664
transform 1 0 24748 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_253
timestamp 1632082664
transform 1 0 24380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_286
timestamp 1632082664
transform 1 0 27416 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1632082664
transform 1 0 27600 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_80_274
timestamp 1632082664
transform 1 0 26312 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1632082664
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1632082664
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_309
timestamp 1632082664
transform 1 0 29532 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1632082664
transform 1 0 28336 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1632082664
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_304
timestamp 1632082664
transform 1 0 29072 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_312
timestamp 1632082664
transform 1 0 29808 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_79_293
timestamp 1632082664
transform 1 0 28060 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 1632082664
transform 1 0 30268 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp 1632082664
transform 1 0 30176 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_80_333
timestamp 1632082664
transform 1 0 31740 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_332
timestamp 1632082664
transform 1 0 31648 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_353
timestamp 1632082664
transform 1 0 33580 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1632082664
transform 1 0 33488 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0943_
timestamp 1632082664
transform 1 0 32108 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1632082664
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1632082664
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_349
timestamp 1632082664
transform 1 0 33212 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_365
timestamp 1632082664
transform 1 0 34684 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_373
timestamp 1632082664
transform 1 0 35420 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1632082664
transform 1 0 35328 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0952_
timestamp 1632082664
transform 1 0 35604 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1632082664
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_368
timestamp 1632082664
transform 1 0 34960 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_80_361
timestamp 1632082664
transform 1 0 34316 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_393
timestamp 1632082664
transform 1 0 37260 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0956_
timestamp 1632082664
transform 1 0 37444 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1632082664
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_391
timestamp 1632082664
transform 1 0 37076 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_388
timestamp 1632082664
transform 1 0 36800 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_411
timestamp 1632082664
transform 1 0 38916 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1632082664
transform 1 0 37996 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_80_421
timestamp 1632082664
transform 1 0 39836 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_437
timestamp 1632082664
transform 1 0 41308 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0961_
timestamp 1632082664
transform 1 0 39836 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0960_
timestamp 1632082664
transform 1 0 40572 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1632082664
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1632082664
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_417
timestamp 1632082664
transform 1 0 39468 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0966_
timestamp 1632082664
transform 1 0 42412 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0964_
timestamp 1632082664
transform 1 0 42412 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1632082664
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_445
timestamp 1632082664
transform 1 0 42044 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_79_445
timestamp 1632082664
transform 1 0 42044 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_465
timestamp 1632082664
transform 1 0 43884 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0971_
timestamp 1632082664
transform 1 0 44988 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0970_
timestamp 1632082664
transform 1 0 44252 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1632082664
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_465
timestamp 1632082664
transform 1 0 43884 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_80_473
timestamp 1632082664
transform 1 0 44620 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1632082664
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0975_
timestamp 1632082664
transform 1 0 46828 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_79_485
timestamp 1632082664
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_493
timestamp 1632082664
transform 1 0 46460 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0976_
timestamp 1632082664
transform 1 0 47564 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_80_513
timestamp 1632082664
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1632082664
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1632082664
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1632082664
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1632082664
transform 1 0 50232 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0486_
timestamp 1632082664
transform 1 0 50508 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_79_521
timestamp 1632082664
transform 1 0 49036 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1632082664
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1632082664
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_533
timestamp 1632082664
transform 1 0 50140 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_533
timestamp 1632082664
transform 1 0 50140 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_550
timestamp 1632082664
transform 1 0 51704 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_558
timestamp 1632082664
transform 1 0 52440 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1632082664
transform 1 0 52716 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1632082664
transform 1 0 52348 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1632082664
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_553
timestamp 1632082664
transform 1 0 51980 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1632082664
transform 1 0 54556 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_80_573
timestamp 1632082664
transform 1 0 53820 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_577
timestamp 1632082664
transform 1 0 54188 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1632082664
transform 1 0 55292 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_79_597
timestamp 1632082664
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1632082664
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_80_585
timestamp 1632082664
transform 1 0 54924 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1632082664
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_617
timestamp 1632082664
transform 1 0 57868 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_605
timestamp 1632082664
transform 1 0 56764 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_617
timestamp 1632082664
transform 1 0 57868 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1632082664
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1632082664
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_629
timestamp 1632082664
transform 1 0 58972 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_629
timestamp 1632082664
transform 1 0 58972 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1632082664
transform -1 0 59340 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1632082664
transform -1 0 59340 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_3
timestamp 1632082664
transform 1 0 1380 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0774_
timestamp 1632082664
transform 1 0 2392 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1632082664
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_81_11
timestamp 1632082664
transform 1 0 2116 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0775_
timestamp 1632082664
transform 1 0 4232 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_81_30
timestamp 1632082664
transform 1 0 3864 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_50
timestamp 1632082664
transform 1 0 5704 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0782_
timestamp 1632082664
transform 1 0 6348 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1632082664
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0785_
timestamp 1632082664
transform 1 0 8188 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_81_73
timestamp 1632082664
transform 1 0 7820 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1632082664
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1632082664
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0797_
timestamp 1632082664
transform 1 0 11500 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1632082664
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1632082664
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_141
timestamp 1632082664
transform 1 0 14076 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_129
timestamp 1632082664
transform 1 0 12972 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0702_
timestamp 1632082664
transform 1 0 14720 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_81_147
timestamp 1632082664
transform 1 0 14628 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_164
timestamp 1632082664
transform 1 0 16192 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0698_
timestamp 1632082664
transform 1 0 16744 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_81_186
timestamp 1632082664
transform 1 0 18216 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1632082664
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_169
timestamp 1632082664
transform 1 0 16652 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0373_
timestamp 1632082664
transform 1 0 19596 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_81_198
timestamp 1632082664
transform 1 0 19320 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1632082664
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_81_225
timestamp 1632082664
transform 1 0 21804 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1632082664
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1632082664
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_250
timestamp 1632082664
transform 1 0 24104 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1101_
timestamp 1632082664
transform 1 0 22632 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_81_233
timestamp 1632082664
transform 1 0 22540 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_258
timestamp 1632082664
transform 1 0 24840 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1632082664
transform 1 0 25024 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1632082664
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1632082664
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_276
timestamp 1632082664
transform 1 0 26496 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_293
timestamp 1632082664
transform 1 0 28060 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1077_
timestamp 1632082664
transform 1 0 28796 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1632082664
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_317
timestamp 1632082664
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0942_
timestamp 1632082664
transform 1 0 32108 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1632082664
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1632082664
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_353
timestamp 1632082664
transform 1 0 33580 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0947_
timestamp 1632082664
transform 1 0 33948 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_81_373
timestamp 1632082664
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1632082664
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0954_
timestamp 1632082664
transform 1 0 37260 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1632082664
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1632082664
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0959_
timestamp 1632082664
transform 1 0 39100 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_81_409
timestamp 1632082664
transform 1 0 38732 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_429
timestamp 1632082664
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1632082664
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0965_
timestamp 1632082664
transform 1 0 42412 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1632082664
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1632082664
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0967_
timestamp 1632082664
transform 1 0 44252 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_81_465
timestamp 1632082664
transform 1 0 43884 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1632082664
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_485
timestamp 1632082664
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0974_
timestamp 1632082664
transform 1 0 47564 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1632082664
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1632082664
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0485_
timestamp 1632082664
transform 1 0 50140 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_81_521
timestamp 1632082664
transform 1 0 49036 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_561
timestamp 1632082664
transform 1 0 52716 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_81_549
timestamp 1632082664
transform 1 0 51612 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1632082664
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_81_557
timestamp 1632082664
transform 1 0 52348 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_81_569
timestamp 1632082664
transform 1 0 53452 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1632082664
transform 1 0 53636 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 1632082664
transform 1 0 55568 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_81_591
timestamp 1632082664
transform 1 0 55476 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_587
timestamp 1632082664
transform 1 0 55108 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_608
timestamp 1632082664
transform 1 0 57040 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_617
timestamp 1632082664
transform 1 0 57868 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1632082664
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_629
timestamp 1632082664
transform 1 0 58972 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1632082664
transform -1 0 59340 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_3
timestamp 1632082664
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_15
timestamp 1632082664
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1632082664
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0776_
timestamp 1632082664
transform 1 0 3772 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1632082664
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1632082664
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0778_
timestamp 1632082664
transform 1 0 5612 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_82_45
timestamp 1632082664
transform 1 0 5244 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1632082664
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_82_65
timestamp 1632082664
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1632082664
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_97
timestamp 1632082664
transform 1 0 10028 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0796_
timestamp 1632082664
transform 1 0 10580 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_82_85
timestamp 1632082664
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1632082664
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_119
timestamp 1632082664
transform 1 0 12052 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_141
timestamp 1632082664
transform 1 0 14076 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_82_131
timestamp 1632082664
transform 1 0 13156 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1632082664
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1632082664
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_165
timestamp 1632082664
transform 1 0 16284 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0701_
timestamp 1632082664
transform 1 0 14812 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_82_187
timestamp 1632082664
transform 1 0 18308 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0697_
timestamp 1632082664
transform 1 0 16836 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0375_
timestamp 1632082664
transform 1 0 19504 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1632082664
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1632082664
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_82_197
timestamp 1632082664
transform 1 0 19228 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_216
timestamp 1632082664
transform 1 0 20976 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_228
timestamp 1632082664
transform 1 0 22080 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1099_
timestamp 1632082664
transform 1 0 22448 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_82_248
timestamp 1632082664
transform 1 0 23920 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_253
timestamp 1632082664
transform 1 0 24380 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1632082664
transform 1 0 25392 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1632082664
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_82_261
timestamp 1632082664
transform 1 0 25116 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_280
timestamp 1632082664
transform 1 0 26864 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 1632082664
transform 1 0 27600 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_82_309
timestamp 1632082664
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1632082664
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_304
timestamp 1632082664
transform 1 0 29072 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0941_
timestamp 1632082664
transform 1 0 31096 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_82_325
timestamp 1632082664
transform 1 0 31004 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_321
timestamp 1632082664
transform 1 0 30636 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_354
timestamp 1632082664
transform 1 0 33672 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_342
timestamp 1632082664
transform 1 0 32568 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_362
timestamp 1632082664
transform 1 0 34408 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0948_
timestamp 1632082664
transform 1 0 34684 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1632082664
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0951_
timestamp 1632082664
transform 1 0 36524 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_82_381
timestamp 1632082664
transform 1 0 36156 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1632082664
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_82_401
timestamp 1632082664
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0958_
timestamp 1632082664
transform 1 0 39836 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1632082664
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1632082664
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_437
timestamp 1632082664
transform 1 0 41308 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0963_
timestamp 1632082664
transform 1 0 41676 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_82_457
timestamp 1632082664
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1632082664
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0972_
timestamp 1632082664
transform 1 0 44988 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1632082664
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1632082664
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_493
timestamp 1632082664
transform 1 0 46460 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_505
timestamp 1632082664
transform 1 0 47564 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0481_
timestamp 1632082664
transform 1 0 48208 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_82_511
timestamp 1632082664
transform 1 0 48116 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0483_
timestamp 1632082664
transform 1 0 50600 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1632082664
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_537
timestamp 1632082664
transform 1 0 50508 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_533
timestamp 1632082664
transform 1 0 50140 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_528
timestamp 1632082664
transform 1 0 49680 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0490_
timestamp 1632082664
transform 1 0 52532 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_82_558
timestamp 1632082664
transform 1 0 52440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_554
timestamp 1632082664
transform 1 0 52072 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_575
timestamp 1632082664
transform 1 0 54004 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_601
timestamp 1632082664
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_589
timestamp 1632082664
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1632082664
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1632082664
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_613
timestamp 1632082664
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_625
timestamp 1632082664
transform 1 0 58604 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_629
timestamp 1632082664
transform 1 0 58972 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1632082664
transform -1 0 59340 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_83_15
timestamp 1632082664
transform 1 0 2484 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_3
timestamp 1632082664
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1632082664
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0777_
timestamp 1632082664
transform 1 0 3496 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_83_23
timestamp 1632082664
transform 1 0 3220 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_83_54
timestamp 1632082664
transform 1 0 6072 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0783_
timestamp 1632082664
transform 1 0 6348 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_83_42
timestamp 1632082664
transform 1 0 4968 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1632082664
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_73
timestamp 1632082664
transform 1 0 7820 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_97
timestamp 1632082664
transform 1 0 10028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_85
timestamp 1632082664
transform 1 0 8924 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_26_clk
timestamp 1632082664
transform 1 0 11868 0 -1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1632082664
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_113
timestamp 1632082664
transform 1 0 11500 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_83_109
timestamp 1632082664
transform 1 0 11132 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0800_
timestamp 1632082664
transform 1 0 14076 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_83_137
timestamp 1632082664
transform 1 0 13708 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_157
timestamp 1632082664
transform 1 0 15548 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_165
timestamp 1632082664
transform 1 0 16284 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0696_
timestamp 1632082664
transform 1 0 16928 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1632082664
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_83_169
timestamp 1632082664
transform 1 0 16652 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0376_
timestamp 1632082664
transform 1 0 19504 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_83_188
timestamp 1632082664
transform 1 0 18400 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_216
timestamp 1632082664
transform 1 0 20976 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_225
timestamp 1632082664
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1632082664
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1097_
timestamp 1632082664
transform 1 0 23000 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_83_237
timestamp 1632082664
transform 1 0 22908 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_254
timestamp 1632082664
transform 1 0 24472 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1093_
timestamp 1632082664
transform 1 0 25024 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_83_281
timestamp 1632082664
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1632082664
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_276
timestamp 1632082664
transform 1 0 26496 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_293
timestamp 1632082664
transform 1 0 28060 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 1632082664
transform 1 0 28612 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_83_327
timestamp 1632082664
transform 1 0 31188 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_315
timestamp 1632082664
transform 1 0 30084 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0940_
timestamp 1632082664
transform 1 0 32384 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1632082664
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1632082664
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_83_337
timestamp 1632082664
transform 1 0 32108 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0944_
timestamp 1632082664
transform 1 0 34224 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_83_356
timestamp 1632082664
transform 1 0 33856 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0953_
timestamp 1632082664
transform 1 0 37260 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_83_376
timestamp 1632082664
transform 1 0 35696 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1632082664
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_388
timestamp 1632082664
transform 1 0 36800 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_409
timestamp 1632082664
transform 1 0 38732 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_49_clk
timestamp 1632082664
transform 1 0 39652 0 -1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_83_417
timestamp 1632082664
transform 1 0 39468 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_83_449
timestamp 1632082664
transform 1 0 42412 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_83_439
timestamp 1632082664
transform 1 0 41492 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0443_
timestamp 1632082664
transform 1 0 43056 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1632082664
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_83_455
timestamp 1632082664
transform 1 0 42964 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1632082664
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0969_
timestamp 1632082664
transform 1 0 44896 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_83_472
timestamp 1632082664
transform 1 0 44528 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_492
timestamp 1632082664
transform 1 0 46368 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_63_clk
timestamp 1632082664
transform 1 0 48760 0 -1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_83_505
timestamp 1632082664
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1632082664
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_83_517
timestamp 1632082664
transform 1 0 48668 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_538
timestamp 1632082664
transform 1 0 50600 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_550
timestamp 1632082664
transform 1 0 51704 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_558
timestamp 1632082664
transform 1 0 52440 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0487_
timestamp 1632082664
transform 1 0 52716 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1632082664
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_577
timestamp 1632082664
transform 1 0 54188 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_601
timestamp 1632082664
transform 1 0 56396 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_589
timestamp 1632082664
transform 1 0 55292 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_617
timestamp 1632082664
transform 1 0 57868 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1632082664
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_83_613
timestamp 1632082664
transform 1 0 57500 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_83_629
timestamp 1632082664
transform 1 0 58972 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1632082664
transform -1 0 59340 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_3
timestamp 1632082664
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_15
timestamp 1632082664
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1632082664
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_29
timestamp 1632082664
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1632082664
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_84_41
timestamp 1632082664
transform 1 0 4876 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1632082664
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0780_
timestamp 1632082664
transform 1 0 4968 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_84_58
timestamp 1632082664
transform 1 0 6440 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_84_82
timestamp 1632082664
transform 1 0 8648 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_84_70
timestamp 1632082664
transform 1 0 7544 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0812_
timestamp 1632082664
transform 1 0 9384 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1632082664
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_84_89
timestamp 1632082664
transform 1 0 9292 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_85
timestamp 1632082664
transform 1 0 8924 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_106
timestamp 1632082664
transform 1 0 10856 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0798_
timestamp 1632082664
transform 1 0 11500 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_84_112
timestamp 1632082664
transform 1 0 11408 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_84_141
timestamp 1632082664
transform 1 0 14076 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_84_129
timestamp 1632082664
transform 1 0 12972 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1632082664
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_84_137
timestamp 1632082664
transform 1 0 13708 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_84_163
timestamp 1632082664
transform 1 0 16100 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0802_
timestamp 1632082664
transform 1 0 14628 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_84_171
timestamp 1632082664
transform 1 0 16836 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0695_
timestamp 1632082664
transform 1 0 17020 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1632082664
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_84_197
timestamp 1632082664
transform 1 0 19228 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0377_
timestamp 1632082664
transform 1 0 19412 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1632082664
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1632082664
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_40_clk
timestamp 1632082664
transform 1 0 21252 0 1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_84_215
timestamp 1632082664
transform 1 0 20884 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_239
timestamp 1632082664
transform 1 0 23092 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_39_clk
timestamp 1632082664
transform 1 0 25668 0 1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_84_265
timestamp 1632082664
transform 1 0 25484 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_84_253
timestamp 1632082664
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1632082664
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1632082664
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_287
timestamp 1632082664
transform 1 0 27508 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_309
timestamp 1632082664
transform 1 0 29532 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_84_299
timestamp 1632082664
transform 1 0 28612 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1632082664
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1632082664
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0939_
timestamp 1632082664
transform 1 0 30360 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_84_317
timestamp 1632082664
transform 1 0 30268 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_354
timestamp 1632082664
transform 1 0 33672 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0937_
timestamp 1632082664
transform 1 0 32200 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_84_334
timestamp 1632082664
transform 1 0 31832 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_362
timestamp 1632082664
transform 1 0 34408 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0949_
timestamp 1632082664
transform 1 0 34684 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1632082664
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0950_
timestamp 1632082664
transform 1 0 36524 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_84_381
timestamp 1632082664
transform 1 0 36156 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1632082664
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_84_401
timestamp 1632082664
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0962_
timestamp 1632082664
transform 1 0 39836 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_84_437
timestamp 1632082664
transform 1 0 41308 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1632082664
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1632082664
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0439_
timestamp 1632082664
transform 1 0 42412 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_84_465
timestamp 1632082664
transform 1 0 43884 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0973_
timestamp 1632082664
transform 1 0 45080 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1632082664
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_84_477
timestamp 1632082664
transform 1 0 44988 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_84_473
timestamp 1632082664
transform 1 0 44620 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_494
timestamp 1632082664
transform 1 0 46552 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_506
timestamp 1632082664
transform 1 0 47656 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0480_
timestamp 1632082664
transform 1 0 48208 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0482_
timestamp 1632082664
transform 1 0 50140 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1632082664
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_528
timestamp 1632082664
transform 1 0 49680 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0488_
timestamp 1632082664
transform 1 0 51980 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_84_549
timestamp 1632082664
transform 1 0 51612 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1632082664
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_84_569
timestamp 1632082664
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0496_
timestamp 1632082664
transform 1 0 55292 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1632082664
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1632082664
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_617
timestamp 1632082664
transform 1 0 57868 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_605
timestamp 1632082664
transform 1 0 56764 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_629
timestamp 1632082664
transform 1 0 58972 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1632082664
transform -1 0 59340 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_85_3
timestamp 1632082664
transform 1 0 1380 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1632082664
transform 1 0 1380 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0833_
timestamp 1632082664
transform 1 0 1564 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0831_
timestamp 1632082664
transform 1 0 2116 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1632082664
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1632082664
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_86_41
timestamp 1632082664
transform 1 0 4876 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_86_21
timestamp 1632082664
transform 1 0 3036 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0830_
timestamp 1632082664
transform 1 0 3956 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_86_29
timestamp 1632082664
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1632082664
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1632082664
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_27
timestamp 1632082664
transform 1 0 3588 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_27_clk
timestamp 1632082664
transform 1 0 6808 0 -1 48960
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_85_47
timestamp 1632082664
transform 1 0 5428 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0828_
timestamp 1632082664
transform 1 0 5428 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1632082664
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_61
timestamp 1632082664
transform 1 0 6716 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1632082664
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_57
timestamp 1632082664
transform 1 0 6348 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_75
timestamp 1632082664
transform 1 0 8004 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_63
timestamp 1632082664
transform 1 0 6900 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1632082664
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_82
timestamp 1632082664
transform 1 0 8648 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_102
timestamp 1632082664
transform 1 0 10488 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0810_
timestamp 1632082664
transform 1 0 9016 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0809_
timestamp 1632082664
transform 1 0 8924 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_86_101
timestamp 1632082664
transform 1 0 10396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1632082664
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_86_113
timestamp 1632082664
transform 1 0 11500 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_85_113
timestamp 1632082664
transform 1 0 11500 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_110
timestamp 1632082664
transform 1 0 11224 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0806_
timestamp 1632082664
transform 1 0 12144 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0799_
timestamp 1632082664
transform 1 0 11684 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1632082664
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_86_119
timestamp 1632082664
transform 1 0 12052 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0805_
timestamp 1632082664
transform 1 0 14076 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0801_
timestamp 1632082664
transform 1 0 13524 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1632082664
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_136
timestamp 1632082664
transform 1 0 13616 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_131
timestamp 1632082664
transform 1 0 13156 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_157
timestamp 1632082664
transform 1 0 15548 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_151
timestamp 1632082664
transform 1 0 14996 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_163
timestamp 1632082664
transform 1 0 16100 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_169
timestamp 1632082664
transform 1 0 16652 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0694_
timestamp 1632082664
transform 1 0 16928 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0692_
timestamp 1632082664
transform 1 0 17204 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1632082664
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1632082664
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_85_169
timestamp 1632082664
transform 1 0 16652 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0379_
timestamp 1632082664
transform 1 0 19688 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0378_
timestamp 1632082664
transform 1 0 19596 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_85_188
timestamp 1632082664
transform 1 0 18400 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1632082664
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_86_201
timestamp 1632082664
transform 1 0 19596 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1632082664
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_200
timestamp 1632082664
transform 1 0 19504 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_197
timestamp 1632082664
transform 1 0 19228 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_191
timestamp 1632082664
transform 1 0 18676 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_225
timestamp 1632082664
transform 1 0 21804 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1632082664
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_86_218
timestamp 1632082664
transform 1 0 21160 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1632082664
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1632082664
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_86_230
timestamp 1632082664
transform 1 0 22264 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1102_
timestamp 1632082664
transform 1 0 22448 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1098_
timestamp 1632082664
transform 1 0 22448 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_85_248
timestamp 1632082664
transform 1 0 23920 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_85_231
timestamp 1632082664
transform 1 0 22356 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_248
timestamp 1632082664
transform 1 0 23920 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_253
timestamp 1632082664
transform 1 0 24380 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1095_
timestamp 1632082664
transform 1 0 25024 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1094_
timestamp 1632082664
transform 1 0 25024 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1632082664
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_86_259
timestamp 1632082664
transform 1 0 24932 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_288
timestamp 1632082664
transform 1 0 27600 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_276
timestamp 1632082664
transform 1 0 26496 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_281
timestamp 1632082664
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1632082664
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_276
timestamp 1632082664
transform 1 0 26496 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_300
timestamp 1632082664
transform 1 0 28704 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_85_305
timestamp 1632082664
transform 1 0 29164 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_293
timestamp 1632082664
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1632082664
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_309
timestamp 1632082664
transform 1 0 29532 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0938_
timestamp 1632082664
transform 1 0 30176 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0934_
timestamp 1632082664
transform 1 0 31740 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0932_
timestamp 1632082664
transform 1 0 29900 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_86_329
timestamp 1632082664
transform 1 0 31372 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_332
timestamp 1632082664
transform 1 0 31648 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_85_313
timestamp 1632082664
transform 1 0 29900 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0936_
timestamp 1632082664
transform 1 0 32108 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_86_349
timestamp 1632082664
transform 1 0 33212 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1632082664
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_353
timestamp 1632082664
transform 1 0 33580 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_50_clk
timestamp 1632082664
transform 1 0 35512 0 1 48960
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_86_365
timestamp 1632082664
transform 1 0 34684 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0945_
timestamp 1632082664
transform 1 0 33948 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_85_373
timestamp 1632082664
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1632082664
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_86_373
timestamp 1632082664
transform 1 0 35420 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_86_361
timestamp 1632082664
transform 1 0 34316 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1632082664
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0955_
timestamp 1632082664
transform 1 0 37260 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_86_394
timestamp 1632082664
transform 1 0 37352 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1632082664
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1632082664
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_406
timestamp 1632082664
transform 1 0 38456 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_409
timestamp 1632082664
transform 1 0 38732 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_421
timestamp 1632082664
transform 1 0 39836 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_86_418
timestamp 1632082664
transform 1 0 39560 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0436_
timestamp 1632082664
transform 1 0 40388 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0433_
timestamp 1632082664
transform 1 0 39836 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1632082664
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_437
timestamp 1632082664
transform 1 0 41308 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_449
timestamp 1632082664
transform 1 0 42412 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0438_
timestamp 1632082664
transform 1 0 43148 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0437_
timestamp 1632082664
transform 1 0 41676 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_86_457
timestamp 1632082664
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1632082664
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1632082664
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_443
timestamp 1632082664
transform 1 0 41860 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1632082664
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0446_
timestamp 1632082664
transform 1 0 44988 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0444_
timestamp 1632082664
transform 1 0 44988 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1632082664
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1632082664
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_473
timestamp 1632082664
transform 1 0 44620 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_493
timestamp 1632082664
transform 1 0 46460 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_493
timestamp 1632082664
transform 1 0 46460 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_505
timestamp 1632082664
transform 1 0 47564 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0478_
timestamp 1632082664
transform 1 0 48208 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0477_
timestamp 1632082664
transform 1 0 48760 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_85_505
timestamp 1632082664
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1632082664
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_86_511
timestamp 1632082664
transform 1 0 48116 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_517
timestamp 1632082664
transform 1 0 48668 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_85_501
timestamp 1632082664
transform 1 0 47196 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0479_
timestamp 1632082664
transform 1 0 50140 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_85_534
timestamp 1632082664
transform 1 0 50232 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1632082664
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_528
timestamp 1632082664
transform 1 0 49680 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_558
timestamp 1632082664
transform 1 0 52440 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0489_
timestamp 1632082664
transform 1 0 52716 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_86_549
timestamp 1632082664
transform 1 0 51612 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_546
timestamp 1632082664
transform 1 0 51336 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1632082664
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_561
timestamp 1632082664
transform 1 0 52716 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_62_clk
timestamp 1632082664
transform 1 0 53176 0 -1 48960
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_86_577
timestamp 1632082664
transform 1 0 54188 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_565
timestamp 1632082664
transform 1 0 53084 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0494_
timestamp 1632082664
transform 1 0 55292 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0492_
timestamp 1632082664
transform 1 0 55384 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1632082664
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_586
timestamp 1632082664
transform 1 0 55016 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_86_585
timestamp 1632082664
transform 1 0 54924 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_85_606
timestamp 1632082664
transform 1 0 56856 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_614
timestamp 1632082664
transform 1 0 57592 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0504_
timestamp 1632082664
transform 1 0 57132 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_85_617
timestamp 1632082664
transform 1 0 57868 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1632082664
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_625
timestamp 1632082664
transform 1 0 58604 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_605
timestamp 1632082664
transform 1 0 56764 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_629
timestamp 1632082664
transform 1 0 58972 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_629
timestamp 1632082664
transform 1 0 58972 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1632082664
transform -1 0 59340 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1632082664
transform -1 0 59340 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_87_3
timestamp 1632082664
transform 1 0 1380 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0832_
timestamp 1632082664
transform 1 0 1564 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1632082664
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0829_
timestamp 1632082664
transform 1 0 4416 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_87_21
timestamp 1632082664
transform 1 0 3036 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_33
timestamp 1632082664
transform 1 0 4140 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0827_
timestamp 1632082664
transform 1 0 6348 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1632082664
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_52
timestamp 1632082664
transform 1 0 5888 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_87_73
timestamp 1632082664
transform 1 0 7820 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_102
timestamp 1632082664
transform 1 0 10488 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0811_
timestamp 1632082664
transform 1 0 9016 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_87_85
timestamp 1632082664
transform 1 0 8924 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_110
timestamp 1632082664
transform 1 0 11224 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_87_113
timestamp 1632082664
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1632082664
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_87_125
timestamp 1632082664
transform 1 0 12604 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0804_
timestamp 1632082664
transform 1 0 12880 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_87_144
timestamp 1632082664
transform 1 0 14352 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0807_
timestamp 1632082664
transform 1 0 14720 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_87_164
timestamp 1632082664
transform 1 0 16192 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_33_clk
timestamp 1632082664
transform 1 0 17020 0 -1 50048
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1632082664
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_169
timestamp 1632082664
transform 1 0 16652 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_193
timestamp 1632082664
transform 1 0 18860 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0380_
timestamp 1632082664
transform 1 0 19688 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_87_201
timestamp 1632082664
transform 1 0 19596 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_218
timestamp 1632082664
transform 1 0 21160 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_87_225
timestamp 1632082664
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1632082664
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_237
timestamp 1632082664
transform 1 0 22908 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0390_
timestamp 1632082664
transform 1 0 23092 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 1632082664
transform 1 0 24932 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_87_255
timestamp 1632082664
transform 1 0 24564 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0926_
timestamp 1632082664
transform 1 0 26956 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1632082664
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1632082664
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_275
timestamp 1632082664
transform 1 0 26404 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0928_
timestamp 1632082664
transform 1 0 28796 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_87_297
timestamp 1632082664
transform 1 0 28428 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1632082664
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_87_317
timestamp 1632082664
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_51_clk
timestamp 1632082664
transform 1 0 32476 0 -1 50048
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1632082664
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1632082664
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_337
timestamp 1632082664
transform 1 0 32108 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0422_
timestamp 1632082664
transform 1 0 34684 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_87_361
timestamp 1632082664
transform 1 0 34316 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_381
timestamp 1632082664
transform 1 0 36156 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0427_
timestamp 1632082664
transform 1 0 37260 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1632082664
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_87_389
timestamp 1632082664
transform 1 0 36892 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0432_
timestamp 1632082664
transform 1 0 39100 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_87_409
timestamp 1632082664
transform 1 0 38732 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_87_429
timestamp 1632082664
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_56_clk
timestamp 1632082664
transform 1 0 43148 0 -1 50048
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1632082664
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_87_449
timestamp 1632082664
transform 1 0 42412 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1632082664
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1632082664
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_477
timestamp 1632082664
transform 1 0 44988 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1632082664
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0442_
timestamp 1632082664
transform 1 0 45356 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0476_
timestamp 1632082664
transform 1 0 48760 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_87_505
timestamp 1632082664
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1632082664
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_87_517
timestamp 1632082664
transform 1 0 48668 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1632082664
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0475_
timestamp 1632082664
transform 1 0 50600 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_87_534
timestamp 1632082664
transform 1 0 50232 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_87_554
timestamp 1632082664
transform 1 0 52072 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1632082664
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_561
timestamp 1632082664
transform 1 0 52716 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0491_
timestamp 1632082664
transform 1 0 53084 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_87_581
timestamp 1632082664
transform 1 0 54556 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0493_
timestamp 1632082664
transform 1 0 54924 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_87_601
timestamp 1632082664
transform 1 0 56396 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_617
timestamp 1632082664
transform 1 0 57868 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1632082664
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_87_613
timestamp 1632082664
transform 1 0 57500 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_87_629
timestamp 1632082664
transform 1 0 58972 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1632082664
transform -1 0 59340 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0834_
timestamp 1632082664
transform 1 0 1840 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_88_7
timestamp 1632082664
transform 1 0 1748 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_3
timestamp 1632082664
transform 1 0 1380 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1632082664
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_28_clk
timestamp 1632082664
transform 1 0 4140 0 1 50048
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1632082664
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_29
timestamp 1632082664
transform 1 0 3772 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_24
timestamp 1632082664
transform 1 0 3312 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0823_
timestamp 1632082664
transform 1 0 6348 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_88_53
timestamp 1632082664
transform 1 0 5980 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_88_73
timestamp 1632082664
transform 1 0 7820 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_81
timestamp 1632082664
transform 1 0 8556 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_88_85
timestamp 1632082664
transform 1 0 8924 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_93
timestamp 1632082664
transform 1 0 9660 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0813_
timestamp 1632082664
transform 1 0 9844 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1632082664
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_111
timestamp 1632082664
transform 1 0 11316 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0808_
timestamp 1632082664
transform 1 0 12144 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_88_119
timestamp 1632082664
transform 1 0 12052 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0687_
timestamp 1632082664
transform 1 0 14168 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1632082664
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_88_141
timestamp 1632082664
transform 1 0 14076 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_136
timestamp 1632082664
transform 1 0 13616 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0689_
timestamp 1632082664
transform 1 0 16008 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_88_158
timestamp 1632082664
transform 1 0 15640 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_178
timestamp 1632082664
transform 1 0 17480 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_197
timestamp 1632082664
transform 1 0 19228 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_88_190
timestamp 1632082664
transform 1 0 18584 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0381_
timestamp 1632082664
transform 1 0 19872 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1632082664
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_88_203
timestamp 1632082664
transform 1 0 19780 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0382_
timestamp 1632082664
transform 1 0 21712 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_88_220
timestamp 1632082664
transform 1 0 21344 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_240
timestamp 1632082664
transform 1 0 23184 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0392_
timestamp 1632082664
transform 1 0 24380 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_88_269
timestamp 1632082664
transform 1 0 25852 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1632082664
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0925_
timestamp 1632082664
transform 1 0 26956 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_88_297
timestamp 1632082664
transform 1 0 28428 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0930_
timestamp 1632082664
transform 1 0 29532 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1632082664
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_88_305
timestamp 1632082664
transform 1 0 29164 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0933_
timestamp 1632082664
transform 1 0 31372 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_88_325
timestamp 1632082664
transform 1 0 31004 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_345
timestamp 1632082664
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1632082664
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0421_
timestamp 1632082664
transform 1 0 34684 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1632082664
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1632082664
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0424_
timestamp 1632082664
transform 1 0 36524 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_88_381
timestamp 1632082664
transform 1 0 36156 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1632082664
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_88_401
timestamp 1632082664
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0431_
timestamp 1632082664
transform 1 0 39836 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1632082664
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1632082664
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_437
timestamp 1632082664
transform 1 0 41308 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0435_
timestamp 1632082664
transform 1 0 41676 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_88_457
timestamp 1632082664
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1632082664
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0447_
timestamp 1632082664
transform 1 0 44988 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1632082664
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1632082664
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0448_
timestamp 1632082664
transform 1 0 46828 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_88_493
timestamp 1632082664
transform 1 0 46460 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_513
timestamp 1632082664
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_533
timestamp 1632082664
transform 1 0 50140 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1632082664
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0474_
timestamp 1632082664
transform 1 0 50692 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1632082664
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1632082664
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_555
timestamp 1632082664
transform 1 0 52164 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_579
timestamp 1632082664
transform 1 0 54372 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_567
timestamp 1632082664
transform 1 0 53268 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_589
timestamp 1632082664
transform 1 0 55292 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0497_
timestamp 1632082664
transform 1 0 56028 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1632082664
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1632082664
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_613
timestamp 1632082664
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_625
timestamp 1632082664
transform 1 0 58604 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_629
timestamp 1632082664
transform 1 0 58972 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1632082664
transform -1 0 59340 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_89_3
timestamp 1632082664
transform 1 0 1380 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0835_
timestamp 1632082664
transform 1 0 2024 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_89_9
timestamp 1632082664
transform 1 0 1932 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1632082664
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_89_26
timestamp 1632082664
transform 1 0 3496 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_34
timestamp 1632082664
transform 1 0 4232 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0826_
timestamp 1632082664
transform 1 0 4416 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_89_57
timestamp 1632082664
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1632082664
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_52
timestamp 1632082664
transform 1 0 5888 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0820_
timestamp 1632082664
transform 1 0 7728 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_89_69
timestamp 1632082664
transform 1 0 7452 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0817_
timestamp 1632082664
transform 1 0 9568 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_89_88
timestamp 1632082664
transform 1 0 9200 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_89_113
timestamp 1632082664
transform 1 0 11500 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0815_
timestamp 1632082664
transform 1 0 11684 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1632082664
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_108
timestamp 1632082664
transform 1 0 11040 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_89_131
timestamp 1632082664
transform 1 0 13156 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_139
timestamp 1632082664
transform 1 0 13892 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0686_
timestamp 1632082664
transform 1 0 14076 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_89_157
timestamp 1632082664
transform 1 0 15548 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_89_165
timestamp 1632082664
transform 1 0 16284 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0690_
timestamp 1632082664
transform 1 0 16652 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_89_185
timestamp 1632082664
transform 1 0 18124 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1632082664
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_89_197
timestamp 1632082664
transform 1 0 19228 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0383_
timestamp 1632082664
transform 1 0 19872 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_89_203
timestamp 1632082664
transform 1 0 19780 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0386_
timestamp 1632082664
transform 1 0 21804 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1632082664
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_220
timestamp 1632082664
transform 1 0 21344 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0388_
timestamp 1632082664
transform 1 0 23644 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_89_241
timestamp 1632082664
transform 1 0 23276 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_261
timestamp 1632082664
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1632082664
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0923_
timestamp 1632082664
transform 1 0 26956 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1632082664
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1632082664
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0927_
timestamp 1632082664
transform 1 0 28796 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_89_297
timestamp 1632082664
transform 1 0 28428 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1632082664
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_89_317
timestamp 1632082664
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0417_
timestamp 1632082664
transform 1 0 33212 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_89_337
timestamp 1632082664
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1632082664
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1632082664
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0420_
timestamp 1632082664
transform 1 0 35052 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_89_365
timestamp 1632082664
transform 1 0 34684 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1632082664
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0426_
timestamp 1632082664
transform 1 0 37260 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1632082664
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1632082664
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0428_
timestamp 1632082664
transform 1 0 39100 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_89_409
timestamp 1632082664
transform 1 0 38732 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_429
timestamp 1632082664
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1632082664
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0441_
timestamp 1632082664
transform 1 0 42412 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1632082664
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1632082664
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0445_
timestamp 1632082664
transform 1 0 44252 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_89_465
timestamp 1632082664
transform 1 0 43884 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1632082664
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_89_485
timestamp 1632082664
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0450_
timestamp 1632082664
transform 1 0 47564 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1632082664
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1632082664
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_89_533
timestamp 1632082664
transform 1 0 50140 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0472_
timestamp 1632082664
transform 1 0 50784 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_89_521
timestamp 1632082664
transform 1 0 49036 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_89_539
timestamp 1632082664
transform 1 0 50692 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_561
timestamp 1632082664
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1632082664
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_556
timestamp 1632082664
transform 1 0 52256 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_573
timestamp 1632082664
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_585
timestamp 1632082664
transform 1 0 54924 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0498_
timestamp 1632082664
transform 1 0 55752 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_89_593
timestamp 1632082664
transform 1 0 55660 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_89_610
timestamp 1632082664
transform 1 0 57224 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_89_617
timestamp 1632082664
transform 1 0 57868 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1632082664
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_89_629
timestamp 1632082664
transform 1 0 58972 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1632082664
transform -1 0 59340 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0837_
timestamp 1632082664
transform 1 0 1840 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_90_7
timestamp 1632082664
transform 1 0 1748 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_3
timestamp 1632082664
transform 1 0 1380 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1632082664
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_29
timestamp 1632082664
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1632082664
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_24
timestamp 1632082664
transform 1 0 3312 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_90_41
timestamp 1632082664
transform 1 0 4876 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0824_
timestamp 1632082664
transform 1 0 5152 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_90_60
timestamp 1632082664
transform 1 0 6624 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0821_
timestamp 1632082664
transform 1 0 6992 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_90_80
timestamp 1632082664
transform 1 0 8464 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_90_97
timestamp 1632082664
transform 1 0 10028 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0816_
timestamp 1632082664
transform 1 0 10212 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_90_85
timestamp 1632082664
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1632082664
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0683_
timestamp 1632082664
transform 1 0 12052 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_90_115
timestamp 1632082664
transform 1 0 11684 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0685_
timestamp 1632082664
transform 1 0 14076 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1632082664
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1632082664
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_135
timestamp 1632082664
transform 1 0 13524 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0688_
timestamp 1632082664
transform 1 0 15916 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_90_157
timestamp 1632082664
transform 1 0 15548 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_90_177
timestamp 1632082664
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_clk
timestamp 1632082664
transform 1 0 19964 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1632082664
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_90_197
timestamp 1632082664
transform 1 0 19228 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1632082664
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1632082664
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_208
timestamp 1632082664
transform 1 0 20240 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0384_
timestamp 1632082664
transform 1 0 20700 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_90_229
timestamp 1632082664
transform 1 0 22172 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_212
timestamp 1632082664
transform 1 0 20608 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_241
timestamp 1632082664
transform 1 0 23276 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_90_249
timestamp 1632082664
transform 1 0 24012 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0389_
timestamp 1632082664
transform 1 0 24380 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_90_269
timestamp 1632082664
transform 1 0 25852 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1632082664
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_38_clk
timestamp 1632082664
transform 1 0 27232 0 1 51136
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_90_281
timestamp 1632082664
transform 1 0 26956 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0931_
timestamp 1632082664
transform 1 0 29532 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1632082664
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_304
timestamp 1632082664
transform 1 0 29072 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_90_325
timestamp 1632082664
transform 1 0 31004 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_337
timestamp 1632082664
transform 1 0 32108 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0416_
timestamp 1632082664
transform 1 0 32752 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_90_343
timestamp 1632082664
transform 1 0 32660 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0419_
timestamp 1632082664
transform 1 0 34684 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1632082664
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_360
timestamp 1632082664
transform 1 0 34224 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0425_
timestamp 1632082664
transform 1 0 36524 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_90_381
timestamp 1632082664
transform 1 0 36156 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1632082664
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_90_401
timestamp 1632082664
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0434_
timestamp 1632082664
transform 1 0 39836 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_90_437
timestamp 1632082664
transform 1 0 41308 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1632082664
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1632082664
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_449
timestamp 1632082664
transform 1 0 42412 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_477
timestamp 1632082664
transform 1 0 44988 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_461
timestamp 1632082664
transform 1 0 43516 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1632082664
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_90_473
timestamp 1632082664
transform 1 0 44620 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0449_
timestamp 1632082664
transform 1 0 45816 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_90_485
timestamp 1632082664
transform 1 0 45724 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0452_
timestamp 1632082664
transform 1 0 47656 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_90_502
timestamp 1632082664
transform 1 0 47288 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_90_533
timestamp 1632082664
transform 1 0 50140 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_90_522
timestamp 1632082664
transform 1 0 49128 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_530
timestamp 1632082664
transform 1 0 49864 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0471_
timestamp 1632082664
transform 1 0 50876 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1632082664
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_90_557
timestamp 1632082664
transform 1 0 52348 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_90_579
timestamp 1632082664
transform 1 0 54372 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0505_
timestamp 1632082664
transform 1 0 52900 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_61_clk
timestamp 1632082664
transform 1 0 55844 0 1 51136
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_90_589
timestamp 1632082664
transform 1 0 55292 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1632082664
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1632082664
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_615
timestamp 1632082664
transform 1 0 57684 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1632082664
transform -1 0 59340 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_90_627
timestamp 1632082664
transform 1 0 58788 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_91_3
timestamp 1632082664
transform 1 0 1380 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0838_
timestamp 1632082664
transform 1 0 2024 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_91_9
timestamp 1632082664
transform 1 0 1932 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1632082664
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_38
timestamp 1632082664
transform 1 0 4600 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_26
timestamp 1632082664
transform 1 0 3496 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_50
timestamp 1632082664
transform 1 0 5704 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_91_57
timestamp 1632082664
transform 1 0 6348 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0822_
timestamp 1632082664
transform 1 0 6532 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1632082664
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_75
timestamp 1632082664
transform 1 0 8004 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0818_
timestamp 1632082664
transform 1 0 9568 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_91_91
timestamp 1632082664
transform 1 0 9476 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_87
timestamp 1632082664
transform 1 0 9108 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0680_
timestamp 1632082664
transform 1 0 11500 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1632082664
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_108
timestamp 1632082664
transform 1 0 11040 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_clk
timestamp 1632082664
transform 1 0 13340 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0684_
timestamp 1632082664
transform 1 0 14076 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_91_140
timestamp 1632082664
transform 1 0 13984 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_136
timestamp 1632082664
transform 1 0 13616 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_129
timestamp 1632082664
transform 1 0 12972 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_91_157
timestamp 1632082664
transform 1 0 15548 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_165
timestamp 1632082664
transform 1 0 16284 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0691_
timestamp 1632082664
transform 1 0 16652 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_91_185
timestamp 1632082664
transform 1 0 18124 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1632082664
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0906_
timestamp 1632082664
transform 1 0 19228 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_91_213
timestamp 1632082664
transform 1 0 20700 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0387_
timestamp 1632082664
transform 1 0 21804 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1632082664
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_91_221
timestamp 1632082664
transform 1 0 21436 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0391_
timestamp 1632082664
transform 1 0 23644 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_91_241
timestamp 1632082664
transform 1 0 23276 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_91_261
timestamp 1632082664
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1632082664
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0922_
timestamp 1632082664
transform 1 0 26956 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1632082664
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1632082664
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0929_
timestamp 1632082664
transform 1 0 28796 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_91_297
timestamp 1632082664
transform 1 0 28428 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1632082664
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_91_317
timestamp 1632082664
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_337
timestamp 1632082664
transform 1 0 32108 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0415_
timestamp 1632082664
transform 1 0 33120 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1632082664
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1632082664
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_91_345
timestamp 1632082664
transform 1 0 32844 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_91_364
timestamp 1632082664
transform 1 0 34592 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0423_
timestamp 1632082664
transform 1 0 35144 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_91_386
timestamp 1632082664
transform 1 0 36616 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1632082664
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_393
timestamp 1632082664
transform 1 0 37260 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0430_
timestamp 1632082664
transform 1 0 37720 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_91_414
timestamp 1632082664
transform 1 0 39192 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_91_397
timestamp 1632082664
transform 1 0 37628 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_clk
timestamp 1632082664
transform 1 0 40296 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_429
timestamp 1632082664
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1632082664
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_91_449
timestamp 1632082664
transform 1 0 42412 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0584_
timestamp 1632082664
transform 1 0 43148 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1632082664
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1632082664
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_473
timestamp 1632082664
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_clk
timestamp 1632082664
transform 1 0 46828 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_485
timestamp 1632082664
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_500
timestamp 1632082664
transform 1 0 47104 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0453_
timestamp 1632082664
transform 1 0 47564 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1632082664
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_91_533
timestamp 1632082664
transform 1 0 50140 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0470_
timestamp 1632082664
transform 1 0 50784 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_91_521
timestamp 1632082664
transform 1 0 49036 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_91_539
timestamp 1632082664
transform 1 0 50692 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1632082664
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_561
timestamp 1632082664
transform 1 0 52716 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_556
timestamp 1632082664
transform 1 0 52256 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0507_
timestamp 1632082664
transform 1 0 53084 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_91_581
timestamp 1632082664
transform 1 0 54556 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0499_
timestamp 1632082664
transform 1 0 55936 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_91_593
timestamp 1632082664
transform 1 0 55660 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_617
timestamp 1632082664
transform 1 0 57868 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1632082664
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_612
timestamp 1632082664
transform 1 0 57408 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_629
timestamp 1632082664
transform 1 0 58972 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1632082664
transform -1 0 59340 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_93_3
timestamp 1632082664
transform 1 0 1380 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0840_
timestamp 1632082664
transform 1 0 2116 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0839_
timestamp 1632082664
transform 1 0 1840 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_92_7
timestamp 1632082664
transform 1 0 1748 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_3
timestamp 1632082664
transform 1 0 1380 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1632082664
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1632082664
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_92_29
timestamp 1632082664
transform 1 0 3772 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0845_
timestamp 1632082664
transform 1 0 4416 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0841_
timestamp 1632082664
transform 1 0 3956 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1632082664
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_92_35
timestamp 1632082664
transform 1 0 4324 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_27
timestamp 1632082664
transform 1 0 3588 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_24
timestamp 1632082664
transform 1 0 3312 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_93_47
timestamp 1632082664
transform 1 0 5428 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_57
timestamp 1632082664
transform 1 0 6348 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0850_
timestamp 1632082664
transform 1 0 6532 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_92_52
timestamp 1632082664
transform 1 0 5888 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1632082664
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1632082664
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_76
timestamp 1632082664
transform 1 0 8096 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_75
timestamp 1632082664
transform 1 0 8004 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_64
timestamp 1632082664
transform 1 0 6992 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_103
timestamp 1632082664
transform 1 0 10580 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_85
timestamp 1632082664
transform 1 0 8924 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0819_
timestamp 1632082664
transform 1 0 9108 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_93_99
timestamp 1632082664
transform 1 0 10212 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_87
timestamp 1632082664
transform 1 0 9108 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1632082664
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_111
timestamp 1632082664
transform 1 0 11316 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0679_
timestamp 1632082664
transform 1 0 11500 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_93_113
timestamp 1632082664
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1632082664
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1632082664
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_125
timestamp 1632082664
transform 1 0 12604 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_32_clk
timestamp 1632082664
transform 1 0 13064 0 -1 53312
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_92_129
timestamp 1632082664
transform 1 0 12972 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0681_
timestamp 1632082664
transform 1 0 14076 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1632082664
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_93_129
timestamp 1632082664
transform 1 0 12972 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_92_137
timestamp 1632082664
transform 1 0 13708 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_93_162
timestamp 1632082664
transform 1 0 16008 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_93_150
timestamp 1632082664
transform 1 0 14904 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_157
timestamp 1632082664
transform 1 0 15548 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0901_
timestamp 1632082664
transform 1 0 17112 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0900_
timestamp 1632082664
transform 1 0 16652 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1632082664
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_92_173
timestamp 1632082664
transform 1 0 17020 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_185
timestamp 1632082664
transform 1 0 18124 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_169
timestamp 1632082664
transform 1 0 16652 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_92_190
timestamp 1632082664
transform 1 0 18584 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_92_197
timestamp 1632082664
transform 1 0 19228 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0905_
timestamp 1632082664
transform 1 0 19964 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0903_
timestamp 1632082664
transform 1 0 18492 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_93_205
timestamp 1632082664
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1632082664
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1632082664
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1104_
timestamp 1632082664
transform 1 0 21804 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_93_225
timestamp 1632082664
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1632082664
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1632082664
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_221
timestamp 1632082664
transform 1 0 21436 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_92_241
timestamp 1632082664
transform 1 0 23276 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0920_
timestamp 1632082664
transform 1 0 23184 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_93_237
timestamp 1632082664
transform 1 0 22908 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_92_249
timestamp 1632082664
transform 1 0 24012 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0394_
timestamp 1632082664
transform 1 0 25024 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0393_
timestamp 1632082664
transform 1 0 24840 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1632082664
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_92_257
timestamp 1632082664
transform 1 0 24748 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_256
timestamp 1632082664
transform 1 0 24656 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_253
timestamp 1632082664
transform 1 0 24380 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0921_
timestamp 1632082664
transform 1 0 26680 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_93_281
timestamp 1632082664
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1632082664
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_276
timestamp 1632082664
transform 1 0 26496 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_274
timestamp 1632082664
transform 1 0 26312 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_306
timestamp 1632082664
transform 1 0 29256 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0404_
timestamp 1632082664
transform 1 0 29440 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_93_293
timestamp 1632082664
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_309
timestamp 1632082664
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_294
timestamp 1632082664
transform 1 0 28152 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1632082664
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_93_305
timestamp 1632082664
transform 1 0 29164 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_92_333
timestamp 1632082664
transform 1 0 31740 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_324
timestamp 1632082664
transform 1 0 30912 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_321
timestamp 1632082664
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_92_341
timestamp 1632082664
transform 1 0 32476 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0412_
timestamp 1632082664
transform 1 0 32660 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0409_
timestamp 1632082664
transform 1 0 32108 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1632082664
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_353
timestamp 1632082664
transform 1 0 33580 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0414_
timestamp 1632082664
transform 1 0 33948 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_93_373
timestamp 1632082664
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_365
timestamp 1632082664
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1632082664
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1632082664
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_359
timestamp 1632082664
transform 1 0 34132 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1632082664
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_93_393
timestamp 1632082664
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_389
timestamp 1632082664
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_377
timestamp 1632082664
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1632082664
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1632082664
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1632082664
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0592_
timestamp 1632082664
transform 1 0 38640 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_92_401
timestamp 1632082664
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_405
timestamp 1632082664
transform 1 0 38364 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_92_421
timestamp 1632082664
transform 1 0 39836 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0589_
timestamp 1632082664
transform 1 0 40388 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0586_
timestamp 1632082664
transform 1 0 40480 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1632082664
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1632082664
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_424
timestamp 1632082664
transform 1 0 40112 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_93_449
timestamp 1632082664
transform 1 0 42412 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0581_
timestamp 1632082664
transform 1 0 43056 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_92_443
timestamp 1632082664
transform 1 0 41860 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1632082664
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_92_455
timestamp 1632082664
transform 1 0 42964 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_444
timestamp 1632082664
transform 1 0 41952 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_93_457
timestamp 1632082664
transform 1 0 43148 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0579_
timestamp 1632082664
transform 1 0 43424 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_92_477
timestamp 1632082664
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1632082664
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_476
timestamp 1632082664
transform 1 0 44896 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_472
timestamp 1632082664
transform 1 0 44528 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_93_496
timestamp 1632082664
transform 1 0 46736 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_92_489
timestamp 1632082664
transform 1 0 46092 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0578_
timestamp 1632082664
transform 1 0 45264 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0454_
timestamp 1632082664
transform 1 0 46920 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_92_497
timestamp 1632082664
transform 1 0 46828 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0455_
timestamp 1632082664
transform 1 0 47564 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_92_514
timestamp 1632082664
transform 1 0 48392 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1632082664
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_92_526
timestamp 1632082664
transform 1 0 49496 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_92_533
timestamp 1632082664
transform 1 0 50140 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_541
timestamp 1632082664
transform 1 0 50876 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_93_533
timestamp 1632082664
transform 1 0 50140 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_521
timestamp 1632082664
transform 1 0 49036 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1632082664
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_561
timestamp 1632082664
transform 1 0 52716 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_92_559
timestamp 1632082664
transform 1 0 52532 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0469_
timestamp 1632082664
transform 1 0 51060 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_93_545
timestamp 1632082664
transform 1 0 51244 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1632082664
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_93_557
timestamp 1632082664
transform 1 0 52348 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_93_569
timestamp 1632082664
transform 1 0 53452 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0509_
timestamp 1632082664
transform 1 0 53636 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0508_
timestamp 1632082664
transform 1 0 53360 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_92_567
timestamp 1632082664
transform 1 0 53268 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_587
timestamp 1632082664
transform 1 0 55108 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_92_589
timestamp 1632082664
transform 1 0 55292 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0502_
timestamp 1632082664
transform 1 0 55936 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0500_
timestamp 1632082664
transform 1 0 56304 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1632082664
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_93_595
timestamp 1632082664
transform 1 0 55844 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_584
timestamp 1632082664
transform 1 0 54832 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_92_597
timestamp 1632082664
transform 1 0 56028 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_617
timestamp 1632082664
transform 1 0 57868 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_616
timestamp 1632082664
transform 1 0 57776 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1632082664
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_612
timestamp 1632082664
transform 1 0 57408 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_628
timestamp 1632082664
transform 1 0 58880 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_93_629
timestamp 1632082664
transform 1 0 58972 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1632082664
transform -1 0 59340 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1632082664
transform -1 0 59340 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_3
timestamp 1632082664
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_15
timestamp 1632082664
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1632082664
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0843_
timestamp 1632082664
transform 1 0 3772 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1632082664
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1632082664
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0844_
timestamp 1632082664
transform 1 0 5612 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_94_45
timestamp 1632082664
transform 1 0 5244 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1632082664
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_94_65
timestamp 1632082664
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1632082664
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_85
timestamp 1632082664
transform 1 0 8924 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_93
timestamp 1632082664
transform 1 0 9660 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0676_
timestamp 1632082664
transform 1 0 9844 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1632082664
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0678_
timestamp 1632082664
transform 1 0 11684 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_94_111
timestamp 1632082664
transform 1 0 11316 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_94_131
timestamp 1632082664
transform 1 0 13156 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1632082664
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_94_145
timestamp 1632082664
transform 1 0 14444 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1632082664
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_141
timestamp 1632082664
transform 1 0 14076 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0898_
timestamp 1632082664
transform 1 0 16376 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0896_
timestamp 1632082664
transform 1 0 14536 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_94_162
timestamp 1632082664
transform 1 0 16008 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_182
timestamp 1632082664
transform 1 0 17848 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_94_194
timestamp 1632082664
transform 1 0 18952 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0904_
timestamp 1632082664
transform 1 0 19228 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1632082664
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0907_
timestamp 1632082664
transform 1 0 21068 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_94_213
timestamp 1632082664
transform 1 0 20700 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1632082664
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_94_233
timestamp 1632082664
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0395_
timestamp 1632082664
transform 1 0 25944 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_94_253
timestamp 1632082664
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1632082664
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_94_269
timestamp 1632082664
transform 1 0 25852 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1632082664
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_265
timestamp 1632082664
transform 1 0 25484 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_286
timestamp 1632082664
transform 1 0 27416 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_298
timestamp 1632082664
transform 1 0 28520 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_306
timestamp 1632082664
transform 1 0 29256 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0403_
timestamp 1632082664
transform 1 0 29532 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1632082664
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0405_
timestamp 1632082664
transform 1 0 31372 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_94_325
timestamp 1632082664
transform 1 0 31004 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_345
timestamp 1632082664
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1632082664
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0413_
timestamp 1632082664
transform 1 0 34684 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1632082664
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1632082664
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_94_393
timestamp 1632082664
transform 1 0 37260 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_94_381
timestamp 1632082664
transform 1 0 36156 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0595_
timestamp 1632082664
transform 1 0 37904 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_94_399
timestamp 1632082664
transform 1 0 37812 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_416
timestamp 1632082664
transform 1 0 39376 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0587_
timestamp 1632082664
transform 1 0 41216 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_94_421
timestamp 1632082664
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1632082664
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_94_433
timestamp 1632082664
transform 1 0 40940 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0582_
timestamp 1632082664
transform 1 0 43056 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_94_452
timestamp 1632082664
transform 1 0 42688 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1632082664
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_472
timestamp 1632082664
transform 1 0 44528 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_94_477
timestamp 1632082664
transform 1 0 44988 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_57_clk
timestamp 1632082664
transform 1 0 47104 0 1 53312
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _0577_
timestamp 1632082664
transform 1 0 45264 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_94_496
timestamp 1632082664
transform 1 0 46736 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_520
timestamp 1632082664
transform 1 0 48944 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_533
timestamp 1632082664
transform 1 0 50140 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_541
timestamp 1632082664
transform 1 0 50876 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1632082664
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0466_
timestamp 1632082664
transform 1 0 51060 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_94_559
timestamp 1632082664
transform 1 0 52532 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_94_579
timestamp 1632082664
transform 1 0 54372 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0468_
timestamp 1632082664
transform 1 0 52900 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_94_589
timestamp 1632082664
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1632082664
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1632082664
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_601
timestamp 1632082664
transform 1 0 56396 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_94_621
timestamp 1632082664
transform 1 0 58236 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0501_
timestamp 1632082664
transform 1 0 56764 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_94_629
timestamp 1632082664
transform 1 0 58972 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1632082664
transform -1 0 59340 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0842_
timestamp 1632082664
transform 1 0 2852 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_95_3
timestamp 1632082664
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_15
timestamp 1632082664
transform 1 0 2484 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1632082664
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_35
timestamp 1632082664
transform 1 0 4324 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_47
timestamp 1632082664
transform 1 0 5428 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0848_
timestamp 1632082664
transform 1 0 6348 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1632082664
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1632082664
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_73
timestamp 1632082664
transform 1 0 7820 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_85
timestamp 1632082664
transform 1 0 8924 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0675_
timestamp 1632082664
transform 1 0 9568 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_95_91
timestamp 1632082664
transform 1 0 9476 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0677_
timestamp 1632082664
transform 1 0 11500 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1632082664
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_108
timestamp 1632082664
transform 1 0 11040 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_141
timestamp 1632082664
transform 1 0 14076 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_95_129
timestamp 1632082664
transform 1 0 12972 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0895_
timestamp 1632082664
transform 1 0 14628 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_95_163
timestamp 1632082664
transform 1 0 16100 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_185
timestamp 1632082664
transform 1 0 18124 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0899_
timestamp 1632082664
transform 1 0 16652 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1632082664
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1632082664
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_34_clk
timestamp 1632082664
transform 1 0 18676 0 -1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _0909_
timestamp 1632082664
transform 1 0 21804 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_95_211
timestamp 1632082664
transform 1 0 20516 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1632082664
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1632082664
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0914_
timestamp 1632082664
transform 1 0 23644 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_95_241
timestamp 1632082664
transform 1 0 23276 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_95_261
timestamp 1632082664
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1632082664
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0397_
timestamp 1632082664
transform 1 0 26956 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1632082664
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1632082664
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0401_
timestamp 1632082664
transform 1 0 28796 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_95_297
timestamp 1632082664
transform 1 0 28428 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1632082664
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_95_317
timestamp 1632082664
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0406_
timestamp 1632082664
transform 1 0 32108 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1632082664
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1632082664
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_353
timestamp 1632082664
transform 1 0 33580 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0411_
timestamp 1632082664
transform 1 0 33948 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_95_373
timestamp 1632082664
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1632082664
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_95_393
timestamp 1632082664
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1632082664
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1632082664
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0593_
timestamp 1632082664
transform 1 0 38640 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_95_405
timestamp 1632082664
transform 1 0 38364 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0588_
timestamp 1632082664
transform 1 0 40480 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_95_424
timestamp 1632082664
transform 1 0 40112 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_95_449
timestamp 1632082664
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1632082664
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_444
timestamp 1632082664
transform 1 0 41952 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0580_
timestamp 1632082664
transform 1 0 43792 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_95_461
timestamp 1632082664
transform 1 0 43516 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0576_
timestamp 1632082664
transform 1 0 45632 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_95_500
timestamp 1632082664
transform 1 0 47104 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_480
timestamp 1632082664
transform 1 0 45264 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0456_
timestamp 1632082664
transform 1 0 47564 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1632082664
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0459_
timestamp 1632082664
transform 1 0 49496 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_95_525
timestamp 1632082664
transform 1 0 49404 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_521
timestamp 1632082664
transform 1 0 49036 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_554
timestamp 1632082664
transform 1 0 52072 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0467_
timestamp 1632082664
transform 1 0 52716 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_95_542
timestamp 1632082664
transform 1 0 50968 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1632082664
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_577
timestamp 1632082664
transform 1 0 54188 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_589
timestamp 1632082664
transform 1 0 55292 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0510_
timestamp 1632082664
transform 1 0 55476 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_95_607
timestamp 1632082664
transform 1 0 56948 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_617
timestamp 1632082664
transform 1 0 57868 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1632082664
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1632082664
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_95_629
timestamp 1632082664
transform 1 0 58972 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1632082664
transform -1 0 59340 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_3
timestamp 1632082664
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_15
timestamp 1632082664
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1632082664
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_96_41
timestamp 1632082664
transform 1 0 4876 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_96_29
timestamp 1632082664
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1632082664
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1632082664
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0846_
timestamp 1632082664
transform 1 0 5060 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_96_59
timestamp 1632082664
transform 1 0 6532 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0849_
timestamp 1632082664
transform 1 0 6900 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1632082664
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_79
timestamp 1632082664
transform 1 0 8372 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_96_85
timestamp 1632082664
transform 1 0 8924 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0674_
timestamp 1632082664
transform 1 0 9476 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1632082664
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_119
timestamp 1632082664
transform 1 0 12052 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_107
timestamp 1632082664
transform 1 0 10948 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_131
timestamp 1632082664
transform 1 0 13156 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0894_
timestamp 1632082664
transform 1 0 14076 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1632082664
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1632082664
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0897_
timestamp 1632082664
transform 1 0 15916 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_96_157
timestamp 1632082664
transform 1 0 15548 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_177
timestamp 1632082664
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_197
timestamp 1632082664
transform 1 0 19228 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1632082664
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0908_
timestamp 1632082664
transform 1 0 19872 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1632082664
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_96_203
timestamp 1632082664
transform 1 0 19780 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1632082664
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0910_
timestamp 1632082664
transform 1 0 21712 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_96_220
timestamp 1632082664
transform 1 0 21344 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_240
timestamp 1632082664
transform 1 0 23184 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_269
timestamp 1632082664
transform 1 0 25852 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0917_
timestamp 1632082664
transform 1 0 24380 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1632082664
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0398_
timestamp 1632082664
transform 1 0 26864 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_96_277
timestamp 1632082664
transform 1 0 26588 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0400_
timestamp 1632082664
transform 1 0 29532 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_96_296
timestamp 1632082664
transform 1 0 28336 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1632082664
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_325
timestamp 1632082664
transform 1 0 31004 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_52_clk
timestamp 1632082664
transform 1 0 32384 0 1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_96_337
timestamp 1632082664
transform 1 0 32108 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_96_365
timestamp 1632082664
transform 1 0 34684 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0597_
timestamp 1632082664
transform 1 0 35236 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1632082664
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_360
timestamp 1632082664
transform 1 0 34224 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0596_
timestamp 1632082664
transform 1 0 37076 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_96_387
timestamp 1632082664
transform 1 0 36708 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_407
timestamp 1632082664
transform 1 0 38548 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_96_421
timestamp 1632082664
transform 1 0 39836 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0590_
timestamp 1632082664
transform 1 0 40020 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1632082664
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1632082664
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0585_
timestamp 1632082664
transform 1 0 42964 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_96_439
timestamp 1632082664
transform 1 0 41492 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_451
timestamp 1632082664
transform 1 0 42596 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_96_477
timestamp 1632082664
transform 1 0 44988 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1632082664
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1632082664
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_471
timestamp 1632082664
transform 1 0 44436 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0575_
timestamp 1632082664
transform 1 0 45816 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_96_485
timestamp 1632082664
transform 1 0 45724 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0457_
timestamp 1632082664
transform 1 0 47656 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_96_502
timestamp 1632082664
transform 1 0 47288 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_96_522
timestamp 1632082664
transform 1 0 49128 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_530
timestamp 1632082664
transform 1 0 49864 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0461_
timestamp 1632082664
transform 1 0 50140 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1632082664
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0465_
timestamp 1632082664
transform 1 0 51980 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_96_549
timestamp 1632082664
transform 1 0 51612 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1632082664
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_96_569
timestamp 1632082664
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_601
timestamp 1632082664
transform 1 0 56396 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_96_589
timestamp 1632082664
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1632082664
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1632082664
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_96_624
timestamp 1632082664
transform 1 0 58512 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0503_
timestamp 1632082664
transform 1 0 57040 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_96_607
timestamp 1632082664
transform 1 0 56948 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1632082664
transform -1 0 59340 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_3
timestamp 1632082664
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_15
timestamp 1632082664
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1632082664
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_97_27
timestamp 1632082664
transform 1 0 3588 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0855_
timestamp 1632082664
transform 1 0 3772 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_97_45
timestamp 1632082664
transform 1 0 5244 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0851_
timestamp 1632082664
transform 1 0 6808 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1632082664
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_97_61
timestamp 1632082664
transform 1 0 6716 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_57
timestamp 1632082664
transform 1 0 6348 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_97_53
timestamp 1632082664
transform 1 0 5980 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_97_78
timestamp 1632082664
transform 1 0 8280 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0673_
timestamp 1632082664
transform 1 0 9292 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_97_86
timestamp 1632082664
transform 1 0 9016 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1632082664
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_97_113
timestamp 1632082664
transform 1 0 11500 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0892_
timestamp 1632082664
transform 1 0 12328 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1632082664
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_97_121
timestamp 1632082664
transform 1 0 12236 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1632082664
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0889_
timestamp 1632082664
transform 1 0 14168 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_97_138
timestamp 1632082664
transform 1 0 13800 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_97_158
timestamp 1632082664
transform 1 0 15640 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_166
timestamp 1632082664
transform 1 0 16376 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0666_
timestamp 1632082664
transform 1 0 17756 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_97_169
timestamp 1632082664
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1632082664
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0668_
timestamp 1632082664
transform 1 0 19596 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_97_197
timestamp 1632082664
transform 1 0 19228 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1632082664
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0911_
timestamp 1632082664
transform 1 0 21804 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1632082664
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1632082664
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0915_
timestamp 1632082664
transform 1 0 23644 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_97_241
timestamp 1632082664
transform 1 0 23276 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_97_261
timestamp 1632082664
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1632082664
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0399_
timestamp 1632082664
transform 1 0 27324 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1632082664
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1632082664
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_281
timestamp 1632082664
transform 1 0 26956 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0402_
timestamp 1632082664
transform 1 0 29164 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_97_301
timestamp 1632082664
transform 1 0 28796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_97_321
timestamp 1632082664
transform 1 0 30636 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_333
timestamp 1632082664
transform 1 0 31740 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0408_
timestamp 1632082664
transform 1 0 32108 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_97_353
timestamp 1632082664
transform 1 0 33580 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1632082664
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_97_365
timestamp 1632082664
transform 1 0 34684 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0598_
timestamp 1632082664
transform 1 0 35328 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_97_371
timestamp 1632082664
transform 1 0 35236 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_393
timestamp 1632082664
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1632082664
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_388
timestamp 1632082664
transform 1 0 36800 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0591_
timestamp 1632082664
transform 1 0 38640 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_97_405
timestamp 1632082664
transform 1 0 38364 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0566_
timestamp 1632082664
transform 1 0 40480 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_97_424
timestamp 1632082664
transform 1 0 40112 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_97_449
timestamp 1632082664
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1632082664
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_444
timestamp 1632082664
transform 1 0 41952 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0574_
timestamp 1632082664
transform 1 0 45080 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_97_461
timestamp 1632082664
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_97_477
timestamp 1632082664
transform 1 0 44988 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_473
timestamp 1632082664
transform 1 0 44620 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_97_494
timestamp 1632082664
transform 1 0 46552 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_502
timestamp 1632082664
transform 1 0 47288 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0458_
timestamp 1632082664
transform 1 0 48024 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1632082664
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_97_509
timestamp 1632082664
transform 1 0 47932 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_505
timestamp 1632082664
transform 1 0 47564 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0460_
timestamp 1632082664
transform 1 0 49864 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_97_526
timestamp 1632082664
transform 1 0 49496 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_558
timestamp 1632082664
transform 1 0 52440 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0464_
timestamp 1632082664
transform 1 0 52716 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_97_546
timestamp 1632082664
transform 1 0 51336 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1632082664
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0511_
timestamp 1632082664
transform 1 0 54556 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_97_577
timestamp 1632082664
transform 1 0 54188 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_97_597
timestamp 1632082664
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1632082664
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_97_617
timestamp 1632082664
transform 1 0 57868 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1632082664
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1632082664
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_97_629
timestamp 1632082664
transform 1 0 58972 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1632082664
transform -1 0 59340 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_3
timestamp 1632082664
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_15
timestamp 1632082664
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1632082664
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_29
timestamp 1632082664
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1632082664
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_98_41
timestamp 1632082664
transform 1 0 4876 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1632082664
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_29_clk
timestamp 1632082664
transform 1 0 4968 0 1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_98_62
timestamp 1632082664
transform 1 0 6808 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_74
timestamp 1632082664
transform 1 0 7912 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_82
timestamp 1632082664
transform 1 0 8648 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0672_
timestamp 1632082664
transform 1 0 8924 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_98_101
timestamp 1632082664
transform 1 0 10396 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1632082664
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_113
timestamp 1632082664
transform 1 0 11500 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0893_
timestamp 1632082664
transform 1 0 12144 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_98_119
timestamp 1632082664
transform 1 0 12052 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_141
timestamp 1632082664
transform 1 0 14076 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1632082664
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_136
timestamp 1632082664
transform 1 0 13616 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0888_
timestamp 1632082664
transform 1 0 14628 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_98_163
timestamp 1632082664
transform 1 0 16100 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0665_
timestamp 1632082664
transform 1 0 17296 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_98_175
timestamp 1632082664
transform 1 0 17204 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_197
timestamp 1632082664
transform 1 0 19228 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0659_
timestamp 1632082664
transform 1 0 19872 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1632082664
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_98_203
timestamp 1632082664
transform 1 0 19780 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_192
timestamp 1632082664
transform 1 0 18768 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0912_
timestamp 1632082664
transform 1 0 21712 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_98_220
timestamp 1632082664
transform 1 0 21344 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_240
timestamp 1632082664
transform 1 0 23184 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0918_
timestamp 1632082664
transform 1 0 24380 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_98_269
timestamp 1632082664
transform 1 0 25852 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1632082664
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_281
timestamp 1632082664
transform 1 0 26956 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0640_
timestamp 1632082664
transform 1 0 27140 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_98_299
timestamp 1632082664
transform 1 0 28612 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_309
timestamp 1632082664
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1632082664
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1632082664
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_321
timestamp 1632082664
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_333
timestamp 1632082664
transform 1 0 31740 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_353
timestamp 1632082664
transform 1 0 33580 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0410_
timestamp 1632082664
transform 1 0 32108 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_98_365
timestamp 1632082664
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1632082664
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_98_361
timestamp 1632082664
transform 1 0 34316 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0599_
timestamp 1632082664
transform 1 0 35788 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_98_393
timestamp 1632082664
transform 1 0 37260 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1632082664
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0600_
timestamp 1632082664
transform 1 0 37628 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_98_421
timestamp 1632082664
transform 1 0 39836 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0565_
timestamp 1632082664
transform 1 0 40020 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1632082664
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1632082664
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_55_clk
timestamp 1632082664
transform 1 0 41860 0 1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_98_439
timestamp 1632082664
transform 1 0 41492 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0571_
timestamp 1632082664
transform 1 0 44988 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_98_463
timestamp 1632082664
transform 1 0 43700 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1632082664
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1632082664
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_493
timestamp 1632082664
transform 1 0 46460 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0545_
timestamp 1632082664
transform 1 0 48024 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_98_509
timestamp 1632082664
transform 1 0 47932 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_505
timestamp 1632082664
transform 1 0 47564 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_98_526
timestamp 1632082664
transform 1 0 49496 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0463_
timestamp 1632082664
transform 1 0 50140 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1632082664
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_561
timestamp 1632082664
transform 1 0 52716 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_98_549
timestamp 1632082664
transform 1 0 51612 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0519_
timestamp 1632082664
transform 1 0 53360 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_98_567
timestamp 1632082664
transform 1 0 53268 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_60_clk
timestamp 1632082664
transform 1 0 56120 0 1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_98_589
timestamp 1632082664
transform 1 0 55292 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1632082664
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_98_597
timestamp 1632082664
transform 1 0 56028 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_584
timestamp 1632082664
transform 1 0 54832 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_618
timestamp 1632082664
transform 1 0 57960 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1632082664
transform -1 0 59340 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_3
timestamp 1632082664
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_15
timestamp 1632082664
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_3
timestamp 1632082664
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_15
timestamp 1632082664
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1632082664
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1632082664
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0857_
timestamp 1632082664
transform 1 0 3772 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0856_
timestamp 1632082664
transform 1 0 3588 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1632082664
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1632082664
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_99_57
timestamp 1632082664
transform 1 0 6348 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_100_57
timestamp 1632082664
transform 1 0 6348 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_99_43
timestamp 1632082664
transform 1 0 5060 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_45
timestamp 1632082664
transform 1 0 5244 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1632082664
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1632082664
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0853_
timestamp 1632082664
transform 1 0 6900 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0852_
timestamp 1632082664
transform 1 0 6900 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0670_
timestamp 1632082664
transform 1 0 8740 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1632082664
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_79
timestamp 1632082664
transform 1 0 8372 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_79
timestamp 1632082664
transform 1 0 8372 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0669_
timestamp 1632082664
transform 1 0 8924 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_99_99
timestamp 1632082664
transform 1 0 10212 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_101
timestamp 1632082664
transform 1 0 10396 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1632082664
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_99_125
timestamp 1632082664
transform 1 0 12604 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0877_
timestamp 1632082664
transform 1 0 11500 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_99_113
timestamp 1632082664
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1632082664
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1632082664
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_129
timestamp 1632082664
transform 1 0 12972 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0890_
timestamp 1632082664
transform 1 0 12788 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0885_
timestamp 1632082664
transform 1 0 14444 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1632082664
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_143
timestamp 1632082664
transform 1 0 14260 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_141
timestamp 1632082664
transform 1 0 14076 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_100_137
timestamp 1632082664
transform 1 0 13708 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0887_
timestamp 1632082664
transform 1 0 14720 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_100_161
timestamp 1632082664
transform 1 0 15916 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_99_147
timestamp 1632082664
transform 1 0 14628 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_164
timestamp 1632082664
transform 1 0 16192 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0663_
timestamp 1632082664
transform 1 0 17296 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0662_
timestamp 1632082664
transform 1 0 18032 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_99_169
timestamp 1632082664
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1632082664
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_99_181
timestamp 1632082664
transform 1 0 17756 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_100_173
timestamp 1632082664
transform 1 0 17020 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_100_197
timestamp 1632082664
transform 1 0 19228 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0658_
timestamp 1632082664
transform 1 0 19872 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0657_
timestamp 1632082664
transform 1 0 19872 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1632082664
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_100_203
timestamp 1632082664
transform 1 0 19780 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_200
timestamp 1632082664
transform 1 0 19504 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_192
timestamp 1632082664
transform 1 0 18768 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_225
timestamp 1632082664
transform 1 0 21804 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_100_220
timestamp 1632082664
transform 1 0 21344 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1632082664
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_220
timestamp 1632082664
transform 1 0 21344 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0652_
timestamp 1632082664
transform 1 0 22356 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0648_
timestamp 1632082664
transform 1 0 22448 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_99_247
timestamp 1632082664
transform 1 0 23828 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_248
timestamp 1632082664
transform 1 0 23920 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_36_clk
timestamp 1632082664
transform 1 0 24748 0 1 56576
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _0916_
timestamp 1632082664
transform 1 0 24196 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_99_267
timestamp 1632082664
transform 1 0 25668 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1632082664
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_253
timestamp 1632082664
transform 1 0 24380 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_281
timestamp 1632082664
transform 1 0 26956 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_100_277
timestamp 1632082664
transform 1 0 26588 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_285
timestamp 1632082664
transform 1 0 27324 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0637_
timestamp 1632082664
transform 1 0 27508 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1632082664
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1632082664
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_99_289
timestamp 1632082664
transform 1 0 27692 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_37_clk
timestamp 1632082664
transform 1 0 27968 0 -1 56576
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_100_309
timestamp 1632082664
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1632082664
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1632082664
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_312
timestamp 1632082664
transform 1 0 29808 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_303
timestamp 1632082664
transform 1 0 28980 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0919_
timestamp 1632082664
transform 1 0 30176 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0622_
timestamp 1632082664
transform 1 0 30912 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_99_332
timestamp 1632082664
transform 1 0 31648 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_100_321
timestamp 1632082664
transform 1 0 30636 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_99_337
timestamp 1632082664
transform 1 0 32108 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0620_
timestamp 1632082664
transform 1 0 32752 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0619_
timestamp 1632082664
transform 1 0 32844 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1632082664
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_340
timestamp 1632082664
transform 1 0 32384 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0618_
timestamp 1632082664
transform 1 0 34684 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0617_
timestamp 1632082664
transform 1 0 34684 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1632082664
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_361
timestamp 1632082664
transform 1 0 34316 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_360
timestamp 1632082664
transform 1 0 34224 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_381
timestamp 1632082664
transform 1 0 36156 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0602_
timestamp 1632082664
transform 1 0 37260 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_100_381
timestamp 1632082664
transform 1 0 36156 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1632082664
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_393
timestamp 1632082664
transform 1 0 37260 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_99_389
timestamp 1632082664
transform 1 0 36892 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_100_409
timestamp 1632082664
transform 1 0 38732 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0601_
timestamp 1632082664
transform 1 0 37628 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_99_413
timestamp 1632082664
transform 1 0 39100 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_421
timestamp 1632082664
transform 1 0 39836 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_425
timestamp 1632082664
transform 1 0 40204 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0563_
timestamp 1632082664
transform 1 0 40388 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0562_
timestamp 1632082664
transform 1 0 40848 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1632082664
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_100_429
timestamp 1632082664
transform 1 0 40572 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_100_417
timestamp 1632082664
transform 1 0 39468 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0567_
timestamp 1632082664
transform 1 0 42412 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0564_
timestamp 1632082664
transform 1 0 42688 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1632082664
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1632082664
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_443
timestamp 1632082664
transform 1 0 41860 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_448
timestamp 1632082664
transform 1 0 42320 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_468
timestamp 1632082664
transform 1 0 44160 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0573_
timestamp 1632082664
transform 1 0 44988 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0569_
timestamp 1632082664
transform 1 0 44252 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1632082664
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_465
timestamp 1632082664
transform 1 0 43884 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1632082664
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_99_485
timestamp 1632082664
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_493
timestamp 1632082664
transform 1 0 46460 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_505
timestamp 1632082664
transform 1 0 47564 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0543_
timestamp 1632082664
transform 1 0 48208 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0538_
timestamp 1632082664
transform 1 0 48944 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_99_505
timestamp 1632082664
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1632082664
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1632082664
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_100_511
timestamp 1632082664
transform 1 0 48116 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_99_517
timestamp 1632082664
transform 1 0 48668 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0535_
timestamp 1632082664
transform 1 0 50784 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_100_533
timestamp 1632082664
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1632082664
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_536
timestamp 1632082664
transform 1 0 50416 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_528
timestamp 1632082664
transform 1 0 49680 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0531_
timestamp 1632082664
transform 1 0 51520 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_99_561
timestamp 1632082664
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1632082664
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_556
timestamp 1632082664
transform 1 0 52256 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_100_545
timestamp 1632082664
transform 1 0 51244 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0522_
timestamp 1632082664
transform 1 0 53360 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0512_
timestamp 1632082664
transform 1 0 54280 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_99_577
timestamp 1632082664
transform 1 0 54188 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_573
timestamp 1632082664
transform 1 0 53820 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_564
timestamp 1632082664
transform 1 0 52992 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0513_
timestamp 1632082664
transform 1 0 55292 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_99_594
timestamp 1632082664
transform 1 0 55752 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1632082664
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_584
timestamp 1632082664
transform 1 0 54832 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_606
timestamp 1632082664
transform 1 0 56856 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_614
timestamp 1632082664
transform 1 0 57592 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0515_
timestamp 1632082664
transform 1 0 57132 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_99_617
timestamp 1632082664
transform 1 0 57868 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1632082664
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_625
timestamp 1632082664
transform 1 0 58604 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_605
timestamp 1632082664
transform 1 0 56764 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_629
timestamp 1632082664
transform 1 0 58972 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_100_629
timestamp 1632082664
transform 1 0 58972 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1632082664
transform -1 0 59340 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1632082664
transform -1 0 59340 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_3
timestamp 1632082664
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_15
timestamp 1632082664
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1632082664
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0859_
timestamp 1632082664
transform 1 0 3588 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_101_57
timestamp 1632082664
transform 1 0 6348 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_43
timestamp 1632082664
transform 1 0 5060 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1632082664
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_101_55
timestamp 1632082664
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_30_clk
timestamp 1632082664
transform 1 0 8740 0 -1 57664
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _0854_
timestamp 1632082664
transform 1 0 6900 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_101_79
timestamp 1632082664
transform 1 0 8372 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_103
timestamp 1632082664
transform 1 0 10580 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0874_
timestamp 1632082664
transform 1 0 11500 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1632082664
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_101_111
timestamp 1632082664
transform 1 0 11316 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0884_
timestamp 1632082664
transform 1 0 14076 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_101_129
timestamp 1632082664
transform 1 0 12972 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_157
timestamp 1632082664
transform 1 0 15548 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_165
timestamp 1632082664
transform 1 0 16284 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0661_
timestamp 1632082664
transform 1 0 18032 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_101_169
timestamp 1632082664
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1632082664
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_181
timestamp 1632082664
transform 1 0 17756 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0653_
timestamp 1632082664
transform 1 0 19872 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_101_200
timestamp 1632082664
transform 1 0 19504 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_101_225
timestamp 1632082664
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1632082664
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_220
timestamp 1632082664
transform 1 0 21344 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0647_
timestamp 1632082664
transform 1 0 23184 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_101_237
timestamp 1632082664
transform 1 0 22908 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0643_
timestamp 1632082664
transform 1 0 25024 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_101_256
timestamp 1632082664
transform 1 0 24656 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_281
timestamp 1632082664
transform 1 0 26956 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0636_
timestamp 1632082664
transform 1 0 27600 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1632082664
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_101_287
timestamp 1632082664
transform 1 0 27508 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_276
timestamp 1632082664
transform 1 0 26496 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_101_304
timestamp 1632082664
transform 1 0 29072 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0624_
timestamp 1632082664
transform 1 0 30176 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_101_332
timestamp 1632082664
transform 1 0 31648 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_337
timestamp 1632082664
transform 1 0 32108 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0621_
timestamp 1632082664
transform 1 0 32844 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1632082664
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0615_
timestamp 1632082664
transform 1 0 34684 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_101_361
timestamp 1632082664
transform 1 0 34316 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_381
timestamp 1632082664
transform 1 0 36156 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_101_393
timestamp 1632082664
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1632082664
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_389
timestamp 1632082664
transform 1 0 36892 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_54_clk
timestamp 1632082664
transform 1 0 39008 0 -1 57664
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_101_405
timestamp 1632082664
transform 1 0 38364 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_411
timestamp 1632082664
transform 1 0 38916 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_432
timestamp 1632082664
transform 1 0 40848 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0568_
timestamp 1632082664
transform 1 0 42412 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1632082664
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_444
timestamp 1632082664
transform 1 0 41952 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0570_
timestamp 1632082664
transform 1 0 44252 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_101_465
timestamp 1632082664
transform 1 0 43884 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_497
timestamp 1632082664
transform 1 0 46828 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_485
timestamp 1632082664
transform 1 0 45724 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0541_
timestamp 1632082664
transform 1 0 48944 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_101_505
timestamp 1632082664
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1632082664
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_101_503
timestamp 1632082664
transform 1 0 47380 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_517
timestamp 1632082664
transform 1 0 48668 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0534_
timestamp 1632082664
transform 1 0 50784 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_101_536
timestamp 1632082664
transform 1 0 50416 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1632082664
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_561
timestamp 1632082664
transform 1 0 52716 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_556
timestamp 1632082664
transform 1 0 52256 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_59_clk
timestamp 1632082664
transform 1 0 53084 0 -1 57664
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _0514_
timestamp 1632082664
transform 1 0 55292 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_101_585
timestamp 1632082664
transform 1 0 54924 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_605
timestamp 1632082664
transform 1 0 56764 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_101_617
timestamp 1632082664
transform 1 0 57868 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1632082664
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_613
timestamp 1632082664
transform 1 0 57500 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_101_629
timestamp 1632082664
transform 1 0 58972 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1632082664
transform -1 0 59340 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_102_3
timestamp 1632082664
transform 1 0 1380 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_15
timestamp 1632082664
transform 1 0 2484 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1632082664
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0860_
timestamp 1632082664
transform 1 0 3772 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1632082664
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1632082664
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0862_
timestamp 1632082664
transform 1 0 5612 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_102_45
timestamp 1632082664
transform 1 0 5244 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1632082664
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_102_65
timestamp 1632082664
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1632082664
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0872_
timestamp 1632082664
transform 1 0 8924 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1632082664
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_101
timestamp 1632082664
transform 1 0 10396 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0873_
timestamp 1632082664
transform 1 0 10764 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_102_121
timestamp 1632082664
transform 1 0 12236 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_31_clk
timestamp 1632082664
transform 1 0 14444 0 1 57664
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_102_133
timestamp 1632082664
transform 1 0 13340 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1632082664
transform 1 0 13984 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_102_139
timestamp 1632082664
transform 1 0 13892 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_141
timestamp 1632082664
transform 1 0 14076 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_102_165
timestamp 1632082664
transform 1 0 16284 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0664_
timestamp 1632082664
transform 1 0 17296 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_102_173
timestamp 1632082664
transform 1 0 17020 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_102_197
timestamp 1632082664
transform 1 0 19228 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1632082664
transform 1 0 19136 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_192
timestamp 1632082664
transform 1 0 18768 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_35_clk
timestamp 1632082664
transform 1 0 20424 0 1 57664
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_102_209
timestamp 1632082664
transform 1 0 20332 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_102_242
timestamp 1632082664
transform 1 0 23368 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_102_250
timestamp 1632082664
transform 1 0 24104 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_102_230
timestamp 1632082664
transform 1 0 22264 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0639_
timestamp 1632082664
transform 1 0 25760 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_102_253
timestamp 1632082664
transform 1 0 24380 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1632082664
transform 1 0 24288 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_102_265
timestamp 1632082664
transform 1 0 25484 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0635_
timestamp 1632082664
transform 1 0 27600 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_102_284
timestamp 1632082664
transform 1 0 27232 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_102_309
timestamp 1632082664
transform 1 0 29532 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1632082664
transform 1 0 29440 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_304
timestamp 1632082664
transform 1 0 29072 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0623_
timestamp 1632082664
transform 1 0 30912 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_102_321
timestamp 1632082664
transform 1 0 30636 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0614_
timestamp 1632082664
transform 1 0 32752 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_102_340
timestamp 1632082664
transform 1 0 32384 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_102_365
timestamp 1632082664
transform 1 0 34684 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0612_
timestamp 1632082664
transform 1 0 35328 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1632082664
transform 1 0 34592 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_102_371
timestamp 1632082664
transform 1 0 35236 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_360
timestamp 1632082664
transform 1 0 34224 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0603_
timestamp 1632082664
transform 1 0 37168 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_102_388
timestamp 1632082664
transform 1 0 36800 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_102_408
timestamp 1632082664
transform 1 0 38640 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_421
timestamp 1632082664
transform 1 0 39836 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0560_
timestamp 1632082664
transform 1 0 40388 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1632082664
transform 1 0 39744 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0556_
timestamp 1632082664
transform 1 0 43056 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_102_443
timestamp 1632082664
transform 1 0 41860 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_455
timestamp 1632082664
transform 1 0 42964 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_477
timestamp 1632082664
transform 1 0 44988 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1632082664
transform 1 0 44896 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_472
timestamp 1632082664
transform 1 0 44528 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0547_
timestamp 1632082664
transform 1 0 46368 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_102_489
timestamp 1632082664
transform 1 0 46092 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0537_
timestamp 1632082664
transform 1 0 48208 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_102_508
timestamp 1632082664
transform 1 0 47840 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_102_533
timestamp 1632082664
transform 1 0 50140 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1632082664
transform 1 0 50048 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_528
timestamp 1632082664
transform 1 0 49680 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0532_
timestamp 1632082664
transform 1 0 51520 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_102_545
timestamp 1632082664
transform 1 0 51244 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0525_
timestamp 1632082664
transform 1 0 53360 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_102_564
timestamp 1632082664
transform 1 0 52992 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0518_
timestamp 1632082664
transform 1 0 55292 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1632082664
transform 1 0 55200 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_584
timestamp 1632082664
transform 1 0 54832 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0516_
timestamp 1632082664
transform 1 0 57132 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_102_625
timestamp 1632082664
transform 1 0 58604 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_605
timestamp 1632082664
transform 1 0 56764 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_629
timestamp 1632082664
transform 1 0 58972 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1632082664
transform -1 0 59340 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_3
timestamp 1632082664
transform 1 0 1380 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_15
timestamp 1632082664
transform 1 0 2484 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1632082664
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_103_27
timestamp 1632082664
transform 1 0 3588 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0861_
timestamp 1632082664
transform 1 0 4140 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_103_49
timestamp 1632082664
transform 1 0 5612 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0864_
timestamp 1632082664
transform 1 0 6348 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1632082664
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1632082664
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0868_
timestamp 1632082664
transform 1 0 8188 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_103_73
timestamp 1632082664
transform 1 0 7820 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_103_93
timestamp 1632082664
transform 1 0 9660 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_105
timestamp 1632082664
transform 1 0 10764 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0876_
timestamp 1632082664
transform 1 0 11500 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1632082664
transform 1 0 11408 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_103_111
timestamp 1632082664
transform 1 0 11316 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0881_
timestamp 1632082664
transform 1 0 13340 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_103_129
timestamp 1632082664
transform 1 0 12972 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_103_161
timestamp 1632082664
transform 1 0 15916 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_103_149
timestamp 1632082664
transform 1 0 14812 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0667_
timestamp 1632082664
transform 1 0 18032 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_103_169
timestamp 1632082664
transform 1 0 16652 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1632082664
transform 1 0 16560 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_103_167
timestamp 1632082664
transform 1 0 16468 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_103_181
timestamp 1632082664
transform 1 0 17756 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0655_
timestamp 1632082664
transform 1 0 19872 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_103_200
timestamp 1632082664
transform 1 0 19504 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_103_225
timestamp 1632082664
transform 1 0 21804 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1632082664
transform 1 0 21712 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_220
timestamp 1632082664
transform 1 0 21344 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_103_233
timestamp 1632082664
transform 1 0 22540 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0646_
timestamp 1632082664
transform 1 0 22724 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0644_
timestamp 1632082664
transform 1 0 24564 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_103_251
timestamp 1632082664
transform 1 0 24196 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_103_281
timestamp 1632082664
transform 1 0 26956 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_103_271
timestamp 1632082664
transform 1 0 26036 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_103_289
timestamp 1632082664
transform 1 0 27692 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0634_
timestamp 1632082664
transform 1 0 27876 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1632082664
transform 1 0 26864 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_103_279
timestamp 1632082664
transform 1 0 26772 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_103_307
timestamp 1632082664
transform 1 0 29348 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0628_
timestamp 1632082664
transform 1 0 30176 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_103_315
timestamp 1632082664
transform 1 0 30084 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_332
timestamp 1632082664
transform 1 0 31648 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_103_349
timestamp 1632082664
transform 1 0 33212 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_103_337
timestamp 1632082664
transform 1 0 32108 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1632082664
transform 1 0 32016 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_53_clk
timestamp 1632082664
transform 1 0 33856 0 -1 58752
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_103_355
timestamp 1632082664
transform 1 0 33764 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_103_393
timestamp 1632082664
transform 1 0 37260 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0604_
timestamp 1632082664
transform 1 0 37444 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_103_376
timestamp 1632082664
transform 1 0 35696 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1632082664
transform 1 0 37168 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_388
timestamp 1632082664
transform 1 0 36800 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_103_411
timestamp 1632082664
transform 1 0 38916 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0558_
timestamp 1632082664
transform 1 0 40480 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_103_427
timestamp 1632082664
transform 1 0 40388 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_423
timestamp 1632082664
transform 1 0 40020 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_103_449
timestamp 1632082664
transform 1 0 42412 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1632082664
transform 1 0 42320 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_444
timestamp 1632082664
transform 1 0 41952 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0553_
timestamp 1632082664
transform 1 0 43792 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_103_461
timestamp 1632082664
transform 1 0 43516 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0549_
timestamp 1632082664
transform 1 0 45632 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_103_500
timestamp 1632082664
transform 1 0 47104 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_103_480
timestamp 1632082664
transform 1 0 45264 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_58_clk
timestamp 1632082664
transform 1 0 47932 0 -1 58752
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1632082664
transform 1 0 47472 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_505
timestamp 1632082664
transform 1 0 47564 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_103_529
timestamp 1632082664
transform 1 0 49772 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0533_
timestamp 1632082664
transform 1 0 50784 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_103_537
timestamp 1632082664
transform 1 0 50508 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_561
timestamp 1632082664
transform 1 0 52716 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1632082664
transform 1 0 52624 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_556
timestamp 1632082664
transform 1 0 52256 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0524_
timestamp 1632082664
transform 1 0 54096 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_103_573
timestamp 1632082664
transform 1 0 53820 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0521_
timestamp 1632082664
transform 1 0 55936 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_103_592
timestamp 1632082664
transform 1 0 55568 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_103_617
timestamp 1632082664
transform 1 0 57868 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1632082664
transform 1 0 57776 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_612
timestamp 1632082664
transform 1 0 57408 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_629
timestamp 1632082664
transform 1 0 58972 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1632082664
transform -1 0 59340 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_104_3
timestamp 1632082664
transform 1 0 1380 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_15
timestamp 1632082664
transform 1 0 2484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1632082664
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0863_
timestamp 1632082664
transform 1 0 4876 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_104_29
timestamp 1632082664
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1632082664
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1632082664
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0865_
timestamp 1632082664
transform 1 0 6716 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_104_57
timestamp 1632082664
transform 1 0 6348 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1632082664
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1632082664
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0871_
timestamp 1632082664
transform 1 0 8924 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1632082664
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_104_101
timestamp 1632082664
transform 1 0 10396 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0875_
timestamp 1632082664
transform 1 0 10764 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_104_121
timestamp 1632082664
transform 1 0 12236 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_133
timestamp 1632082664
transform 1 0 13340 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0883_
timestamp 1632082664
transform 1 0 14076 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1632082664
transform 1 0 13984 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_104_139
timestamp 1632082664
transform 1 0 13892 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0886_
timestamp 1632082664
transform 1 0 15916 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_104_157
timestamp 1632082664
transform 1 0 15548 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_104_177
timestamp 1632082664
transform 1 0 17388 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_189
timestamp 1632082664
transform 1 0 18492 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_104_197
timestamp 1632082664
transform 1 0 19228 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1632082664
transform 1 0 19136 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_104_195
timestamp 1632082664
transform 1 0 19044 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_104_209
timestamp 1632082664
transform 1 0 20332 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0654_
timestamp 1632082664
transform 1 0 20516 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_104_227
timestamp 1632082664
transform 1 0 21988 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0650_
timestamp 1632082664
transform 1 0 22448 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_104_231
timestamp 1632082664
transform 1 0 22356 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_104_248
timestamp 1632082664
transform 1 0 23920 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0642_
timestamp 1632082664
transform 1 0 25760 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_104_253
timestamp 1632082664
transform 1 0 24380 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1632082664
transform 1 0 24288 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_104_265
timestamp 1632082664
transform 1 0 25484 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0633_
timestamp 1632082664
transform 1 0 27600 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_104_284
timestamp 1632082664
transform 1 0 27232 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_104_309
timestamp 1632082664
transform 1 0 29532 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1632082664
transform 1 0 29440 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_104_304
timestamp 1632082664
transform 1 0 29072 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0626_
timestamp 1632082664
transform 1 0 30268 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_104_333
timestamp 1632082664
transform 1 0 31740 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_104_353
timestamp 1632082664
transform 1 0 33580 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0625_
timestamp 1632082664
transform 1 0 32108 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_104_365
timestamp 1632082664
transform 1 0 34684 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_104_373
timestamp 1632082664
transform 1 0 35420 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0611_
timestamp 1632082664
transform 1 0 35604 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1632082664
transform 1 0 34592 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_104_361
timestamp 1632082664
transform 1 0 34316 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_104_391
timestamp 1632082664
transform 1 0 37076 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_104_413
timestamp 1632082664
transform 1 0 39100 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0606_
timestamp 1632082664
transform 1 0 37628 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0557_
timestamp 1632082664
transform 1 0 41216 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_104_421
timestamp 1632082664
transform 1 0 39836 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1632082664
transform 1 0 39744 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_104_419
timestamp 1632082664
transform 1 0 39652 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_104_433
timestamp 1632082664
transform 1 0 40940 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0554_
timestamp 1632082664
transform 1 0 43056 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_104_452
timestamp 1632082664
transform 1 0 42688 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_104_477
timestamp 1632082664
transform 1 0 44988 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1632082664
transform 1 0 44896 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_104_472
timestamp 1632082664
transform 1 0 44528 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0548_
timestamp 1632082664
transform 1 0 46368 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_104_489
timestamp 1632082664
transform 1 0 46092 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0544_
timestamp 1632082664
transform 1 0 48208 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_104_508
timestamp 1632082664
transform 1 0 47840 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_104_533
timestamp 1632082664
transform 1 0 50140 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1632082664
transform 1 0 50048 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_104_528
timestamp 1632082664
transform 1 0 49680 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0530_
timestamp 1632082664
transform 1 0 51520 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_104_545
timestamp 1632082664
transform 1 0 51244 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0526_
timestamp 1632082664
transform 1 0 53360 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_104_564
timestamp 1632082664
transform 1 0 52992 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1182_
timestamp 1632082664
transform 1 0 55292 0 1 58752
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1632082664
transform 1 0 55200 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_104_584
timestamp 1632082664
transform 1 0 54832 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0520_
timestamp 1632082664
transform 1 0 57224 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_104_606
timestamp 1632082664
transform 1 0 56856 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_104_626
timestamp 1632082664
transform 1 0 58696 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1632082664
transform -1 0 59340 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_106_3
timestamp 1632082664
transform 1 0 1380 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_15
timestamp 1632082664
transform 1 0 2484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_3
timestamp 1632082664
transform 1 0 1380 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_15
timestamp 1632082664
transform 1 0 2484 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1632082664
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1632082664
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_106_41
timestamp 1632082664
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_29
timestamp 1632082664
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_39
timestamp 1632082664
transform 1 0 4692 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_27
timestamp 1632082664
transform 1 0 3588 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1632082664
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1632082664
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _0867_
timestamp 1632082664
transform 1 0 6440 0 1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0866_
timestamp 1632082664
transform 1 0 6348 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1632082664
transform 1 0 6256 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1632082664
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_106_57
timestamp 1632082664
transform 1 0 6348 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1632082664
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_51
timestamp 1632082664
transform 1 0 5796 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_106_53
timestamp 1632082664
transform 1 0 5980 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_106_74
timestamp 1632082664
transform 1 0 7912 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_106_82
timestamp 1632082664
transform 1 0 8648 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0870_
timestamp 1632082664
transform 1 0 8188 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_105_73
timestamp 1632082664
transform 1 0 7820 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_106_97
timestamp 1632082664
transform 1 0 10028 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_85
timestamp 1632082664
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_93
timestamp 1632082664
transform 1 0 9660 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1632082664
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_105_105
timestamp 1632082664
transform 1 0 10764 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_106_113
timestamp 1632082664
transform 1 0 11500 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0879_
timestamp 1632082664
transform 1 0 11684 0 1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0878_
timestamp 1632082664
transform 1 0 11500 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1632082664
transform 1 0 11408 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1632082664
transform 1 0 11408 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_105_111
timestamp 1632082664
transform 1 0 11316 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_106_109
timestamp 1632082664
transform 1 0 11132 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_106_131
timestamp 1632082664
transform 1 0 13156 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0882_
timestamp 1632082664
transform 1 0 13340 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_106_141
timestamp 1632082664
transform 1 0 14076 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1632082664
transform 1 0 13984 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_106_139
timestamp 1632082664
transform 1 0 13892 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_129
timestamp 1632082664
transform 1 0 12972 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_105_161
timestamp 1632082664
transform 1 0 15916 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_106_153
timestamp 1632082664
transform 1 0 15180 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_149
timestamp 1632082664
transform 1 0 14812 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_165
timestamp 1632082664
transform 1 0 16284 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_106_181
timestamp 1632082664
transform 1 0 17756 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_169
timestamp 1632082664
transform 1 0 16652 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_181
timestamp 1632082664
transform 1 0 17756 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_169
timestamp 1632082664
transform 1 0 16652 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1632082664
transform 1 0 16560 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1632082664
transform 1 0 16560 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_105_167
timestamp 1632082664
transform 1 0 16468 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_105_193
timestamp 1632082664
transform 1 0 18860 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0656_
timestamp 1632082664
transform 1 0 19872 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_106_197
timestamp 1632082664
transform 1 0 19228 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1632082664
transform 1 0 19136 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_106_193
timestamp 1632082664
transform 1 0 18860 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_105_201
timestamp 1632082664
transform 1 0 19596 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_105_225
timestamp 1632082664
transform 1 0 21804 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_106_225
timestamp 1632082664
transform 1 0 21804 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_209
timestamp 1632082664
transform 1 0 20332 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1632082664
transform 1 0 21712 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1632082664
transform 1 0 21712 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_220
timestamp 1632082664
transform 1 0 21344 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_106_221
timestamp 1632082664
transform 1 0 21436 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0651_
timestamp 1632082664
transform 1 0 22448 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_106_237
timestamp 1632082664
transform 1 0 22908 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_231
timestamp 1632082664
transform 1 0 22356 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_248
timestamp 1632082664
transform 1 0 23920 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_106_249
timestamp 1632082664
transform 1 0 24012 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0645_
timestamp 1632082664
transform 1 0 24288 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_106_265
timestamp 1632082664
transform 1 0 25484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_253
timestamp 1632082664
transform 1 0 24380 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_268
timestamp 1632082664
transform 1 0 25760 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1632082664
transform 1 0 24288 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1632082664
transform -1 0 27324 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_106_281
timestamp 1632082664
transform 1 0 26956 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0641_
timestamp 1632082664
transform 1 0 26956 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_106_289
timestamp 1632082664
transform 1 0 27692 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1632082664
transform 1 0 26864 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1632082664
transform 1 0 26864 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output3
timestamp 1632082664
transform -1 0 27692 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_106_277
timestamp 1632082664
transform 1 0 26588 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_106_301
timestamp 1632082664
transform 1 0 28796 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_105_309
timestamp 1632082664
transform 1 0 29532 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_105_297
timestamp 1632082664
transform 1 0 28428 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1632082664
transform 1 0 29440 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_106_307
timestamp 1632082664
transform 1 0 29348 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_309
timestamp 1632082664
transform 1 0 29532 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_106_329
timestamp 1632082664
transform 1 0 31372 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0632_
timestamp 1632082664
transform 1 0 29900 0 1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0630_
timestamp 1632082664
transform 1 0 30176 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_105_315
timestamp 1632082664
transform 1 0 30084 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_332
timestamp 1632082664
transform 1 0 31648 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_106_353
timestamp 1632082664
transform 1 0 33580 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0631_
timestamp 1632082664
transform 1 0 32108 0 1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0629_
timestamp 1632082664
transform 1 0 32568 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1632082664
transform 1 0 32016 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1632082664
transform 1 0 32016 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_106_335
timestamp 1632082664
transform 1 0 31924 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_105_341
timestamp 1632082664
transform 1 0 32476 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_337
timestamp 1632082664
transform 1 0 32108 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_106_365
timestamp 1632082664
transform 1 0 34684 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0613_
timestamp 1632082664
transform 1 0 34408 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0610_
timestamp 1632082664
transform 1 0 35328 0 1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1632082664
transform 1 0 34592 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_106_371
timestamp 1632082664
transform 1 0 35236 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_358
timestamp 1632082664
transform 1 0 34040 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_106_361
timestamp 1632082664
transform 1 0 34316 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_106_393
timestamp 1632082664
transform 1 0 37260 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_390
timestamp 1632082664
transform 1 0 36984 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0608_
timestamp 1632082664
transform 1 0 37444 0 1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_105_378
timestamp 1632082664
transform 1 0 35880 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1632082664
transform 1 0 37168 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1632082664
transform 1 0 37168 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_388
timestamp 1632082664
transform 1 0 36800 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_105_393
timestamp 1632082664
transform 1 0 37260 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_106_411
timestamp 1632082664
transform 1 0 38916 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0607_
timestamp 1632082664
transform 1 0 37536 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_105_412
timestamp 1632082664
transform 1 0 39008 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_437
timestamp 1632082664
transform 1 0 41308 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0609_
timestamp 1632082664
transform 1 0 39836 0 1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0559_
timestamp 1632082664
transform 1 0 40388 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1632082664
transform 1 0 39744 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_106_419
timestamp 1632082664
transform 1 0 39652 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_105_424
timestamp 1632082664
transform 1 0 40112 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_106_449
timestamp 1632082664
transform 1 0 42412 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_449
timestamp 1632082664
transform 1 0 42412 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1632082664
transform 1 0 42320 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1632082664
transform 1 0 42320 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_105_447
timestamp 1632082664
transform 1 0 42228 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_443
timestamp 1632082664
transform 1 0 41860 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_106_445
timestamp 1632082664
transform 1 0 42044 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0555_
timestamp 1632082664
transform 1 0 43608 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0552_
timestamp 1632082664
transform 1 0 44988 0 1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_106_461
timestamp 1632082664
transform 1 0 43516 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1632082664
transform 1 0 44896 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_105_461
timestamp 1632082664
transform 1 0 43516 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_478
timestamp 1632082664
transform 1 0 45080 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_106_473
timestamp 1632082664
transform 1 0 44620 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_106_493
timestamp 1632082664
transform 1 0 46460 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0551_
timestamp 1632082664
transform 1 0 45540 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_105_482
timestamp 1632082664
transform 1 0 45448 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_499
timestamp 1632082664
transform 1 0 47012 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_106_505
timestamp 1632082664
transform 1 0 47564 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_517
timestamp 1632082664
transform 1 0 48668 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0546_
timestamp 1632082664
transform 1 0 47748 0 1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0542_
timestamp 1632082664
transform 1 0 48852 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_105_505
timestamp 1632082664
transform 1 0 47564 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1632082664
transform 1 0 47472 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1632082664
transform 1 0 47472 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_105_503
timestamp 1632082664
transform 1 0 47380 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_106_501
timestamp 1632082664
transform 1 0 47196 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_106_523
timestamp 1632082664
transform 1 0 49220 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0540_
timestamp 1632082664
transform 1 0 50140 0 1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0536_
timestamp 1632082664
transform 1 0 50784 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1632082664
transform 1 0 50048 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_106_531
timestamp 1632082664
transform 1 0 49956 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_105_539
timestamp 1632082664
transform 1 0 50692 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_535
timestamp 1632082664
transform 1 0 50324 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_106_561
timestamp 1632082664
transform 1 0 52716 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_106_549
timestamp 1632082664
transform 1 0 51612 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_105_561
timestamp 1632082664
transform 1 0 52716 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1632082664
transform 1 0 52624 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1632082664
transform 1 0 52624 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_556
timestamp 1632082664
transform 1 0 52256 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_106_557
timestamp 1632082664
transform 1 0 52348 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0529_
timestamp 1632082664
transform 1 0 53360 0 1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0527_
timestamp 1632082664
transform 1 0 53544 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_106_567
timestamp 1632082664
transform 1 0 53268 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_105_569
timestamp 1632082664
transform 1 0 53452 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_105_586
timestamp 1632082664
transform 1 0 55016 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_594
timestamp 1632082664
transform 1 0 55752 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _0523_
timestamp 1632082664
transform 1 0 55936 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_106_601
timestamp 1632082664
transform 1 0 56396 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_589
timestamp 1632082664
transform 1 0 55292 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1632082664
transform 1 0 55200 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_584
timestamp 1632082664
transform 1 0 54832 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_105_617
timestamp 1632082664
transform 1 0 57868 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1632082664
transform 1 0 57776 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1632082664
transform 1 0 57776 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output4
timestamp 1632082664
transform 1 0 58328 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_621
timestamp 1632082664
transform 1 0 58236 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_617
timestamp 1632082664
transform 1 0 57868 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_105_612
timestamp 1632082664
transform 1 0 57408 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_106_613
timestamp 1632082664
transform 1 0 57500 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_105_629
timestamp 1632082664
transform 1 0 58972 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_626
timestamp 1632082664
transform 1 0 58696 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1632082664
transform -1 0 59340 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1632082664
transform -1 0 59340 0 -1 59840
box -38 -48 314 592
<< labels >>
rlabel metal5 s 1104 20616 59340 20936 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 5298 59340 5618 6 VPWR
port 1 nsew power input
rlabel metal3 s 0 50600 800 50720 6 clk
port 2 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 din
port 3 nsew signal input
rlabel metal2 s 18 0 74 800 6 out_window[0]
port 4 nsew signal tristate
rlabel metal2 s 26146 61860 26202 62660 6 out_window[1]
port 5 nsew signal tristate
rlabel metal2 s 60370 61860 60426 62660 6 out_window[2]
port 6 nsew signal tristate
rlabel metal3 s 59716 11704 60516 11824 6 out_window[3]
port 7 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 60516 62660
<< end >>
