magic
tech sky130A
timestamp 1640659972
<< nwell >>
rect 65035 278750 65595 278895
<< nmos >>
rect 65095 278670 65110 278715
rect 65275 278515 65290 278615
rect 65465 278515 65480 278615
<< pmos >>
rect 65095 278810 65110 278855
rect 65275 278770 65290 278870
rect 65465 278770 65480 278870
<< ndiff >>
rect 65060 278705 65095 278715
rect 65060 278680 65065 278705
rect 65085 278680 65095 278705
rect 65060 278670 65095 278680
rect 65110 278705 65145 278715
rect 65110 278680 65120 278705
rect 65140 278680 65145 278705
rect 65110 278670 65145 278680
rect 65240 278605 65275 278615
rect 65240 278525 65245 278605
rect 65265 278525 65275 278605
rect 65240 278515 65275 278525
rect 65290 278605 65325 278615
rect 65290 278525 65300 278605
rect 65320 278525 65325 278605
rect 65290 278515 65325 278525
rect 65430 278605 65465 278615
rect 65430 278525 65435 278605
rect 65455 278525 65465 278605
rect 65430 278515 65465 278525
rect 65480 278605 65515 278615
rect 65480 278525 65490 278605
rect 65510 278525 65515 278605
rect 65480 278515 65515 278525
<< pdiff >>
rect 65240 278860 65275 278870
rect 65060 278845 65095 278855
rect 65060 278820 65065 278845
rect 65085 278820 65095 278845
rect 65060 278810 65095 278820
rect 65110 278845 65145 278855
rect 65110 278820 65120 278845
rect 65140 278820 65145 278845
rect 65110 278810 65145 278820
rect 65240 278780 65245 278860
rect 65265 278780 65275 278860
rect 65240 278770 65275 278780
rect 65290 278860 65325 278870
rect 65290 278780 65300 278860
rect 65320 278780 65325 278860
rect 65290 278770 65325 278780
rect 65430 278860 65465 278870
rect 65430 278780 65435 278860
rect 65455 278780 65465 278860
rect 65430 278770 65465 278780
rect 65480 278860 65515 278870
rect 65480 278780 65490 278860
rect 65510 278780 65515 278860
rect 65480 278770 65515 278780
<< ndiffc >>
rect 65065 278680 65085 278705
rect 65120 278680 65140 278705
rect 65245 278525 65265 278605
rect 65300 278525 65320 278605
rect 65435 278525 65455 278605
rect 65490 278525 65510 278605
<< pdiffc >>
rect 65065 278820 65085 278845
rect 65120 278820 65140 278845
rect 65245 278780 65265 278860
rect 65300 278780 65320 278860
rect 65435 278780 65455 278860
rect 65490 278780 65510 278860
<< psubdiff >>
rect 65185 278605 65240 278615
rect 65185 278525 65200 278605
rect 65220 278525 65240 278605
rect 65185 278515 65240 278525
rect 65515 278605 65570 278615
rect 65515 278525 65535 278605
rect 65555 278525 65570 278605
rect 65515 278515 65570 278525
<< nsubdiff >>
rect 65185 278860 65240 278870
rect 65185 278780 65200 278860
rect 65220 278780 65240 278860
rect 65185 278770 65240 278780
rect 65515 278860 65570 278870
rect 65515 278780 65535 278860
rect 65555 278780 65570 278860
rect 65515 278770 65570 278780
<< psubdiffcont >>
rect 65200 278525 65220 278605
rect 65535 278525 65555 278605
<< nsubdiffcont >>
rect 65200 278780 65220 278860
rect 65535 278780 65555 278860
<< poly >>
rect 64980 278940 65020 278950
rect 64980 278920 64990 278940
rect 65010 278935 65020 278940
rect 65010 278920 65480 278935
rect 64980 278910 65020 278920
rect 65095 278855 65110 278920
rect 65275 278870 65290 278885
rect 65465 278870 65480 278920
rect 65095 278715 65110 278810
rect 65165 278740 65205 278750
rect 65275 278740 65290 278770
rect 65355 278745 65395 278755
rect 65355 278740 65365 278745
rect 65165 278720 65175 278740
rect 65195 278725 65365 278740
rect 65385 278725 65395 278745
rect 65195 278720 65205 278725
rect 65165 278710 65205 278720
rect 65355 278715 65395 278725
rect 65465 278690 65480 278770
rect 65540 278740 65580 278750
rect 65540 278720 65550 278740
rect 65570 278720 65580 278740
rect 65540 278710 65580 278720
rect 65275 278675 65480 278690
rect 65095 278655 65110 278670
rect 65275 278615 65290 278675
rect 65550 278650 65565 278710
rect 65465 278635 65565 278650
rect 65465 278615 65480 278635
rect 65275 278500 65290 278515
rect 65465 278500 65480 278515
<< polycont >>
rect 64990 278920 65010 278940
rect 65175 278720 65195 278740
rect 65365 278725 65385 278745
rect 65550 278720 65570 278740
<< locali >>
rect 65145 279005 65175 279010
rect 65140 279000 65180 279005
rect 65140 278970 65145 279000
rect 65175 278970 65180 279000
rect 65140 278965 65180 278970
rect 64980 278945 65020 278950
rect 64980 278915 64985 278945
rect 65015 278915 65020 278945
rect 65145 278920 65175 278965
rect 64980 278910 65020 278915
rect 65060 278895 65555 278920
rect 65060 278845 65090 278895
rect 65200 278860 65220 278895
rect 65060 278820 65065 278845
rect 65085 278820 65090 278845
rect 65060 278810 65090 278820
rect 65115 278845 65145 278855
rect 65115 278820 65120 278845
rect 65140 278820 65145 278845
rect 65115 278745 65145 278820
rect 65200 278770 65220 278780
rect 65240 278860 65270 278870
rect 65240 278780 65245 278860
rect 65265 278780 65270 278860
rect 65165 278745 65205 278750
rect 65115 278740 65205 278745
rect 65115 278720 65175 278740
rect 65195 278720 65205 278740
rect 65060 278705 65090 278715
rect 65060 278680 65065 278705
rect 65085 278680 65090 278705
rect 65060 278670 65090 278680
rect 65115 278705 65145 278720
rect 65165 278710 65205 278720
rect 65115 278680 65120 278705
rect 65140 278680 65145 278705
rect 65115 278670 65145 278680
rect 65240 278665 65270 278780
rect 65200 278605 65220 278615
rect 65060 278490 65100 278495
rect 65200 278490 65220 278525
rect 65240 278605 65270 278635
rect 65240 278525 65245 278605
rect 65265 278525 65270 278605
rect 65240 278515 65270 278525
rect 65295 278860 65325 278870
rect 65295 278780 65300 278860
rect 65320 278780 65325 278860
rect 65295 278665 65325 278780
rect 65430 278860 65460 278870
rect 65430 278780 65435 278860
rect 65455 278780 65460 278860
rect 65355 278750 65395 278755
rect 65355 278720 65360 278750
rect 65390 278720 65395 278750
rect 65355 278715 65395 278720
rect 65355 278665 65395 278670
rect 65430 278665 65460 278780
rect 65295 278635 65360 278665
rect 65390 278635 65460 278665
rect 65295 278605 65325 278635
rect 65355 278630 65395 278635
rect 65295 278525 65300 278605
rect 65320 278525 65325 278605
rect 65295 278515 65325 278525
rect 65430 278605 65460 278635
rect 65430 278525 65435 278605
rect 65455 278525 65460 278605
rect 65430 278515 65460 278525
rect 65485 278860 65515 278870
rect 65485 278780 65490 278860
rect 65510 278780 65515 278860
rect 65485 278605 65515 278780
rect 65535 278860 65555 278895
rect 65535 278770 65555 278780
rect 65540 278745 65580 278750
rect 65540 278715 65545 278745
rect 65575 278715 65580 278745
rect 65540 278710 65580 278715
rect 65485 278525 65490 278605
rect 65510 278525 65515 278605
rect 65485 278490 65515 278525
rect 65535 278605 65555 278615
rect 65535 278490 65555 278525
rect 65055 278460 65065 278490
rect 65095 278460 65555 278490
rect 65060 278455 65100 278460
<< viali >>
rect 65145 278970 65175 279000
rect 64985 278940 65015 278945
rect 64985 278920 64990 278940
rect 64990 278920 65010 278940
rect 65010 278920 65015 278940
rect 64985 278915 65015 278920
rect 65065 278680 65085 278705
rect 65240 278635 65270 278665
rect 65360 278745 65390 278750
rect 65360 278725 65365 278745
rect 65365 278725 65385 278745
rect 65385 278725 65390 278745
rect 65360 278720 65390 278725
rect 65360 278635 65390 278665
rect 65545 278740 65575 278745
rect 65545 278720 65550 278740
rect 65550 278720 65570 278740
rect 65570 278720 65575 278740
rect 65545 278715 65575 278720
rect 65065 278460 65095 278490
<< metal1 >>
rect 64975 278945 65025 279060
rect 64975 278915 64985 278945
rect 65015 278915 65025 278945
rect 64975 278905 65025 278915
rect 65055 278705 65105 279060
rect 65135 279000 65185 279060
rect 65135 278970 65145 279000
rect 65175 278970 65185 279000
rect 65135 278960 65185 278970
rect 65350 278750 65400 278760
rect 65535 278750 65585 278755
rect 65350 278720 65360 278750
rect 65390 278745 65585 278750
rect 65390 278720 65545 278745
rect 65350 278710 65400 278720
rect 65535 278715 65545 278720
rect 65575 278715 65585 278745
rect 65535 278705 65585 278715
rect 65055 278680 65065 278705
rect 65085 278680 65105 278705
rect 65055 278490 65105 278680
rect 65230 278670 65280 278675
rect 65230 278630 65235 278670
rect 65275 278630 65280 278670
rect 65230 278625 65280 278630
rect 65350 278665 65840 278675
rect 65350 278635 65360 278665
rect 65390 278635 65840 278665
rect 65350 278625 65840 278635
rect 65055 278460 65065 278490
rect 65095 278460 65105 278490
rect 65055 278455 65105 278460
<< via1 >>
rect 65235 278665 65275 278670
rect 65235 278635 65240 278665
rect 65240 278635 65270 278665
rect 65270 278635 65275 278665
rect 65235 278630 65275 278635
<< metal2 >>
rect 64775 278670 65280 278675
rect 64775 278630 64780 278670
rect 64825 278630 65235 278670
rect 65275 278630 65280 278670
rect 64775 278625 65280 278630
<< via2 >>
rect 64780 278630 64825 278670
<< metal3 >>
rect 64775 278670 64830 278675
rect 64775 278630 64780 278670
rect 64825 278630 64830 278670
rect 64775 278625 64830 278630
<< via3 >>
rect 64780 278630 64825 278670
<< via4 >>
rect 64740 278670 64860 278710
rect 64740 278630 64780 278670
rect 64780 278630 64825 278670
rect 64825 278630 64860 278670
rect 64740 278590 64860 278630
<< metal5 >>
rect 64610 278710 65010 278855
rect 64610 278590 64740 278710
rect 64860 278590 65010 278710
rect 64610 278455 65010 278590
<< labels >>
rlabel metal1 65001 279060 65001 279060 5 SIgnal
rlabel metal1 65079 279059 65079 279059 5 GND
rlabel metal1 65159 279060 65159 279060 5 VDD
<< end >>
